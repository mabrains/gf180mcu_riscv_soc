magic
tech gf180mcuD
magscale 1 10
timestamp 1700584958
<< metal1 >>
rect 1344 98026 38640 98060
rect 1344 97974 4478 98026
rect 4530 97974 4582 98026
rect 4634 97974 4686 98026
rect 4738 97974 35198 98026
rect 35250 97974 35302 98026
rect 35354 97974 35406 98026
rect 35458 97974 38640 98026
rect 1344 97940 38640 97974
rect 14466 97582 14478 97634
rect 14530 97582 14542 97634
rect 15250 97582 15262 97634
rect 15314 97582 15326 97634
rect 13022 97522 13074 97534
rect 13022 97458 13074 97470
rect 1710 97410 1762 97422
rect 1710 97346 1762 97358
rect 4062 97410 4114 97422
rect 4062 97346 4114 97358
rect 6526 97410 6578 97422
rect 6526 97346 6578 97358
rect 9326 97410 9378 97422
rect 9326 97346 9378 97358
rect 11454 97410 11506 97422
rect 11454 97346 11506 97358
rect 15710 97410 15762 97422
rect 15710 97346 15762 97358
rect 16270 97410 16322 97422
rect 16270 97346 16322 97358
rect 16942 97410 16994 97422
rect 16942 97346 16994 97358
rect 18846 97410 18898 97422
rect 18846 97346 18898 97358
rect 1344 97242 38640 97276
rect 1344 97190 19838 97242
rect 19890 97190 19942 97242
rect 19994 97190 20046 97242
rect 20098 97190 38640 97242
rect 1344 97156 38640 97190
rect 14702 96850 14754 96862
rect 32286 96850 32338 96862
rect 7970 96798 7982 96850
rect 8034 96798 8046 96850
rect 8866 96798 8878 96850
rect 8930 96798 8942 96850
rect 13906 96798 13918 96850
rect 13970 96798 13982 96850
rect 31266 96798 31278 96850
rect 31330 96798 31342 96850
rect 34290 96798 34302 96850
rect 34354 96798 34366 96850
rect 35186 96798 35198 96850
rect 35250 96798 35262 96850
rect 14702 96786 14754 96798
rect 32286 96786 32338 96798
rect 9662 96738 9714 96750
rect 9662 96674 9714 96686
rect 10110 96738 10162 96750
rect 10110 96674 10162 96686
rect 12350 96738 12402 96750
rect 12350 96674 12402 96686
rect 15150 96738 15202 96750
rect 15150 96674 15202 96686
rect 6862 96626 6914 96638
rect 6862 96562 6914 96574
rect 30158 96626 30210 96638
rect 30158 96562 30210 96574
rect 33182 96626 33234 96638
rect 33182 96562 33234 96574
rect 1344 96458 38640 96492
rect 1344 96406 4478 96458
rect 4530 96406 4582 96458
rect 4634 96406 4686 96458
rect 4738 96406 35198 96458
rect 35250 96406 35302 96458
rect 35354 96406 35406 96458
rect 35458 96406 38640 96458
rect 1344 96372 38640 96406
rect 15598 96290 15650 96302
rect 15598 96226 15650 96238
rect 19518 96290 19570 96302
rect 19518 96226 19570 96238
rect 23438 96290 23490 96302
rect 23438 96226 23490 96238
rect 16158 96178 16210 96190
rect 16158 96114 16210 96126
rect 9326 96066 9378 96078
rect 2930 96014 2942 96066
rect 2994 96014 3006 96066
rect 3826 96014 3838 96066
rect 3890 96014 3902 96066
rect 6738 96014 6750 96066
rect 6802 96014 6814 96066
rect 7634 96014 7646 96066
rect 7698 96014 7710 96066
rect 10322 96014 10334 96066
rect 10386 96014 10398 96066
rect 13570 96014 13582 96066
rect 13634 96014 13646 96066
rect 14466 96014 14478 96066
rect 14530 96014 14542 96066
rect 17490 96014 17502 96066
rect 17554 96014 17566 96066
rect 18386 96014 18398 96066
rect 18450 96014 18462 96066
rect 21410 96014 21422 96066
rect 21474 96014 21486 96066
rect 22306 96014 22318 96066
rect 22370 96014 22382 96066
rect 29250 96014 29262 96066
rect 29314 96014 29326 96066
rect 30146 96014 30158 96066
rect 30210 96014 30222 96066
rect 32946 96014 32958 96066
rect 33010 96014 33022 96066
rect 33842 96014 33854 96066
rect 33906 96014 33918 96066
rect 9326 96002 9378 96014
rect 25006 95954 25058 95966
rect 8642 95902 8654 95954
rect 8706 95902 8718 95954
rect 24210 95902 24222 95954
rect 24274 95902 24286 95954
rect 25006 95890 25058 95902
rect 25342 95954 25394 95966
rect 25342 95890 25394 95902
rect 26462 95954 26514 95966
rect 26462 95890 26514 95902
rect 26798 95954 26850 95966
rect 26798 95890 26850 95902
rect 5182 95842 5234 95854
rect 5182 95778 5234 95790
rect 5742 95842 5794 95854
rect 5742 95778 5794 95790
rect 11678 95842 11730 95854
rect 11678 95778 11730 95790
rect 12014 95842 12066 95854
rect 12014 95778 12066 95790
rect 20078 95842 20130 95854
rect 20078 95778 20130 95790
rect 20750 95842 20802 95854
rect 20750 95778 20802 95790
rect 23886 95842 23938 95854
rect 23886 95778 23938 95790
rect 25678 95842 25730 95854
rect 27358 95842 27410 95854
rect 26002 95790 26014 95842
rect 26066 95790 26078 95842
rect 25678 95778 25730 95790
rect 27358 95778 27410 95790
rect 31502 95842 31554 95854
rect 31502 95778 31554 95790
rect 35198 95842 35250 95854
rect 35198 95778 35250 95790
rect 1344 95674 38640 95708
rect 1344 95622 19838 95674
rect 19890 95622 19942 95674
rect 19994 95622 20046 95674
rect 20098 95622 38640 95674
rect 1344 95588 38640 95622
rect 6190 95506 6242 95518
rect 6190 95442 6242 95454
rect 9662 95506 9714 95518
rect 9662 95442 9714 95454
rect 12350 95506 12402 95518
rect 12350 95442 12402 95454
rect 15150 95506 15202 95518
rect 15150 95442 15202 95454
rect 16818 95342 16830 95394
rect 16882 95342 16894 95394
rect 6750 95282 6802 95294
rect 14702 95282 14754 95294
rect 3938 95230 3950 95282
rect 4002 95230 4014 95282
rect 4834 95230 4846 95282
rect 4898 95230 4910 95282
rect 7634 95230 7646 95282
rect 7698 95230 7710 95282
rect 13906 95230 13918 95282
rect 13970 95230 13982 95282
rect 6750 95218 6802 95230
rect 14702 95218 14754 95230
rect 16494 95282 16546 95294
rect 22206 95282 22258 95294
rect 17490 95230 17502 95282
rect 17554 95230 17566 95282
rect 18386 95230 18398 95282
rect 18450 95230 18462 95282
rect 21186 95230 21198 95282
rect 21250 95230 21262 95282
rect 16494 95218 16546 95230
rect 22206 95218 22258 95230
rect 24670 95282 24722 95294
rect 33070 95282 33122 95294
rect 35646 95282 35698 95294
rect 25330 95230 25342 95282
rect 25394 95230 25406 95282
rect 26002 95230 26014 95282
rect 26066 95230 26078 95282
rect 28242 95230 28254 95282
rect 28306 95230 28318 95282
rect 29138 95230 29150 95282
rect 29202 95230 29214 95282
rect 34066 95230 34078 95282
rect 34130 95230 34142 95282
rect 36418 95230 36430 95282
rect 36482 95230 36494 95282
rect 24670 95218 24722 95230
rect 33070 95218 33122 95230
rect 35646 95218 35698 95230
rect 9102 95170 9154 95182
rect 9102 95106 9154 95118
rect 19854 95170 19906 95182
rect 19854 95106 19906 95118
rect 23550 95170 23602 95182
rect 23550 95106 23602 95118
rect 30494 95170 30546 95182
rect 30494 95106 30546 95118
rect 19518 95058 19570 95070
rect 19518 94994 19570 95006
rect 27358 95058 27410 95070
rect 27358 94994 27410 95006
rect 35198 95058 35250 95070
rect 35198 94994 35250 95006
rect 37774 95058 37826 95070
rect 37774 94994 37826 95006
rect 1344 94890 38640 94924
rect 1344 94838 4478 94890
rect 4530 94838 4582 94890
rect 4634 94838 4686 94890
rect 4738 94838 35198 94890
rect 35250 94838 35302 94890
rect 35354 94838 35406 94890
rect 35458 94838 38640 94890
rect 1344 94804 38640 94838
rect 4958 94722 5010 94734
rect 4958 94658 5010 94670
rect 20638 94722 20690 94734
rect 20638 94658 20690 94670
rect 25342 94722 25394 94734
rect 25342 94658 25394 94670
rect 34974 94722 35026 94734
rect 34974 94658 35026 94670
rect 5742 94610 5794 94622
rect 5742 94546 5794 94558
rect 6302 94610 6354 94622
rect 6302 94546 6354 94558
rect 15598 94610 15650 94622
rect 26238 94610 26290 94622
rect 15922 94558 15934 94610
rect 15986 94558 15998 94610
rect 22194 94558 22206 94610
rect 22258 94558 22270 94610
rect 15598 94546 15650 94558
rect 26238 94546 26290 94558
rect 16718 94498 16770 94510
rect 2930 94446 2942 94498
rect 2994 94446 3006 94498
rect 3826 94446 3838 94498
rect 3890 94446 3902 94498
rect 16146 94446 16158 94498
rect 16210 94446 16222 94498
rect 16718 94434 16770 94446
rect 18510 94498 18562 94510
rect 22654 94498 22706 94510
rect 19282 94446 19294 94498
rect 19346 94446 19358 94498
rect 21522 94446 21534 94498
rect 21586 94446 21598 94498
rect 22306 94446 22318 94498
rect 22370 94446 22382 94498
rect 18510 94434 18562 94446
rect 22654 94434 22706 94446
rect 25006 94498 25058 94510
rect 25678 94498 25730 94510
rect 28590 94498 28642 94510
rect 32846 94498 32898 94510
rect 25330 94446 25342 94498
rect 25394 94446 25406 94498
rect 27794 94446 27806 94498
rect 27858 94446 27870 94498
rect 29250 94446 29262 94498
rect 29314 94446 29326 94498
rect 30146 94446 30158 94498
rect 30210 94446 30222 94498
rect 33842 94446 33854 94498
rect 33906 94446 33918 94498
rect 25006 94434 25058 94446
rect 25678 94434 25730 94446
rect 28590 94434 28642 94446
rect 32846 94434 32898 94446
rect 1710 94386 1762 94398
rect 1710 94322 1762 94334
rect 16830 94386 16882 94398
rect 16830 94322 16882 94334
rect 21982 94386 22034 94398
rect 21982 94322 22034 94334
rect 22766 94386 22818 94398
rect 22766 94322 22818 94334
rect 24334 94386 24386 94398
rect 24334 94322 24386 94334
rect 25790 94386 25842 94398
rect 25790 94322 25842 94334
rect 17278 94274 17330 94286
rect 17278 94210 17330 94222
rect 17726 94274 17778 94286
rect 17726 94210 17778 94222
rect 21310 94274 21362 94286
rect 21310 94210 21362 94222
rect 23214 94274 23266 94286
rect 23214 94210 23266 94222
rect 24110 94274 24162 94286
rect 24110 94210 24162 94222
rect 24670 94274 24722 94286
rect 24670 94210 24722 94222
rect 31502 94274 31554 94286
rect 31502 94210 31554 94222
rect 1344 94106 38640 94140
rect 1344 94054 19838 94106
rect 19890 94054 19942 94106
rect 19994 94054 20046 94106
rect 20098 94054 38640 94106
rect 1344 94020 38640 94054
rect 4622 93938 4674 93950
rect 4622 93874 4674 93886
rect 9102 93938 9154 93950
rect 23326 93938 23378 93950
rect 16258 93886 16270 93938
rect 16322 93886 16334 93938
rect 20626 93886 20638 93938
rect 20690 93886 20702 93938
rect 9102 93874 9154 93886
rect 23326 93874 23378 93886
rect 13246 93826 13298 93838
rect 13246 93762 13298 93774
rect 4174 93714 4226 93726
rect 3378 93662 3390 93714
rect 3442 93662 3454 93714
rect 4174 93650 4226 93662
rect 6750 93714 6802 93726
rect 13358 93714 13410 93726
rect 7634 93662 7646 93714
rect 7698 93662 7710 93714
rect 12002 93662 12014 93714
rect 12066 93662 12078 93714
rect 6750 93650 6802 93662
rect 13358 93650 13410 93662
rect 16606 93714 16658 93726
rect 16606 93650 16658 93662
rect 16830 93714 16882 93726
rect 20302 93714 20354 93726
rect 17490 93662 17502 93714
rect 17554 93662 17566 93714
rect 18386 93662 18398 93714
rect 18450 93662 18462 93714
rect 16830 93650 16882 93662
rect 20302 93650 20354 93662
rect 20974 93714 21026 93726
rect 25230 93714 25282 93726
rect 21970 93662 21982 93714
rect 22034 93662 22046 93714
rect 23874 93662 23886 93714
rect 23938 93662 23950 93714
rect 26002 93662 26014 93714
rect 26066 93662 26078 93714
rect 28802 93662 28814 93714
rect 28866 93662 28878 93714
rect 29586 93662 29598 93714
rect 29650 93662 29662 93714
rect 33170 93662 33182 93714
rect 33234 93662 33246 93714
rect 33842 93662 33854 93714
rect 33906 93662 33918 93714
rect 20974 93650 21026 93662
rect 25230 93650 25282 93662
rect 9662 93602 9714 93614
rect 20078 93602 20130 93614
rect 24558 93602 24610 93614
rect 12674 93550 12686 93602
rect 12738 93550 12750 93602
rect 23986 93550 23998 93602
rect 24050 93550 24062 93602
rect 9662 93538 9714 93550
rect 20078 93538 20130 93550
rect 24558 93538 24610 93550
rect 2046 93490 2098 93502
rect 19518 93490 19570 93502
rect 12338 93438 12350 93490
rect 12402 93438 12414 93490
rect 2046 93426 2098 93438
rect 19518 93426 19570 93438
rect 27358 93490 27410 93502
rect 27358 93426 27410 93438
rect 30830 93490 30882 93502
rect 30830 93426 30882 93438
rect 35198 93490 35250 93502
rect 35198 93426 35250 93438
rect 1344 93322 38640 93356
rect 1344 93270 4478 93322
rect 4530 93270 4582 93322
rect 4634 93270 4686 93322
rect 4738 93270 35198 93322
rect 35250 93270 35302 93322
rect 35354 93270 35406 93322
rect 35458 93270 38640 93322
rect 1344 93236 38640 93270
rect 4958 93154 5010 93166
rect 4958 93090 5010 93102
rect 10782 93154 10834 93166
rect 10782 93090 10834 93102
rect 19294 93154 19346 93166
rect 19294 93090 19346 93102
rect 23438 93154 23490 93166
rect 24446 93154 24498 93166
rect 24098 93102 24110 93154
rect 24162 93102 24174 93154
rect 23438 93090 23490 93102
rect 24446 93090 24498 93102
rect 25678 93154 25730 93166
rect 25678 93090 25730 93102
rect 5742 93042 5794 93054
rect 5742 92978 5794 92990
rect 9326 93042 9378 93054
rect 18622 93042 18674 93054
rect 17266 92990 17278 93042
rect 17330 92990 17342 93042
rect 9326 92978 9378 92990
rect 18622 92978 18674 92990
rect 20750 93042 20802 93054
rect 20750 92978 20802 92990
rect 31502 93042 31554 93054
rect 31502 92978 31554 92990
rect 6974 92930 7026 92942
rect 12910 92930 12962 92942
rect 2930 92878 2942 92930
rect 2994 92878 3006 92930
rect 3826 92878 3838 92930
rect 3890 92878 3902 92930
rect 7746 92878 7758 92930
rect 7810 92878 7822 92930
rect 12114 92878 12126 92930
rect 12178 92878 12190 92930
rect 6974 92866 7026 92878
rect 12910 92866 12962 92878
rect 17054 92930 17106 92942
rect 21310 92930 21362 92942
rect 24670 92930 24722 92942
rect 17938 92878 17950 92930
rect 18002 92878 18014 92930
rect 22306 92878 22318 92930
rect 22370 92878 22382 92930
rect 29250 92878 29262 92930
rect 29314 92878 29326 92930
rect 30146 92878 30158 92930
rect 30210 92878 30222 92930
rect 31826 92878 31838 92930
rect 31890 92878 31902 92930
rect 32722 92878 32734 92930
rect 32786 92878 32798 92930
rect 17054 92866 17106 92878
rect 21310 92866 21362 92878
rect 24670 92866 24722 92878
rect 9662 92818 9714 92830
rect 9662 92754 9714 92766
rect 10334 92818 10386 92830
rect 10334 92754 10386 92766
rect 13470 92818 13522 92830
rect 13470 92754 13522 92766
rect 13806 92818 13858 92830
rect 13806 92754 13858 92766
rect 14142 92818 14194 92830
rect 14142 92754 14194 92766
rect 14590 92818 14642 92830
rect 14590 92754 14642 92766
rect 19406 92818 19458 92830
rect 19406 92754 19458 92766
rect 25566 92818 25618 92830
rect 26674 92766 26686 92818
rect 26738 92766 26750 92818
rect 27458 92766 27470 92818
rect 27522 92766 27534 92818
rect 25566 92754 25618 92766
rect 25118 92706 25170 92718
rect 25118 92642 25170 92654
rect 26126 92706 26178 92718
rect 26126 92642 26178 92654
rect 34078 92706 34130 92718
rect 34078 92642 34130 92654
rect 1344 92538 38640 92572
rect 1344 92486 19838 92538
rect 19890 92486 19942 92538
rect 19994 92486 20046 92538
rect 20098 92486 38640 92538
rect 1344 92452 38640 92486
rect 5630 92370 5682 92382
rect 5630 92306 5682 92318
rect 8766 92370 8818 92382
rect 23214 92370 23266 92382
rect 10770 92318 10782 92370
rect 10834 92318 10846 92370
rect 8766 92306 8818 92318
rect 23214 92306 23266 92318
rect 9998 92258 10050 92270
rect 4834 92206 4846 92258
rect 4898 92206 4910 92258
rect 9998 92194 10050 92206
rect 10222 92258 10274 92270
rect 10222 92194 10274 92206
rect 13470 92258 13522 92270
rect 13470 92194 13522 92206
rect 14702 92258 14754 92270
rect 14702 92194 14754 92206
rect 15150 92258 15202 92270
rect 15150 92194 15202 92206
rect 20750 92258 20802 92270
rect 37886 92258 37938 92270
rect 26114 92206 26126 92258
rect 26178 92206 26190 92258
rect 20750 92194 20802 92206
rect 37886 92194 37938 92206
rect 12350 92146 12402 92158
rect 14366 92146 14418 92158
rect 2930 92094 2942 92146
rect 2994 92094 3006 92146
rect 3826 92094 3838 92146
rect 3890 92094 3902 92146
rect 6514 92094 6526 92146
rect 6578 92094 6590 92146
rect 7298 92094 7310 92146
rect 7362 92094 7374 92146
rect 10882 92094 10894 92146
rect 10946 92094 10958 92146
rect 12674 92094 12686 92146
rect 12738 92094 12750 92146
rect 12350 92082 12402 92094
rect 14366 92082 14418 92094
rect 20974 92146 21026 92158
rect 25342 92146 25394 92158
rect 38222 92146 38274 92158
rect 21634 92094 21646 92146
rect 21698 92094 21710 92146
rect 27346 92094 27358 92146
rect 27410 92094 27422 92146
rect 33170 92094 33182 92146
rect 33234 92094 33246 92146
rect 33842 92094 33854 92146
rect 33906 92094 33918 92146
rect 20974 92082 21026 92094
rect 25342 92082 25394 92094
rect 38222 92082 38274 92094
rect 22318 92034 22370 92046
rect 22318 91970 22370 91982
rect 23326 92034 23378 92046
rect 23326 91970 23378 91982
rect 24222 92034 24274 92046
rect 24222 91970 24274 91982
rect 24670 92034 24722 92046
rect 37662 92034 37714 92046
rect 26114 91982 26126 92034
rect 26178 91982 26190 92034
rect 27794 91982 27806 92034
rect 27858 91982 27870 92034
rect 24670 91970 24722 91982
rect 37662 91970 37714 91982
rect 10334 91922 10386 91934
rect 10334 91858 10386 91870
rect 14590 91922 14642 91934
rect 14590 91858 14642 91870
rect 35198 91922 35250 91934
rect 35198 91858 35250 91870
rect 1344 91754 38640 91788
rect 1344 91702 4478 91754
rect 4530 91702 4582 91754
rect 4634 91702 4686 91754
rect 4738 91702 35198 91754
rect 35250 91702 35302 91754
rect 35354 91702 35406 91754
rect 35458 91702 38640 91754
rect 1344 91668 38640 91702
rect 4958 91586 5010 91598
rect 4958 91522 5010 91534
rect 12238 91586 12290 91598
rect 32510 91586 32562 91598
rect 12562 91534 12574 91586
rect 12626 91534 12638 91586
rect 14018 91534 14030 91586
rect 14082 91583 14094 91586
rect 14578 91583 14590 91586
rect 14082 91537 14590 91583
rect 14082 91534 14094 91537
rect 14578 91534 14590 91537
rect 14642 91534 14654 91586
rect 12238 91522 12290 91534
rect 32510 91522 32562 91534
rect 8878 91474 8930 91486
rect 8878 91410 8930 91422
rect 14254 91474 14306 91486
rect 14254 91410 14306 91422
rect 14702 91474 14754 91486
rect 14702 91410 14754 91422
rect 11566 91362 11618 91374
rect 2930 91310 2942 91362
rect 2994 91310 3006 91362
rect 3826 91310 3838 91362
rect 3890 91310 3902 91362
rect 11566 91298 11618 91310
rect 12014 91362 12066 91374
rect 12014 91298 12066 91310
rect 13582 91362 13634 91374
rect 13794 91310 13806 91362
rect 13858 91310 13870 91362
rect 27682 91310 27694 91362
rect 27746 91310 27758 91362
rect 33842 91310 33854 91362
rect 33906 91310 33918 91362
rect 34514 91310 34526 91362
rect 34578 91310 34590 91362
rect 13582 91298 13634 91310
rect 13470 91250 13522 91262
rect 23762 91198 23774 91250
rect 23826 91198 23838 91250
rect 13470 91186 13522 91198
rect 5742 91138 5794 91150
rect 5742 91074 5794 91086
rect 11678 91138 11730 91150
rect 11678 91074 11730 91086
rect 1344 90970 38640 91004
rect 1344 90918 19838 90970
rect 19890 90918 19942 90970
rect 19994 90918 20046 90970
rect 20098 90918 38640 90970
rect 1344 90884 38640 90918
rect 12574 90802 12626 90814
rect 12574 90738 12626 90750
rect 24110 90690 24162 90702
rect 29710 90690 29762 90702
rect 26002 90638 26014 90690
rect 26066 90638 26078 90690
rect 24110 90626 24162 90638
rect 29710 90626 29762 90638
rect 30158 90690 30210 90702
rect 30158 90626 30210 90638
rect 22990 90578 23042 90590
rect 3154 90526 3166 90578
rect 3218 90526 3230 90578
rect 3826 90526 3838 90578
rect 3890 90526 3902 90578
rect 12338 90526 12350 90578
rect 12402 90526 12414 90578
rect 22990 90514 23042 90526
rect 25678 90578 25730 90590
rect 25678 90514 25730 90526
rect 30270 90578 30322 90590
rect 30270 90514 30322 90526
rect 5742 90466 5794 90478
rect 5742 90402 5794 90414
rect 21758 90466 21810 90478
rect 21758 90402 21810 90414
rect 22206 90466 22258 90478
rect 22206 90402 22258 90414
rect 22654 90466 22706 90478
rect 22654 90402 22706 90414
rect 23550 90466 23602 90478
rect 23550 90402 23602 90414
rect 24782 90466 24834 90478
rect 24782 90402 24834 90414
rect 25454 90466 25506 90478
rect 25454 90402 25506 90414
rect 26574 90466 26626 90478
rect 26574 90402 26626 90414
rect 27022 90466 27074 90478
rect 27022 90402 27074 90414
rect 27470 90466 27522 90478
rect 27470 90402 27522 90414
rect 27918 90466 27970 90478
rect 27918 90402 27970 90414
rect 28254 90466 28306 90478
rect 28254 90402 28306 90414
rect 5182 90354 5234 90366
rect 5182 90290 5234 90302
rect 12686 90354 12738 90366
rect 30158 90354 30210 90366
rect 26226 90302 26238 90354
rect 26290 90351 26302 90354
rect 26562 90351 26574 90354
rect 26290 90305 26574 90351
rect 26290 90302 26302 90305
rect 26562 90302 26574 90305
rect 26626 90302 26638 90354
rect 12686 90290 12738 90302
rect 30158 90290 30210 90302
rect 1344 90186 38640 90220
rect 1344 90134 4478 90186
rect 4530 90134 4582 90186
rect 4634 90134 4686 90186
rect 4738 90134 35198 90186
rect 35250 90134 35302 90186
rect 35354 90134 35406 90186
rect 35458 90134 38640 90186
rect 1344 90100 38640 90134
rect 30258 89966 30270 90018
rect 30322 89966 30334 90018
rect 10782 89906 10834 89918
rect 10782 89842 10834 89854
rect 21646 89906 21698 89918
rect 27346 89854 27358 89906
rect 27410 89854 27422 89906
rect 30482 89854 30494 89906
rect 30546 89854 30558 89906
rect 21646 89842 21698 89854
rect 8430 89794 8482 89806
rect 19966 89794 20018 89806
rect 3378 89742 3390 89794
rect 3442 89742 3454 89794
rect 4274 89742 4286 89794
rect 4338 89742 4350 89794
rect 7298 89742 7310 89794
rect 7362 89742 7374 89794
rect 7970 89742 7982 89794
rect 8034 89742 8046 89794
rect 9314 89742 9326 89794
rect 9378 89742 9390 89794
rect 8430 89730 8482 89742
rect 19966 89730 20018 89742
rect 22766 89794 22818 89806
rect 27010 89742 27022 89794
rect 27074 89742 27086 89794
rect 30370 89742 30382 89794
rect 30434 89742 30446 89794
rect 22766 89730 22818 89742
rect 22094 89682 22146 89694
rect 22094 89618 22146 89630
rect 23886 89682 23938 89694
rect 23886 89618 23938 89630
rect 26574 89682 26626 89694
rect 26574 89618 26626 89630
rect 2046 89570 2098 89582
rect 2046 89506 2098 89518
rect 4846 89570 4898 89582
rect 4846 89506 4898 89518
rect 5742 89570 5794 89582
rect 5742 89506 5794 89518
rect 15934 89570 15986 89582
rect 15934 89506 15986 89518
rect 16494 89570 16546 89582
rect 16494 89506 16546 89518
rect 17278 89570 17330 89582
rect 17278 89506 17330 89518
rect 19518 89570 19570 89582
rect 19518 89506 19570 89518
rect 22542 89570 22594 89582
rect 22542 89506 22594 89518
rect 22654 89570 22706 89582
rect 22654 89506 22706 89518
rect 22990 89570 23042 89582
rect 22990 89506 23042 89518
rect 23326 89570 23378 89582
rect 23326 89506 23378 89518
rect 23438 89570 23490 89582
rect 23438 89506 23490 89518
rect 23662 89570 23714 89582
rect 23662 89506 23714 89518
rect 24222 89570 24274 89582
rect 25118 89570 25170 89582
rect 24546 89518 24558 89570
rect 24610 89518 24622 89570
rect 24222 89506 24274 89518
rect 25118 89506 25170 89518
rect 25790 89570 25842 89582
rect 25790 89506 25842 89518
rect 26014 89570 26066 89582
rect 26014 89506 26066 89518
rect 26126 89570 26178 89582
rect 26126 89506 26178 89518
rect 26238 89570 26290 89582
rect 26238 89506 26290 89518
rect 28030 89570 28082 89582
rect 28030 89506 28082 89518
rect 28478 89570 28530 89582
rect 28478 89506 28530 89518
rect 29262 89570 29314 89582
rect 29262 89506 29314 89518
rect 1344 89402 38640 89436
rect 1344 89350 19838 89402
rect 19890 89350 19942 89402
rect 19994 89350 20046 89402
rect 20098 89350 38640 89402
rect 1344 89316 38640 89350
rect 24670 89234 24722 89246
rect 24670 89170 24722 89182
rect 16718 89122 16770 89134
rect 16718 89058 16770 89070
rect 12910 89010 12962 89022
rect 16830 89010 16882 89022
rect 20750 89010 20802 89022
rect 23998 89010 24050 89022
rect 6850 88958 6862 89010
rect 6914 88958 6926 89010
rect 7522 88958 7534 89010
rect 7586 88958 7598 89010
rect 13346 88958 13358 89010
rect 13410 88958 13422 89010
rect 17490 88958 17502 89010
rect 17554 88958 17566 89010
rect 21970 88958 21982 89010
rect 22034 88958 22046 89010
rect 23538 88958 23550 89010
rect 23602 88958 23614 89010
rect 12910 88946 12962 88958
rect 16830 88946 16882 88958
rect 20750 88946 20802 88958
rect 23998 88946 24050 88958
rect 24446 89010 24498 89022
rect 25218 88958 25230 89010
rect 25282 88958 25294 89010
rect 37874 88958 37886 89010
rect 37938 88958 37950 89010
rect 24446 88946 24498 88958
rect 9102 88898 9154 88910
rect 22766 88898 22818 88910
rect 14018 88846 14030 88898
rect 14082 88846 14094 88898
rect 16146 88846 16158 88898
rect 16210 88846 16222 88898
rect 18274 88846 18286 88898
rect 18338 88846 18350 88898
rect 20402 88846 20414 88898
rect 20466 88846 20478 88898
rect 21186 88846 21198 88898
rect 21250 88846 21262 88898
rect 9102 88834 9154 88846
rect 22766 88834 22818 88846
rect 24558 88898 24610 88910
rect 31054 88898 31106 88910
rect 30146 88846 30158 88898
rect 30210 88846 30222 88898
rect 36530 88846 36542 88898
rect 36594 88846 36606 88898
rect 24558 88834 24610 88846
rect 31054 88834 31106 88846
rect 16718 88786 16770 88798
rect 16718 88722 16770 88734
rect 1344 88618 38640 88652
rect 1344 88566 4478 88618
rect 4530 88566 4582 88618
rect 4634 88566 4686 88618
rect 4738 88566 35198 88618
rect 35250 88566 35302 88618
rect 35354 88566 35406 88618
rect 35458 88566 38640 88618
rect 1344 88532 38640 88566
rect 2158 88450 2210 88462
rect 2158 88386 2210 88398
rect 21758 88450 21810 88462
rect 22082 88398 22094 88450
rect 22146 88398 22158 88450
rect 24994 88398 25006 88450
rect 25058 88398 25070 88450
rect 21758 88386 21810 88398
rect 12798 88338 12850 88350
rect 15474 88286 15486 88338
rect 15538 88286 15550 88338
rect 16930 88286 16942 88338
rect 16994 88286 17006 88338
rect 24882 88286 24894 88338
rect 24946 88286 24958 88338
rect 29922 88286 29934 88338
rect 29986 88286 29998 88338
rect 32050 88286 32062 88338
rect 32114 88286 32126 88338
rect 12798 88274 12850 88286
rect 4286 88226 4338 88238
rect 3266 88174 3278 88226
rect 3330 88174 3342 88226
rect 4286 88162 4338 88174
rect 7086 88226 7138 88238
rect 9662 88226 9714 88238
rect 12574 88226 12626 88238
rect 7858 88174 7870 88226
rect 7922 88174 7934 88226
rect 10546 88174 10558 88226
rect 10610 88174 10622 88226
rect 7086 88162 7138 88174
rect 9662 88162 9714 88174
rect 12574 88162 12626 88174
rect 14030 88226 14082 88238
rect 19518 88226 19570 88238
rect 15250 88174 15262 88226
rect 15314 88174 15326 88226
rect 16146 88174 16158 88226
rect 16210 88174 16222 88226
rect 14030 88162 14082 88174
rect 19518 88162 19570 88174
rect 19854 88226 19906 88238
rect 19854 88162 19906 88174
rect 20638 88226 20690 88238
rect 20638 88162 20690 88174
rect 21534 88226 21586 88238
rect 22418 88174 22430 88226
rect 22482 88174 22494 88226
rect 24770 88174 24782 88226
rect 24834 88174 24846 88226
rect 28578 88174 28590 88226
rect 28642 88174 28654 88226
rect 29250 88174 29262 88226
rect 29314 88174 29326 88226
rect 21534 88162 21586 88174
rect 14366 88114 14418 88126
rect 14366 88050 14418 88062
rect 14702 88114 14754 88126
rect 35646 88114 35698 88126
rect 27794 88062 27806 88114
rect 27858 88062 27870 88114
rect 14702 88050 14754 88062
rect 35646 88050 35698 88062
rect 4734 88002 4786 88014
rect 4734 87938 4786 87950
rect 9438 88002 9490 88014
rect 9438 87938 9490 87950
rect 12014 88002 12066 88014
rect 13806 88002 13858 88014
rect 12226 87950 12238 88002
rect 12290 87950 12302 88002
rect 12014 87938 12066 87950
rect 13806 87938 13858 87950
rect 14254 88002 14306 88014
rect 19742 88002 19794 88014
rect 19170 87950 19182 88002
rect 19234 87950 19246 88002
rect 14254 87938 14306 87950
rect 19742 87938 19794 87950
rect 20302 88002 20354 88014
rect 20302 87938 20354 87950
rect 20750 88002 20802 88014
rect 32510 88002 32562 88014
rect 25554 87950 25566 88002
rect 25618 87950 25630 88002
rect 20750 87938 20802 87950
rect 32510 87938 32562 87950
rect 35086 88002 35138 88014
rect 35086 87938 35138 87950
rect 35310 88002 35362 88014
rect 35310 87938 35362 87950
rect 35534 88002 35586 88014
rect 35534 87938 35586 87950
rect 1344 87834 38640 87868
rect 1344 87782 19838 87834
rect 19890 87782 19942 87834
rect 19994 87782 20046 87834
rect 20098 87782 38640 87834
rect 1344 87748 38640 87782
rect 9102 87666 9154 87678
rect 9102 87602 9154 87614
rect 11902 87666 11954 87678
rect 11902 87602 11954 87614
rect 14366 87666 14418 87678
rect 14366 87602 14418 87614
rect 15262 87666 15314 87678
rect 15262 87602 15314 87614
rect 15710 87666 15762 87678
rect 15710 87602 15762 87614
rect 17502 87666 17554 87678
rect 17502 87602 17554 87614
rect 20078 87666 20130 87678
rect 20078 87602 20130 87614
rect 22766 87666 22818 87678
rect 22766 87602 22818 87614
rect 22990 87666 23042 87678
rect 22990 87602 23042 87614
rect 23214 87666 23266 87678
rect 23214 87602 23266 87614
rect 23550 87666 23602 87678
rect 23550 87602 23602 87614
rect 23774 87666 23826 87678
rect 23774 87602 23826 87614
rect 16718 87554 16770 87566
rect 19070 87554 19122 87566
rect 24334 87554 24386 87566
rect 13570 87502 13582 87554
rect 13634 87502 13646 87554
rect 18162 87502 18174 87554
rect 18226 87502 18238 87554
rect 18722 87502 18734 87554
rect 18786 87502 18798 87554
rect 21074 87502 21086 87554
rect 21138 87502 21150 87554
rect 16718 87490 16770 87502
rect 19070 87490 19122 87502
rect 24334 87490 24386 87502
rect 24558 87554 24610 87566
rect 31166 87554 31218 87566
rect 27234 87502 27246 87554
rect 27298 87502 27310 87554
rect 35634 87502 35646 87554
rect 35698 87502 35710 87554
rect 24558 87490 24610 87502
rect 31166 87490 31218 87502
rect 4286 87442 4338 87454
rect 12350 87442 12402 87454
rect 13918 87442 13970 87454
rect 3266 87390 3278 87442
rect 3330 87390 3342 87442
rect 6850 87390 6862 87442
rect 6914 87390 6926 87442
rect 7746 87390 7758 87442
rect 7810 87390 7822 87442
rect 9650 87390 9662 87442
rect 9714 87390 9726 87442
rect 10546 87390 10558 87442
rect 10610 87390 10622 87442
rect 13010 87390 13022 87442
rect 13074 87390 13086 87442
rect 4286 87378 4338 87390
rect 12350 87378 12402 87390
rect 13918 87378 13970 87390
rect 15598 87442 15650 87454
rect 19630 87442 19682 87454
rect 16258 87390 16270 87442
rect 16322 87390 16334 87442
rect 17826 87390 17838 87442
rect 17890 87390 17902 87442
rect 15598 87378 15650 87390
rect 19630 87378 19682 87390
rect 20638 87442 20690 87454
rect 24222 87442 24274 87454
rect 20962 87390 20974 87442
rect 21026 87390 21038 87442
rect 21186 87390 21198 87442
rect 21250 87390 21262 87442
rect 22194 87390 22206 87442
rect 22258 87390 22270 87442
rect 20638 87378 20690 87390
rect 24222 87378 24274 87390
rect 24670 87442 24722 87454
rect 31054 87442 31106 87454
rect 25666 87390 25678 87442
rect 25730 87390 25742 87442
rect 30818 87390 30830 87442
rect 30882 87390 30894 87442
rect 24670 87378 24722 87390
rect 31054 87378 31106 87390
rect 32062 87442 32114 87454
rect 32062 87378 32114 87390
rect 32958 87442 33010 87454
rect 32958 87378 33010 87390
rect 33406 87442 33458 87454
rect 33406 87378 33458 87390
rect 33630 87442 33682 87454
rect 33630 87378 33682 87390
rect 34526 87442 34578 87454
rect 34850 87390 34862 87442
rect 34914 87390 34926 87442
rect 34526 87378 34578 87390
rect 4734 87330 4786 87342
rect 4734 87266 4786 87278
rect 5182 87330 5234 87342
rect 5182 87266 5234 87278
rect 23102 87330 23154 87342
rect 23102 87266 23154 87278
rect 23662 87330 23714 87342
rect 23662 87266 23714 87278
rect 32510 87330 32562 87342
rect 32510 87266 32562 87278
rect 33518 87330 33570 87342
rect 37762 87278 37774 87330
rect 37826 87278 37838 87330
rect 33518 87266 33570 87278
rect 2158 87218 2210 87230
rect 15710 87218 15762 87230
rect 12562 87166 12574 87218
rect 12626 87166 12638 87218
rect 31602 87166 31614 87218
rect 31666 87166 31678 87218
rect 2158 87154 2210 87166
rect 15710 87154 15762 87166
rect 1344 87050 38640 87084
rect 1344 86998 4478 87050
rect 4530 86998 4582 87050
rect 4634 86998 4686 87050
rect 4738 86998 35198 87050
rect 35250 86998 35302 87050
rect 35354 86998 35406 87050
rect 35458 86998 38640 87050
rect 1344 86964 38640 86998
rect 2158 86882 2210 86894
rect 2158 86818 2210 86830
rect 24670 86882 24722 86894
rect 26002 86830 26014 86882
rect 26066 86830 26078 86882
rect 24670 86818 24722 86830
rect 16046 86770 16098 86782
rect 16046 86706 16098 86718
rect 16830 86770 16882 86782
rect 16830 86706 16882 86718
rect 18286 86770 18338 86782
rect 18286 86706 18338 86718
rect 19182 86770 19234 86782
rect 19182 86706 19234 86718
rect 19854 86770 19906 86782
rect 29150 86770 29202 86782
rect 36206 86770 36258 86782
rect 22082 86718 22094 86770
rect 22146 86718 22158 86770
rect 22306 86718 22318 86770
rect 22370 86718 22382 86770
rect 26114 86718 26126 86770
rect 26178 86718 26190 86770
rect 29586 86718 29598 86770
rect 29650 86718 29662 86770
rect 32834 86718 32846 86770
rect 32898 86718 32910 86770
rect 34962 86718 34974 86770
rect 35026 86718 35038 86770
rect 19854 86706 19906 86718
rect 29150 86706 29202 86718
rect 36206 86706 36258 86718
rect 4286 86658 4338 86670
rect 9326 86658 9378 86670
rect 3266 86606 3278 86658
rect 3330 86606 3342 86658
rect 8418 86606 8430 86658
rect 8482 86606 8494 86658
rect 4286 86594 4338 86606
rect 9326 86594 9378 86606
rect 10110 86658 10162 86670
rect 10110 86594 10162 86606
rect 10670 86658 10722 86670
rect 16942 86658 16994 86670
rect 20302 86658 20354 86670
rect 11666 86606 11678 86658
rect 11730 86606 11742 86658
rect 17490 86606 17502 86658
rect 17554 86606 17566 86658
rect 10670 86594 10722 86606
rect 16942 86594 16994 86606
rect 20302 86594 20354 86606
rect 20750 86658 20802 86670
rect 23214 86658 23266 86670
rect 21970 86606 21982 86658
rect 22034 86606 22046 86658
rect 22754 86606 22766 86658
rect 22818 86606 22830 86658
rect 20750 86594 20802 86606
rect 23214 86594 23266 86606
rect 23550 86658 23602 86670
rect 23550 86594 23602 86606
rect 24334 86658 24386 86670
rect 27134 86658 27186 86670
rect 25106 86606 25118 86658
rect 25170 86606 25182 86658
rect 25890 86606 25902 86658
rect 25954 86606 25966 86658
rect 24334 86594 24386 86606
rect 27134 86594 27186 86606
rect 28030 86658 28082 86670
rect 28030 86594 28082 86606
rect 28478 86658 28530 86670
rect 32498 86606 32510 86658
rect 32562 86606 32574 86658
rect 35634 86606 35646 86658
rect 35698 86606 35710 86658
rect 28478 86594 28530 86606
rect 10894 86546 10946 86558
rect 20414 86546 20466 86558
rect 12562 86494 12574 86546
rect 12626 86494 12638 86546
rect 10894 86482 10946 86494
rect 20414 86482 20466 86494
rect 23774 86546 23826 86558
rect 23774 86482 23826 86494
rect 24110 86546 24162 86558
rect 24110 86482 24162 86494
rect 26910 86546 26962 86558
rect 31714 86494 31726 86546
rect 31778 86494 31790 86546
rect 26910 86482 26962 86494
rect 4734 86434 4786 86446
rect 4734 86370 4786 86382
rect 6974 86434 7026 86446
rect 6974 86370 7026 86382
rect 20638 86434 20690 86446
rect 20638 86370 20690 86382
rect 23662 86434 23714 86446
rect 23662 86370 23714 86382
rect 27022 86434 27074 86446
rect 27022 86370 27074 86382
rect 27358 86434 27410 86446
rect 27358 86370 27410 86382
rect 27806 86434 27858 86446
rect 27806 86370 27858 86382
rect 27918 86434 27970 86446
rect 27918 86370 27970 86382
rect 29262 86434 29314 86446
rect 29262 86370 29314 86382
rect 1344 86266 38640 86300
rect 1344 86214 19838 86266
rect 19890 86214 19942 86266
rect 19994 86214 20046 86266
rect 20098 86214 38640 86266
rect 1344 86180 38640 86214
rect 7310 86098 7362 86110
rect 7310 86034 7362 86046
rect 11678 86098 11730 86110
rect 11678 86034 11730 86046
rect 12126 86098 12178 86110
rect 12126 86034 12178 86046
rect 31502 86098 31554 86110
rect 31502 86034 31554 86046
rect 36318 86098 36370 86110
rect 36318 86034 36370 86046
rect 11566 85986 11618 85998
rect 11566 85922 11618 85934
rect 25342 85986 25394 85998
rect 31614 85986 31666 85998
rect 27458 85934 27470 85986
rect 27522 85934 27534 85986
rect 25342 85922 25394 85934
rect 31614 85922 31666 85934
rect 4286 85874 4338 85886
rect 3266 85822 3278 85874
rect 3330 85822 3342 85874
rect 4286 85810 4338 85822
rect 4622 85874 4674 85886
rect 6974 85874 7026 85886
rect 25230 85874 25282 85886
rect 31166 85874 31218 85886
rect 5394 85822 5406 85874
rect 5458 85822 5470 85874
rect 14130 85822 14142 85874
rect 14194 85822 14206 85874
rect 23538 85822 23550 85874
rect 23602 85822 23614 85874
rect 30258 85822 30270 85874
rect 30322 85822 30334 85874
rect 4622 85810 4674 85822
rect 6974 85810 7026 85822
rect 25230 85810 25282 85822
rect 31166 85810 31218 85822
rect 31838 85874 31890 85886
rect 36206 85874 36258 85886
rect 33618 85822 33630 85874
rect 33682 85822 33694 85874
rect 34962 85822 34974 85874
rect 35026 85822 35038 85874
rect 31838 85810 31890 85822
rect 36206 85810 36258 85822
rect 13806 85762 13858 85774
rect 32510 85762 32562 85774
rect 14242 85710 14254 85762
rect 14306 85710 14318 85762
rect 19618 85710 19630 85762
rect 19682 85710 19694 85762
rect 13806 85698 13858 85710
rect 32510 85698 32562 85710
rect 33070 85762 33122 85774
rect 35758 85762 35810 85774
rect 35074 85710 35086 85762
rect 35138 85710 35150 85762
rect 33070 85698 33122 85710
rect 35758 85698 35810 85710
rect 36878 85762 36930 85774
rect 36878 85698 36930 85710
rect 37326 85762 37378 85774
rect 37326 85698 37378 85710
rect 2158 85650 2210 85662
rect 2158 85586 2210 85598
rect 14478 85650 14530 85662
rect 14478 85586 14530 85598
rect 33294 85650 33346 85662
rect 33294 85586 33346 85598
rect 36318 85650 36370 85662
rect 36318 85586 36370 85598
rect 1344 85482 38640 85516
rect 1344 85430 4478 85482
rect 4530 85430 4582 85482
rect 4634 85430 4686 85482
rect 4738 85430 35198 85482
rect 35250 85430 35302 85482
rect 35354 85430 35406 85482
rect 35458 85430 38640 85482
rect 1344 85396 38640 85430
rect 2158 85314 2210 85326
rect 2158 85250 2210 85262
rect 14814 85314 14866 85326
rect 20414 85314 20466 85326
rect 15138 85262 15150 85314
rect 15202 85262 15214 85314
rect 19058 85262 19070 85314
rect 19122 85311 19134 85314
rect 19618 85311 19630 85314
rect 19122 85265 19630 85311
rect 19122 85262 19134 85265
rect 19618 85262 19630 85265
rect 19682 85262 19694 85314
rect 14814 85250 14866 85262
rect 20414 85250 20466 85262
rect 21758 85314 21810 85326
rect 21758 85250 21810 85262
rect 32510 85314 32562 85326
rect 32510 85250 32562 85262
rect 32846 85314 32898 85326
rect 32846 85250 32898 85262
rect 29934 85202 29986 85214
rect 29474 85150 29486 85202
rect 29538 85150 29550 85202
rect 29934 85138 29986 85150
rect 30830 85202 30882 85214
rect 30830 85138 30882 85150
rect 31726 85202 31778 85214
rect 31726 85138 31778 85150
rect 37102 85202 37154 85214
rect 37102 85138 37154 85150
rect 4286 85090 4338 85102
rect 3266 85038 3278 85090
rect 3330 85038 3342 85090
rect 4286 85026 4338 85038
rect 14030 85090 14082 85102
rect 14030 85026 14082 85038
rect 14254 85090 14306 85102
rect 14254 85026 14306 85038
rect 14590 85090 14642 85102
rect 14590 85026 14642 85038
rect 15598 85090 15650 85102
rect 15598 85026 15650 85038
rect 19182 85090 19234 85102
rect 19182 85026 19234 85038
rect 20526 85090 20578 85102
rect 21422 85090 21474 85102
rect 20738 85038 20750 85090
rect 20802 85038 20814 85090
rect 20526 85026 20578 85038
rect 21422 85026 21474 85038
rect 21870 85090 21922 85102
rect 21870 85026 21922 85038
rect 22094 85090 22146 85102
rect 31278 85090 31330 85102
rect 22306 85038 22318 85090
rect 22370 85038 22382 85090
rect 22642 85038 22654 85090
rect 22706 85038 22718 85090
rect 29362 85038 29374 85090
rect 29426 85038 29438 85090
rect 22094 85026 22146 85038
rect 31278 85026 31330 85038
rect 31614 85090 31666 85102
rect 31614 85026 31666 85038
rect 31838 85090 31890 85102
rect 31838 85026 31890 85038
rect 34414 85090 34466 85102
rect 34414 85026 34466 85038
rect 35646 85090 35698 85102
rect 35646 85026 35698 85038
rect 35870 85090 35922 85102
rect 35870 85026 35922 85038
rect 32062 84978 32114 84990
rect 25554 84926 25566 84978
rect 25618 84926 25630 84978
rect 32062 84914 32114 84926
rect 34974 84978 35026 84990
rect 34974 84914 35026 84926
rect 35310 84978 35362 84990
rect 35310 84914 35362 84926
rect 35982 84978 36034 84990
rect 35982 84914 36034 84926
rect 4734 84866 4786 84878
rect 4734 84802 4786 84814
rect 12910 84866 12962 84878
rect 12910 84802 12962 84814
rect 13806 84866 13858 84878
rect 13806 84802 13858 84814
rect 14142 84866 14194 84878
rect 14142 84802 14194 84814
rect 18734 84866 18786 84878
rect 18734 84802 18786 84814
rect 19742 84866 19794 84878
rect 19742 84802 19794 84814
rect 20078 84866 20130 84878
rect 20078 84802 20130 84814
rect 28366 84866 28418 84878
rect 28366 84802 28418 84814
rect 30382 84866 30434 84878
rect 30382 84802 30434 84814
rect 32734 84866 32786 84878
rect 32734 84802 32786 84814
rect 33966 84866 34018 84878
rect 33966 84802 34018 84814
rect 34526 84866 34578 84878
rect 34526 84802 34578 84814
rect 34750 84866 34802 84878
rect 34750 84802 34802 84814
rect 35086 84866 35138 84878
rect 35086 84802 35138 84814
rect 35422 84866 35474 84878
rect 35422 84802 35474 84814
rect 36206 84866 36258 84878
rect 36206 84802 36258 84814
rect 37662 84866 37714 84878
rect 37662 84802 37714 84814
rect 1344 84698 38640 84732
rect 1344 84646 19838 84698
rect 19890 84646 19942 84698
rect 19994 84646 20046 84698
rect 20098 84646 38640 84698
rect 1344 84612 38640 84646
rect 17614 84530 17666 84542
rect 17614 84466 17666 84478
rect 18846 84530 18898 84542
rect 18846 84466 18898 84478
rect 19070 84530 19122 84542
rect 19070 84466 19122 84478
rect 21086 84530 21138 84542
rect 21086 84466 21138 84478
rect 21310 84530 21362 84542
rect 25678 84530 25730 84542
rect 23874 84478 23886 84530
rect 23938 84478 23950 84530
rect 21310 84466 21362 84478
rect 25678 84466 25730 84478
rect 25902 84530 25954 84542
rect 29150 84530 29202 84542
rect 28578 84478 28590 84530
rect 28642 84478 28654 84530
rect 25902 84466 25954 84478
rect 29150 84466 29202 84478
rect 30158 84530 30210 84542
rect 30158 84466 30210 84478
rect 30606 84530 30658 84542
rect 30606 84466 30658 84478
rect 31054 84530 31106 84542
rect 31054 84466 31106 84478
rect 34190 84530 34242 84542
rect 34190 84466 34242 84478
rect 34974 84530 35026 84542
rect 34974 84466 35026 84478
rect 19966 84418 20018 84430
rect 14690 84366 14702 84418
rect 14754 84366 14766 84418
rect 19966 84354 20018 84366
rect 20414 84418 20466 84430
rect 20414 84354 20466 84366
rect 23326 84418 23378 84430
rect 28030 84418 28082 84430
rect 24210 84366 24222 84418
rect 24274 84366 24286 84418
rect 23326 84354 23378 84366
rect 28030 84354 28082 84366
rect 29710 84418 29762 84430
rect 29710 84354 29762 84366
rect 4286 84306 4338 84318
rect 18510 84306 18562 84318
rect 3266 84254 3278 84306
rect 3330 84254 3342 84306
rect 15474 84254 15486 84306
rect 15538 84254 15550 84306
rect 4286 84242 4338 84254
rect 18510 84242 18562 84254
rect 19406 84306 19458 84318
rect 20638 84306 20690 84318
rect 23438 84306 23490 84318
rect 25230 84306 25282 84318
rect 20178 84254 20190 84306
rect 20242 84254 20254 84306
rect 22306 84254 22318 84306
rect 22370 84254 22382 84306
rect 22978 84254 22990 84306
rect 23042 84254 23054 84306
rect 24434 84254 24446 84306
rect 24498 84254 24510 84306
rect 26898 84254 26910 84306
rect 26962 84254 26974 84306
rect 27794 84254 27806 84306
rect 27858 84254 27870 84306
rect 35298 84254 35310 84306
rect 35362 84254 35374 84306
rect 19406 84242 19458 84254
rect 20638 84242 20690 84254
rect 23438 84242 23490 84254
rect 25230 84242 25282 84254
rect 4734 84194 4786 84206
rect 4734 84130 4786 84142
rect 8766 84194 8818 84206
rect 8766 84130 8818 84142
rect 12574 84194 12626 84206
rect 12574 84130 12626 84142
rect 15934 84194 15986 84206
rect 15934 84130 15986 84142
rect 18062 84194 18114 84206
rect 18062 84130 18114 84142
rect 21198 84194 21250 84206
rect 25454 84194 25506 84206
rect 22082 84142 22094 84194
rect 22146 84142 22158 84194
rect 22866 84142 22878 84194
rect 22930 84142 22942 84194
rect 21198 84130 21250 84142
rect 25454 84130 25506 84142
rect 25790 84194 25842 84206
rect 33854 84194 33906 84206
rect 27122 84142 27134 84194
rect 27186 84142 27198 84194
rect 27458 84142 27470 84194
rect 27522 84142 27534 84194
rect 36082 84142 36094 84194
rect 36146 84142 36158 84194
rect 38210 84142 38222 84194
rect 38274 84142 38286 84194
rect 25790 84130 25842 84142
rect 33854 84130 33906 84142
rect 2158 84082 2210 84094
rect 2158 84018 2210 84030
rect 18734 84082 18786 84094
rect 18734 84018 18786 84030
rect 19854 84082 19906 84094
rect 19854 84018 19906 84030
rect 28254 84082 28306 84094
rect 28254 84018 28306 84030
rect 1344 83914 38640 83948
rect 1344 83862 4478 83914
rect 4530 83862 4582 83914
rect 4634 83862 4686 83914
rect 4738 83862 35198 83914
rect 35250 83862 35302 83914
rect 35354 83862 35406 83914
rect 35458 83862 38640 83914
rect 1344 83828 38640 83862
rect 2158 83746 2210 83758
rect 29262 83746 29314 83758
rect 9090 83694 9102 83746
rect 9154 83743 9166 83746
rect 9762 83743 9774 83746
rect 9154 83697 9774 83743
rect 9154 83694 9166 83697
rect 9762 83694 9774 83697
rect 9826 83694 9838 83746
rect 14802 83694 14814 83746
rect 14866 83694 14878 83746
rect 2158 83682 2210 83694
rect 29262 83682 29314 83694
rect 37102 83746 37154 83758
rect 37102 83682 37154 83694
rect 9774 83634 9826 83646
rect 9774 83570 9826 83582
rect 16158 83634 16210 83646
rect 16158 83570 16210 83582
rect 17726 83634 17778 83646
rect 30494 83634 30546 83646
rect 19282 83582 19294 83634
rect 19346 83582 19358 83634
rect 20402 83582 20414 83634
rect 20466 83582 20478 83634
rect 17726 83570 17778 83582
rect 30494 83570 30546 83582
rect 34750 83634 34802 83646
rect 34750 83570 34802 83582
rect 37662 83634 37714 83646
rect 37662 83570 37714 83582
rect 38110 83634 38162 83646
rect 38110 83570 38162 83582
rect 4286 83522 4338 83534
rect 15374 83522 15426 83534
rect 3266 83470 3278 83522
rect 3330 83470 3342 83522
rect 8082 83470 8094 83522
rect 8146 83470 8158 83522
rect 4286 83458 4338 83470
rect 15374 83458 15426 83470
rect 17838 83522 17890 83534
rect 17838 83458 17890 83470
rect 18398 83522 18450 83534
rect 18398 83458 18450 83470
rect 18510 83522 18562 83534
rect 18510 83458 18562 83470
rect 19182 83522 19234 83534
rect 29038 83522 29090 83534
rect 19954 83470 19966 83522
rect 20018 83470 20030 83522
rect 21858 83470 21870 83522
rect 21922 83470 21934 83522
rect 24770 83470 24782 83522
rect 24834 83470 24846 83522
rect 19182 83458 19234 83470
rect 29038 83458 29090 83470
rect 34862 83522 34914 83534
rect 35634 83470 35646 83522
rect 35698 83470 35710 83522
rect 35970 83470 35982 83522
rect 36034 83470 36046 83522
rect 34862 83458 34914 83470
rect 4734 83410 4786 83422
rect 4734 83346 4786 83358
rect 8430 83410 8482 83422
rect 8430 83346 8482 83358
rect 14142 83410 14194 83422
rect 14142 83346 14194 83358
rect 14254 83410 14306 83422
rect 14254 83346 14306 83358
rect 14366 83410 14418 83422
rect 14366 83346 14418 83358
rect 15598 83410 15650 83422
rect 29598 83410 29650 83422
rect 22866 83358 22878 83410
rect 22930 83358 22942 83410
rect 26002 83358 26014 83410
rect 26066 83358 26078 83410
rect 15598 83346 15650 83358
rect 29598 83346 29650 83358
rect 31390 83410 31442 83422
rect 31390 83346 31442 83358
rect 36206 83410 36258 83422
rect 36206 83346 36258 83358
rect 36990 83410 37042 83422
rect 36990 83346 37042 83358
rect 37102 83410 37154 83422
rect 37102 83346 37154 83358
rect 8318 83298 8370 83310
rect 8318 83234 8370 83246
rect 9326 83298 9378 83310
rect 9326 83234 9378 83246
rect 13022 83298 13074 83310
rect 13022 83234 13074 83246
rect 13694 83298 13746 83310
rect 13694 83234 13746 83246
rect 15150 83298 15202 83310
rect 15150 83234 15202 83246
rect 15262 83298 15314 83310
rect 15262 83234 15314 83246
rect 16606 83298 16658 83310
rect 16606 83234 16658 83246
rect 17166 83298 17218 83310
rect 17166 83234 17218 83246
rect 18286 83298 18338 83310
rect 18286 83234 18338 83246
rect 19518 83298 19570 83310
rect 29374 83298 29426 83310
rect 22306 83246 22318 83298
rect 22370 83246 22382 83298
rect 19518 83234 19570 83246
rect 29374 83234 29426 83246
rect 30046 83298 30098 83310
rect 30046 83234 30098 83246
rect 30942 83298 30994 83310
rect 30942 83234 30994 83246
rect 34078 83298 34130 83310
rect 34078 83234 34130 83246
rect 34414 83298 34466 83310
rect 34414 83234 34466 83246
rect 34638 83298 34690 83310
rect 34638 83234 34690 83246
rect 37550 83298 37602 83310
rect 37550 83234 37602 83246
rect 1344 83130 38640 83164
rect 1344 83078 19838 83130
rect 19890 83078 19942 83130
rect 19994 83078 20046 83130
rect 20098 83078 38640 83130
rect 1344 83044 38640 83078
rect 17614 82962 17666 82974
rect 17614 82898 17666 82910
rect 28254 82962 28306 82974
rect 28254 82898 28306 82910
rect 29038 82962 29090 82974
rect 29038 82898 29090 82910
rect 30606 82962 30658 82974
rect 30606 82898 30658 82910
rect 10222 82850 10274 82862
rect 18622 82850 18674 82862
rect 28366 82850 28418 82862
rect 8194 82798 8206 82850
rect 8258 82798 8270 82850
rect 12674 82798 12686 82850
rect 12738 82798 12750 82850
rect 26450 82798 26462 82850
rect 26514 82798 26526 82850
rect 35746 82798 35758 82850
rect 35810 82798 35822 82850
rect 10222 82786 10274 82798
rect 18622 82786 18674 82798
rect 28366 82786 28418 82798
rect 9774 82738 9826 82750
rect 8978 82686 8990 82738
rect 9042 82686 9054 82738
rect 9538 82686 9550 82738
rect 9602 82686 9614 82738
rect 9774 82674 9826 82686
rect 9998 82738 10050 82750
rect 27246 82738 27298 82750
rect 12002 82686 12014 82738
rect 12066 82686 12078 82738
rect 19618 82686 19630 82738
rect 19682 82686 19694 82738
rect 25218 82686 25230 82738
rect 25282 82686 25294 82738
rect 25890 82686 25902 82738
rect 25954 82686 25966 82738
rect 9998 82674 10050 82686
rect 27246 82674 27298 82686
rect 27918 82738 27970 82750
rect 27918 82674 27970 82686
rect 28590 82738 28642 82750
rect 28590 82674 28642 82686
rect 28814 82738 28866 82750
rect 28814 82674 28866 82686
rect 29150 82738 29202 82750
rect 29150 82674 29202 82686
rect 29374 82738 29426 82750
rect 34962 82686 34974 82738
rect 35026 82686 35038 82738
rect 29374 82674 29426 82686
rect 10670 82626 10722 82638
rect 6066 82574 6078 82626
rect 6130 82574 6142 82626
rect 9650 82574 9662 82626
rect 9714 82574 9726 82626
rect 10670 82562 10722 82574
rect 11118 82626 11170 82638
rect 11118 82562 11170 82574
rect 14814 82626 14866 82638
rect 14814 82562 14866 82574
rect 15486 82626 15538 82638
rect 15486 82562 15538 82574
rect 18174 82626 18226 82638
rect 27134 82626 27186 82638
rect 23538 82574 23550 82626
rect 23602 82574 23614 82626
rect 26226 82574 26238 82626
rect 26290 82574 26302 82626
rect 18174 82562 18226 82574
rect 27134 82562 27186 82574
rect 29822 82626 29874 82638
rect 31166 82626 31218 82638
rect 30146 82574 30158 82626
rect 30210 82574 30222 82626
rect 29822 82562 29874 82574
rect 31166 82562 31218 82574
rect 31614 82626 31666 82638
rect 31614 82562 31666 82574
rect 33182 82626 33234 82638
rect 33182 82562 33234 82574
rect 34638 82626 34690 82638
rect 34638 82562 34690 82574
rect 37886 82626 37938 82638
rect 37886 82562 37938 82574
rect 18510 82514 18562 82526
rect 18510 82450 18562 82462
rect 18846 82514 18898 82526
rect 31390 82514 31442 82526
rect 27010 82462 27022 82514
rect 27074 82462 27086 82514
rect 18846 82450 18898 82462
rect 31390 82450 31442 82462
rect 31838 82514 31890 82526
rect 31838 82450 31890 82462
rect 32286 82514 32338 82526
rect 32286 82450 32338 82462
rect 1344 82346 38640 82380
rect 1344 82294 4478 82346
rect 4530 82294 4582 82346
rect 4634 82294 4686 82346
rect 4738 82294 35198 82346
rect 35250 82294 35302 82346
rect 35354 82294 35406 82346
rect 35458 82294 38640 82346
rect 1344 82260 38640 82294
rect 27358 82178 27410 82190
rect 14466 82126 14478 82178
rect 14530 82175 14542 82178
rect 14914 82175 14926 82178
rect 14530 82129 14926 82175
rect 14530 82126 14542 82129
rect 14914 82126 14926 82129
rect 14978 82175 14990 82178
rect 15362 82175 15374 82178
rect 14978 82129 15374 82175
rect 14978 82126 14990 82129
rect 15362 82126 15374 82129
rect 15426 82126 15438 82178
rect 27358 82114 27410 82126
rect 11566 82066 11618 82078
rect 11566 82002 11618 82014
rect 15262 82066 15314 82078
rect 20302 82066 20354 82078
rect 27022 82066 27074 82078
rect 18162 82014 18174 82066
rect 18226 82014 18238 82066
rect 23426 82014 23438 82066
rect 23490 82014 23502 82066
rect 15262 82002 15314 82014
rect 20302 82002 20354 82014
rect 27022 82002 27074 82014
rect 5182 81954 5234 81966
rect 5182 81890 5234 81902
rect 6302 81954 6354 81966
rect 6302 81890 6354 81902
rect 6638 81954 6690 81966
rect 13694 81954 13746 81966
rect 27918 81954 27970 81966
rect 10434 81902 10446 81954
rect 10498 81902 10510 81954
rect 17378 81902 17390 81954
rect 17442 81902 17454 81954
rect 25554 81902 25566 81954
rect 25618 81902 25630 81954
rect 27458 81902 27470 81954
rect 27522 81902 27534 81954
rect 6638 81890 6690 81902
rect 13694 81890 13746 81902
rect 27918 81890 27970 81902
rect 28366 81954 28418 81966
rect 28366 81890 28418 81902
rect 28590 81954 28642 81966
rect 28590 81890 28642 81902
rect 29934 81954 29986 81966
rect 32958 81954 33010 81966
rect 36206 81954 36258 81966
rect 30594 81902 30606 81954
rect 30658 81902 30670 81954
rect 31154 81902 31166 81954
rect 31218 81902 31230 81954
rect 35186 81902 35198 81954
rect 35250 81902 35262 81954
rect 29934 81890 29986 81902
rect 32958 81890 33010 81902
rect 36206 81890 36258 81902
rect 4846 81842 4898 81854
rect 4846 81778 4898 81790
rect 6078 81842 6130 81854
rect 10782 81842 10834 81854
rect 9650 81790 9662 81842
rect 9714 81790 9726 81842
rect 6078 81778 6130 81790
rect 10782 81778 10834 81790
rect 10894 81842 10946 81854
rect 10894 81778 10946 81790
rect 11006 81842 11058 81854
rect 11006 81778 11058 81790
rect 14142 81842 14194 81854
rect 14142 81778 14194 81790
rect 14366 81842 14418 81854
rect 14366 81778 14418 81790
rect 26910 81842 26962 81854
rect 32174 81842 32226 81854
rect 27122 81790 27134 81842
rect 27186 81790 27198 81842
rect 30706 81790 30718 81842
rect 30770 81790 30782 81842
rect 26910 81778 26962 81790
rect 32174 81778 32226 81790
rect 4622 81730 4674 81742
rect 4622 81666 4674 81678
rect 4958 81730 5010 81742
rect 4958 81666 5010 81678
rect 5854 81730 5906 81742
rect 5854 81666 5906 81678
rect 6414 81730 6466 81742
rect 13022 81730 13074 81742
rect 7410 81678 7422 81730
rect 7474 81678 7486 81730
rect 6414 81666 6466 81678
rect 13022 81666 13074 81678
rect 14030 81730 14082 81742
rect 14030 81666 14082 81678
rect 14814 81730 14866 81742
rect 14814 81666 14866 81678
rect 17054 81730 17106 81742
rect 17054 81666 17106 81678
rect 28142 81730 28194 81742
rect 28142 81666 28194 81678
rect 29598 81730 29650 81742
rect 29598 81666 29650 81678
rect 31278 81730 31330 81742
rect 31278 81666 31330 81678
rect 34190 81730 34242 81742
rect 34190 81666 34242 81678
rect 35310 81730 35362 81742
rect 35310 81666 35362 81678
rect 1344 81562 38640 81596
rect 1344 81510 19838 81562
rect 19890 81510 19942 81562
rect 19994 81510 20046 81562
rect 20098 81510 38640 81562
rect 1344 81476 38640 81510
rect 7086 81394 7138 81406
rect 7086 81330 7138 81342
rect 9886 81394 9938 81406
rect 9886 81330 9938 81342
rect 14478 81394 14530 81406
rect 14478 81330 14530 81342
rect 16942 81394 16994 81406
rect 16942 81330 16994 81342
rect 26574 81394 26626 81406
rect 26574 81330 26626 81342
rect 27806 81394 27858 81406
rect 27806 81330 27858 81342
rect 31614 81394 31666 81406
rect 31614 81330 31666 81342
rect 10222 81282 10274 81294
rect 20974 81282 21026 81294
rect 5842 81230 5854 81282
rect 5906 81230 5918 81282
rect 18162 81230 18174 81282
rect 18226 81230 18238 81282
rect 10222 81218 10274 81230
rect 20974 81218 21026 81230
rect 21982 81282 22034 81294
rect 21982 81218 22034 81230
rect 25454 81282 25506 81294
rect 25454 81218 25506 81230
rect 27694 81282 27746 81294
rect 27694 81218 27746 81230
rect 28702 81282 28754 81294
rect 31042 81230 31054 81282
rect 31106 81230 31118 81282
rect 28702 81218 28754 81230
rect 9662 81170 9714 81182
rect 6514 81118 6526 81170
rect 6578 81118 6590 81170
rect 9662 81106 9714 81118
rect 9774 81170 9826 81182
rect 9774 81106 9826 81118
rect 9998 81170 10050 81182
rect 13470 81170 13522 81182
rect 20862 81170 20914 81182
rect 13234 81118 13246 81170
rect 13298 81118 13310 81170
rect 17378 81118 17390 81170
rect 17442 81118 17454 81170
rect 9998 81106 10050 81118
rect 13470 81106 13522 81118
rect 20862 81106 20914 81118
rect 21198 81170 21250 81182
rect 21198 81106 21250 81118
rect 21422 81170 21474 81182
rect 21422 81106 21474 81118
rect 22094 81170 22146 81182
rect 22094 81106 22146 81118
rect 22430 81170 22482 81182
rect 24558 81170 24610 81182
rect 22642 81118 22654 81170
rect 22706 81118 22718 81170
rect 23090 81118 23102 81170
rect 23154 81118 23166 81170
rect 24322 81118 24334 81170
rect 24386 81118 24398 81170
rect 22430 81106 22482 81118
rect 24558 81106 24610 81118
rect 25230 81170 25282 81182
rect 26462 81170 26514 81182
rect 27470 81170 27522 81182
rect 25666 81118 25678 81170
rect 25730 81118 25742 81170
rect 25890 81118 25902 81170
rect 25954 81118 25966 81170
rect 27122 81118 27134 81170
rect 27186 81118 27198 81170
rect 25230 81106 25282 81118
rect 26462 81106 26514 81118
rect 27470 81106 27522 81118
rect 27918 81170 27970 81182
rect 28478 81170 28530 81182
rect 28242 81118 28254 81170
rect 28306 81118 28318 81170
rect 27918 81106 27970 81118
rect 28478 81106 28530 81118
rect 28814 81170 28866 81182
rect 29026 81118 29038 81170
rect 29090 81118 29102 81170
rect 30706 81118 30718 81170
rect 30770 81118 30782 81170
rect 28814 81106 28866 81118
rect 8990 81058 9042 81070
rect 3714 81006 3726 81058
rect 3778 81006 3790 81058
rect 8990 80994 9042 81006
rect 10670 81058 10722 81070
rect 10670 80994 10722 81006
rect 12574 81058 12626 81070
rect 12574 80994 12626 81006
rect 14030 81058 14082 81070
rect 14030 80994 14082 81006
rect 16382 81058 16434 81070
rect 20638 81058 20690 81070
rect 26686 81058 26738 81070
rect 20290 81006 20302 81058
rect 20354 81006 20366 81058
rect 25442 81006 25454 81058
rect 25506 81006 25518 81058
rect 16382 80994 16434 81006
rect 20638 80994 20690 81006
rect 26686 80994 26738 81006
rect 21982 80946 22034 80958
rect 26910 80946 26962 80958
rect 23986 80894 23998 80946
rect 24050 80894 24062 80946
rect 29041 80943 29087 81118
rect 29262 81058 29314 81070
rect 29262 80994 29314 81006
rect 29934 80946 29986 80958
rect 29586 80943 29598 80946
rect 29041 80897 29598 80943
rect 29586 80894 29598 80897
rect 29650 80894 29662 80946
rect 21982 80882 22034 80894
rect 26910 80882 26962 80894
rect 29934 80882 29986 80894
rect 30270 80946 30322 80958
rect 30270 80882 30322 80894
rect 1344 80778 38640 80812
rect 1344 80726 4478 80778
rect 4530 80726 4582 80778
rect 4634 80726 4686 80778
rect 4738 80726 35198 80778
rect 35250 80726 35302 80778
rect 35354 80726 35406 80778
rect 35458 80726 38640 80778
rect 1344 80692 38640 80726
rect 17390 80610 17442 80622
rect 20302 80610 20354 80622
rect 19282 80558 19294 80610
rect 19346 80558 19358 80610
rect 17390 80546 17442 80558
rect 20302 80546 20354 80558
rect 29710 80610 29762 80622
rect 29710 80546 29762 80558
rect 17054 80498 17106 80510
rect 29262 80498 29314 80510
rect 27682 80446 27694 80498
rect 27746 80446 27758 80498
rect 17054 80434 17106 80446
rect 29262 80434 29314 80446
rect 20078 80386 20130 80398
rect 16482 80334 16494 80386
rect 16546 80334 16558 80386
rect 19394 80334 19406 80386
rect 19458 80334 19470 80386
rect 20078 80322 20130 80334
rect 20526 80386 20578 80398
rect 20526 80322 20578 80334
rect 20638 80386 20690 80398
rect 28478 80386 28530 80398
rect 21522 80334 21534 80386
rect 21586 80334 21598 80386
rect 22082 80334 22094 80386
rect 22146 80334 22158 80386
rect 20638 80322 20690 80334
rect 28478 80322 28530 80334
rect 30046 80386 30098 80398
rect 30706 80334 30718 80386
rect 30770 80334 30782 80386
rect 30046 80322 30098 80334
rect 11902 80274 11954 80286
rect 11902 80210 11954 80222
rect 17614 80274 17666 80286
rect 28142 80274 28194 80286
rect 18050 80222 18062 80274
rect 18114 80222 18126 80274
rect 25442 80222 25454 80274
rect 25506 80222 25518 80274
rect 27906 80222 27918 80274
rect 27970 80222 27982 80274
rect 30818 80222 30830 80274
rect 30882 80222 30894 80274
rect 17614 80210 17666 80222
rect 28142 80210 28194 80222
rect 11566 80162 11618 80174
rect 20638 80162 20690 80174
rect 16706 80110 16718 80162
rect 16770 80110 16782 80162
rect 11566 80098 11618 80110
rect 20638 80098 20690 80110
rect 21534 80162 21586 80174
rect 21534 80098 21586 80110
rect 28254 80162 28306 80174
rect 28254 80098 28306 80110
rect 1344 79994 38640 80028
rect 1344 79942 19838 79994
rect 19890 79942 19942 79994
rect 19994 79942 20046 79994
rect 20098 79942 38640 79994
rect 1344 79908 38640 79942
rect 15374 79826 15426 79838
rect 15374 79762 15426 79774
rect 17614 79826 17666 79838
rect 17614 79762 17666 79774
rect 6078 79714 6130 79726
rect 17950 79714 18002 79726
rect 11330 79662 11342 79714
rect 11394 79662 11406 79714
rect 6078 79650 6130 79662
rect 17950 79650 18002 79662
rect 23326 79714 23378 79726
rect 31490 79662 31502 79714
rect 31554 79662 31566 79714
rect 31938 79662 31950 79714
rect 32002 79662 32014 79714
rect 23326 79650 23378 79662
rect 5966 79602 6018 79614
rect 5966 79538 6018 79550
rect 6302 79602 6354 79614
rect 14142 79602 14194 79614
rect 10546 79550 10558 79602
rect 10610 79550 10622 79602
rect 6302 79538 6354 79550
rect 14142 79538 14194 79550
rect 18286 79602 18338 79614
rect 18286 79538 18338 79550
rect 18622 79602 18674 79614
rect 23438 79602 23490 79614
rect 19058 79550 19070 79602
rect 19122 79550 19134 79602
rect 22306 79550 22318 79602
rect 22370 79550 22382 79602
rect 22642 79550 22654 79602
rect 22706 79550 22718 79602
rect 18622 79538 18674 79550
rect 23438 79538 23490 79550
rect 23662 79602 23714 79614
rect 23662 79538 23714 79550
rect 23886 79602 23938 79614
rect 25890 79550 25902 79602
rect 25954 79550 25966 79602
rect 23886 79538 23938 79550
rect 5630 79490 5682 79502
rect 5630 79426 5682 79438
rect 6862 79490 6914 79502
rect 6862 79426 6914 79438
rect 7198 79490 7250 79502
rect 7198 79426 7250 79438
rect 9662 79490 9714 79502
rect 9662 79426 9714 79438
rect 13470 79490 13522 79502
rect 13470 79426 13522 79438
rect 16382 79490 16434 79502
rect 16382 79426 16434 79438
rect 16830 79490 16882 79502
rect 16830 79426 16882 79438
rect 18398 79490 18450 79502
rect 24446 79490 24498 79502
rect 33294 79490 33346 79502
rect 22418 79438 22430 79490
rect 22482 79438 22494 79490
rect 27234 79438 27246 79490
rect 27298 79438 27310 79490
rect 18398 79426 18450 79438
rect 24446 79426 24498 79438
rect 33294 79426 33346 79438
rect 21198 79378 21250 79390
rect 30942 79378 30994 79390
rect 21858 79326 21870 79378
rect 21922 79326 21934 79378
rect 24434 79326 24446 79378
rect 24498 79375 24510 79378
rect 24770 79375 24782 79378
rect 24498 79329 24782 79375
rect 24498 79326 24510 79329
rect 24770 79326 24782 79329
rect 24834 79326 24846 79378
rect 21198 79314 21250 79326
rect 30942 79314 30994 79326
rect 31278 79378 31330 79390
rect 31278 79314 31330 79326
rect 1344 79210 38640 79244
rect 1344 79158 4478 79210
rect 4530 79158 4582 79210
rect 4634 79158 4686 79210
rect 4738 79158 35198 79210
rect 35250 79158 35302 79210
rect 35354 79158 35406 79210
rect 35458 79158 38640 79210
rect 1344 79124 38640 79158
rect 11902 79042 11954 79054
rect 11902 78978 11954 78990
rect 12238 78930 12290 78942
rect 25006 78930 25058 78942
rect 10098 78878 10110 78930
rect 10162 78878 10174 78930
rect 19058 78878 19070 78930
rect 19122 78878 19134 78930
rect 12238 78866 12290 78878
rect 25006 78866 25058 78878
rect 25342 78930 25394 78942
rect 25342 78866 25394 78878
rect 25790 78930 25842 78942
rect 28030 78930 28082 78942
rect 27346 78878 27358 78930
rect 27410 78878 27422 78930
rect 25790 78866 25842 78878
rect 28030 78866 28082 78878
rect 29150 78930 29202 78942
rect 29150 78866 29202 78878
rect 29710 78930 29762 78942
rect 31502 78930 31554 78942
rect 30482 78878 30494 78930
rect 30546 78878 30558 78930
rect 29710 78866 29762 78878
rect 31502 78866 31554 78878
rect 32398 78930 32450 78942
rect 32398 78866 32450 78878
rect 33294 78930 33346 78942
rect 33294 78866 33346 78878
rect 33742 78930 33794 78942
rect 33742 78866 33794 78878
rect 6302 78818 6354 78830
rect 11566 78818 11618 78830
rect 7522 78766 7534 78818
rect 7586 78766 7598 78818
rect 10658 78766 10670 78818
rect 10722 78766 10734 78818
rect 6302 78754 6354 78766
rect 11566 78754 11618 78766
rect 12462 78818 12514 78830
rect 12462 78754 12514 78766
rect 14590 78818 14642 78830
rect 14590 78754 14642 78766
rect 14926 78818 14978 78830
rect 14926 78754 14978 78766
rect 15038 78818 15090 78830
rect 20078 78818 20130 78830
rect 16258 78766 16270 78818
rect 16322 78766 16334 78818
rect 15038 78754 15090 78766
rect 20078 78754 20130 78766
rect 20526 78818 20578 78830
rect 20526 78754 20578 78766
rect 23998 78818 24050 78830
rect 23998 78754 24050 78766
rect 24558 78818 24610 78830
rect 24558 78754 24610 78766
rect 26126 78818 26178 78830
rect 27694 78818 27746 78830
rect 27234 78766 27246 78818
rect 27298 78766 27310 78818
rect 26126 78754 26178 78766
rect 27694 78754 27746 78766
rect 28366 78818 28418 78830
rect 28366 78754 28418 78766
rect 29486 78818 29538 78830
rect 29486 78754 29538 78766
rect 30606 78818 30658 78830
rect 31390 78818 31442 78830
rect 31042 78766 31054 78818
rect 31106 78766 31118 78818
rect 30606 78754 30658 78766
rect 31390 78754 31442 78766
rect 31838 78818 31890 78830
rect 31838 78754 31890 78766
rect 5966 78706 6018 78718
rect 5966 78642 6018 78654
rect 6526 78706 6578 78718
rect 20638 78706 20690 78718
rect 8866 78654 8878 78706
rect 8930 78654 8942 78706
rect 16930 78654 16942 78706
rect 16994 78654 17006 78706
rect 6526 78642 6578 78654
rect 20638 78642 20690 78654
rect 23438 78706 23490 78718
rect 23438 78642 23490 78654
rect 24110 78706 24162 78718
rect 24110 78642 24162 78654
rect 24782 78706 24834 78718
rect 24782 78642 24834 78654
rect 25678 78706 25730 78718
rect 25678 78642 25730 78654
rect 26014 78706 26066 78718
rect 28590 78706 28642 78718
rect 27122 78654 27134 78706
rect 27186 78654 27198 78706
rect 26014 78642 26066 78654
rect 28590 78642 28642 78654
rect 31726 78706 31778 78718
rect 31726 78642 31778 78654
rect 34974 78706 35026 78718
rect 34974 78642 35026 78654
rect 6302 78594 6354 78606
rect 6302 78530 6354 78542
rect 10110 78594 10162 78606
rect 10110 78530 10162 78542
rect 10222 78594 10274 78606
rect 10222 78530 10274 78542
rect 10446 78594 10498 78606
rect 10446 78530 10498 78542
rect 11118 78594 11170 78606
rect 11118 78530 11170 78542
rect 14366 78594 14418 78606
rect 14366 78530 14418 78542
rect 14702 78594 14754 78606
rect 14702 78530 14754 78542
rect 15822 78594 15874 78606
rect 15822 78530 15874 78542
rect 19854 78594 19906 78606
rect 19854 78530 19906 78542
rect 20750 78594 20802 78606
rect 20750 78530 20802 78542
rect 21646 78594 21698 78606
rect 21646 78530 21698 78542
rect 21870 78594 21922 78606
rect 21870 78530 21922 78542
rect 21982 78594 22034 78606
rect 21982 78530 22034 78542
rect 22094 78594 22146 78606
rect 22094 78530 22146 78542
rect 22542 78594 22594 78606
rect 22542 78530 22594 78542
rect 22766 78594 22818 78606
rect 22766 78530 22818 78542
rect 22878 78594 22930 78606
rect 22878 78530 22930 78542
rect 22990 78594 23042 78606
rect 22990 78530 23042 78542
rect 24334 78594 24386 78606
rect 24334 78530 24386 78542
rect 27470 78594 27522 78606
rect 27470 78530 27522 78542
rect 30494 78594 30546 78606
rect 30494 78530 30546 78542
rect 30830 78594 30882 78606
rect 30830 78530 30882 78542
rect 32846 78594 32898 78606
rect 32846 78530 32898 78542
rect 34638 78594 34690 78606
rect 34638 78530 34690 78542
rect 34862 78594 34914 78606
rect 34862 78530 34914 78542
rect 35646 78594 35698 78606
rect 35646 78530 35698 78542
rect 35870 78594 35922 78606
rect 35870 78530 35922 78542
rect 35982 78594 36034 78606
rect 35982 78530 36034 78542
rect 36094 78594 36146 78606
rect 36094 78530 36146 78542
rect 1344 78426 38640 78460
rect 1344 78374 19838 78426
rect 19890 78374 19942 78426
rect 19994 78374 20046 78426
rect 20098 78374 38640 78426
rect 1344 78340 38640 78374
rect 6974 78258 7026 78270
rect 6974 78194 7026 78206
rect 17726 78258 17778 78270
rect 17726 78194 17778 78206
rect 18622 78258 18674 78270
rect 29150 78258 29202 78270
rect 27570 78206 27582 78258
rect 27634 78206 27646 78258
rect 18622 78194 18674 78206
rect 29150 78194 29202 78206
rect 29262 78258 29314 78270
rect 29262 78194 29314 78206
rect 29374 78258 29426 78270
rect 29374 78194 29426 78206
rect 30158 78258 30210 78270
rect 30158 78194 30210 78206
rect 31390 78258 31442 78270
rect 31390 78194 31442 78206
rect 32174 78258 32226 78270
rect 32174 78194 32226 78206
rect 33630 78258 33682 78270
rect 33630 78194 33682 78206
rect 35198 78258 35250 78270
rect 35198 78194 35250 78206
rect 35310 78258 35362 78270
rect 35310 78194 35362 78206
rect 9886 78146 9938 78158
rect 17614 78146 17666 78158
rect 26126 78146 26178 78158
rect 14018 78094 14030 78146
rect 14082 78094 14094 78146
rect 20178 78094 20190 78146
rect 20242 78094 20254 78146
rect 9886 78082 9938 78094
rect 17614 78082 17666 78094
rect 26126 78082 26178 78094
rect 34638 78146 34690 78158
rect 34638 78082 34690 78094
rect 37102 78146 37154 78158
rect 37102 78082 37154 78094
rect 17390 78034 17442 78046
rect 6514 77982 6526 78034
rect 6578 77982 6590 78034
rect 9538 77982 9550 78034
rect 9602 77982 9614 78034
rect 13346 77982 13358 78034
rect 13410 77982 13422 78034
rect 17390 77970 17442 77982
rect 17950 78034 18002 78046
rect 25790 78034 25842 78046
rect 23538 77982 23550 78034
rect 23602 77982 23614 78034
rect 17950 77970 18002 77982
rect 25790 77970 25842 77982
rect 26350 78034 26402 78046
rect 26350 77970 26402 77982
rect 26686 78034 26738 78046
rect 26686 77970 26738 77982
rect 28478 78034 28530 78046
rect 28478 77970 28530 77982
rect 29486 78034 29538 78046
rect 30270 78034 30322 78046
rect 29698 77982 29710 78034
rect 29762 77982 29774 78034
rect 29486 77970 29538 77982
rect 30270 77970 30322 77982
rect 30494 78034 30546 78046
rect 31166 78034 31218 78046
rect 30706 77982 30718 78034
rect 30770 77982 30782 78034
rect 30494 77970 30546 77982
rect 31166 77970 31218 77982
rect 31278 78034 31330 78046
rect 31278 77970 31330 77982
rect 31502 78034 31554 78046
rect 35086 78034 35138 78046
rect 37214 78034 37266 78046
rect 31714 77982 31726 78034
rect 31778 77982 31790 78034
rect 35522 77982 35534 78034
rect 35586 77982 35598 78034
rect 35858 77982 35870 78034
rect 35922 77982 35934 78034
rect 36754 77982 36766 78034
rect 36818 77982 36830 78034
rect 31502 77970 31554 77982
rect 35086 77970 35138 77982
rect 37214 77970 37266 77982
rect 8990 77922 9042 77934
rect 3602 77870 3614 77922
rect 3666 77870 3678 77922
rect 5730 77870 5742 77922
rect 5794 77870 5806 77922
rect 8990 77858 9042 77870
rect 12910 77922 12962 77934
rect 16830 77922 16882 77934
rect 16146 77870 16158 77922
rect 16210 77870 16222 77922
rect 12910 77858 12962 77870
rect 16830 77858 16882 77870
rect 24782 77922 24834 77934
rect 24782 77858 24834 77870
rect 26574 77922 26626 77934
rect 26574 77858 26626 77870
rect 27022 77922 27074 77934
rect 27022 77858 27074 77870
rect 28030 77922 28082 77934
rect 33182 77922 33234 77934
rect 30146 77870 30158 77922
rect 30210 77870 30222 77922
rect 28030 77858 28082 77870
rect 33182 77858 33234 77870
rect 34078 77922 34130 77934
rect 34078 77858 34130 77870
rect 36318 77922 36370 77934
rect 36318 77858 36370 77870
rect 9550 77810 9602 77822
rect 25566 77810 25618 77822
rect 25218 77758 25230 77810
rect 25282 77758 25294 77810
rect 9550 77746 9602 77758
rect 25566 77746 25618 77758
rect 27246 77810 27298 77822
rect 27246 77746 27298 77758
rect 34414 77810 34466 77822
rect 34414 77746 34466 77758
rect 34750 77810 34802 77822
rect 34750 77746 34802 77758
rect 36206 77810 36258 77822
rect 36206 77746 36258 77758
rect 36542 77810 36594 77822
rect 36542 77746 36594 77758
rect 1344 77642 38640 77676
rect 1344 77590 4478 77642
rect 4530 77590 4582 77642
rect 4634 77590 4686 77642
rect 4738 77590 35198 77642
rect 35250 77590 35302 77642
rect 35354 77590 35406 77642
rect 35458 77590 38640 77642
rect 1344 77556 38640 77590
rect 35198 77474 35250 77486
rect 35198 77410 35250 77422
rect 35982 77474 36034 77486
rect 35982 77410 36034 77422
rect 37214 77474 37266 77486
rect 37214 77410 37266 77422
rect 37886 77474 37938 77486
rect 37886 77410 37938 77422
rect 12126 77362 12178 77374
rect 7298 77310 7310 77362
rect 7362 77310 7374 77362
rect 9426 77310 9438 77362
rect 9490 77310 9502 77362
rect 12126 77298 12178 77310
rect 13806 77362 13858 77374
rect 13806 77298 13858 77310
rect 15038 77362 15090 77374
rect 28142 77362 28194 77374
rect 21522 77310 21534 77362
rect 21586 77310 21598 77362
rect 15038 77298 15090 77310
rect 28142 77298 28194 77310
rect 35422 77362 35474 77374
rect 37998 77362 38050 77374
rect 35634 77310 35646 77362
rect 35698 77310 35710 77362
rect 35422 77298 35474 77310
rect 37998 77298 38050 77310
rect 10670 77250 10722 77262
rect 10098 77198 10110 77250
rect 10162 77198 10174 77250
rect 10670 77186 10722 77198
rect 12574 77250 12626 77262
rect 12574 77186 12626 77198
rect 12910 77250 12962 77262
rect 12910 77186 12962 77198
rect 14478 77250 14530 77262
rect 26910 77250 26962 77262
rect 20626 77198 20638 77250
rect 20690 77198 20702 77250
rect 25442 77198 25454 77250
rect 25506 77198 25518 77250
rect 14478 77186 14530 77198
rect 26910 77186 26962 77198
rect 27246 77250 27298 77262
rect 27246 77186 27298 77198
rect 27358 77250 27410 77262
rect 27358 77186 27410 77198
rect 29262 77250 29314 77262
rect 29262 77186 29314 77198
rect 31278 77250 31330 77262
rect 31278 77186 31330 77198
rect 32062 77250 32114 77262
rect 32062 77186 32114 77198
rect 32174 77250 32226 77262
rect 32174 77186 32226 77198
rect 32510 77250 32562 77262
rect 32510 77186 32562 77198
rect 33070 77250 33122 77262
rect 33070 77186 33122 77198
rect 34750 77250 34802 77262
rect 34750 77186 34802 77198
rect 35758 77250 35810 77262
rect 35758 77186 35810 77198
rect 36430 77250 36482 77262
rect 36430 77186 36482 77198
rect 37102 77250 37154 77262
rect 37102 77186 37154 77198
rect 37438 77250 37490 77262
rect 37438 77186 37490 77198
rect 12350 77138 12402 77150
rect 12350 77074 12402 77086
rect 13694 77138 13746 77150
rect 13694 77074 13746 77086
rect 14142 77138 14194 77150
rect 14142 77074 14194 77086
rect 15150 77138 15202 77150
rect 28366 77138 28418 77150
rect 16818 77086 16830 77138
rect 16882 77086 16894 77138
rect 15150 77074 15202 77086
rect 28366 77074 28418 77086
rect 31166 77138 31218 77150
rect 31166 77074 31218 77086
rect 31502 77138 31554 77150
rect 31502 77074 31554 77086
rect 31726 77138 31778 77150
rect 31726 77074 31778 77086
rect 32398 77138 32450 77150
rect 32398 77074 32450 77086
rect 33294 77138 33346 77150
rect 33294 77074 33346 77086
rect 33630 77138 33682 77150
rect 33630 77074 33682 77086
rect 34190 77138 34242 77150
rect 34190 77074 34242 77086
rect 34526 77138 34578 77150
rect 34526 77074 34578 77086
rect 36318 77138 36370 77150
rect 36318 77074 36370 77086
rect 38110 77138 38162 77150
rect 38110 77074 38162 77086
rect 12462 77026 12514 77038
rect 12462 76962 12514 76974
rect 13918 77026 13970 77038
rect 13918 76962 13970 76974
rect 14926 77026 14978 77038
rect 14926 76962 14978 76974
rect 27134 77026 27186 77038
rect 29710 77026 29762 77038
rect 27794 76974 27806 77026
rect 27858 76974 27870 77026
rect 27134 76962 27186 76974
rect 29710 76962 29762 76974
rect 30270 77026 30322 77038
rect 30270 76962 30322 76974
rect 30606 77026 30658 77038
rect 30606 76962 30658 76974
rect 33518 77026 33570 77038
rect 33518 76962 33570 76974
rect 34302 77026 34354 77038
rect 34302 76962 34354 76974
rect 37102 77026 37154 77038
rect 37102 76962 37154 76974
rect 1344 76858 38640 76892
rect 1344 76806 19838 76858
rect 19890 76806 19942 76858
rect 19994 76806 20046 76858
rect 20098 76806 38640 76858
rect 1344 76772 38640 76806
rect 15038 76690 15090 76702
rect 15038 76626 15090 76638
rect 15486 76690 15538 76702
rect 15486 76626 15538 76638
rect 15934 76690 15986 76702
rect 15934 76626 15986 76638
rect 16606 76690 16658 76702
rect 16606 76626 16658 76638
rect 16718 76690 16770 76702
rect 16718 76626 16770 76638
rect 16830 76690 16882 76702
rect 16830 76626 16882 76638
rect 24334 76690 24386 76702
rect 24334 76626 24386 76638
rect 25342 76690 25394 76702
rect 25342 76626 25394 76638
rect 26238 76690 26290 76702
rect 26238 76626 26290 76638
rect 27806 76690 27858 76702
rect 27806 76626 27858 76638
rect 31390 76690 31442 76702
rect 31390 76626 31442 76638
rect 33406 76690 33458 76702
rect 33406 76626 33458 76638
rect 36990 76690 37042 76702
rect 36990 76626 37042 76638
rect 37662 76690 37714 76702
rect 37662 76626 37714 76638
rect 8766 76578 8818 76590
rect 17726 76578 17778 76590
rect 27022 76578 27074 76590
rect 12226 76526 12238 76578
rect 12290 76526 12302 76578
rect 20626 76526 20638 76578
rect 20690 76526 20702 76578
rect 26786 76526 26798 76578
rect 26850 76526 26862 76578
rect 8766 76514 8818 76526
rect 17726 76514 17778 76526
rect 27022 76514 27074 76526
rect 27134 76578 27186 76590
rect 27134 76514 27186 76526
rect 27246 76578 27298 76590
rect 27246 76514 27298 76526
rect 28366 76578 28418 76590
rect 31166 76578 31218 76590
rect 30482 76526 30494 76578
rect 30546 76526 30558 76578
rect 28366 76514 28418 76526
rect 31166 76514 31218 76526
rect 31502 76578 31554 76590
rect 31502 76514 31554 76526
rect 32398 76578 32450 76590
rect 32398 76514 32450 76526
rect 32622 76578 32674 76590
rect 36878 76578 36930 76590
rect 35858 76526 35870 76578
rect 35922 76526 35934 76578
rect 36418 76526 36430 76578
rect 36482 76526 36494 76578
rect 32622 76514 32674 76526
rect 36878 76514 36930 76526
rect 37886 76578 37938 76590
rect 37886 76514 37938 76526
rect 9774 76466 9826 76478
rect 9538 76414 9550 76466
rect 9602 76414 9614 76466
rect 9774 76402 9826 76414
rect 9998 76466 10050 76478
rect 16158 76466 16210 76478
rect 10210 76414 10222 76466
rect 10274 76414 10286 76466
rect 11442 76414 11454 76466
rect 11506 76414 11518 76466
rect 9998 76402 10050 76414
rect 16158 76402 16210 76414
rect 17278 76466 17330 76478
rect 17278 76402 17330 76414
rect 17838 76466 17890 76478
rect 25230 76466 25282 76478
rect 18722 76414 18734 76466
rect 18786 76414 18798 76466
rect 17838 76402 17890 76414
rect 25230 76402 25282 76414
rect 25566 76466 25618 76478
rect 25566 76402 25618 76414
rect 25790 76466 25842 76478
rect 25790 76402 25842 76414
rect 27358 76466 27410 76478
rect 27358 76402 27410 76414
rect 27582 76466 27634 76478
rect 27582 76402 27634 76414
rect 27918 76466 27970 76478
rect 27918 76402 27970 76414
rect 29598 76466 29650 76478
rect 31726 76466 31778 76478
rect 30370 76414 30382 76466
rect 30434 76414 30446 76466
rect 29598 76402 29650 76414
rect 31726 76402 31778 76414
rect 32286 76466 32338 76478
rect 32286 76402 32338 76414
rect 33294 76466 33346 76478
rect 33294 76402 33346 76414
rect 33518 76466 33570 76478
rect 33518 76402 33570 76414
rect 33966 76466 34018 76478
rect 33966 76402 34018 76414
rect 35310 76466 35362 76478
rect 35310 76402 35362 76414
rect 35646 76466 35698 76478
rect 35646 76402 35698 76414
rect 37102 76466 37154 76478
rect 37102 76402 37154 76414
rect 37438 76466 37490 76478
rect 37438 76402 37490 76414
rect 37998 76466 38050 76478
rect 37998 76402 38050 76414
rect 8318 76354 8370 76366
rect 8318 76290 8370 76302
rect 8878 76354 8930 76366
rect 8878 76290 8930 76302
rect 9886 76354 9938 76366
rect 9886 76290 9938 76302
rect 10670 76354 10722 76366
rect 10670 76290 10722 76302
rect 11118 76354 11170 76366
rect 17502 76354 17554 76366
rect 14354 76302 14366 76354
rect 14418 76302 14430 76354
rect 11118 76290 11170 76302
rect 17502 76290 17554 76302
rect 29150 76354 29202 76366
rect 29150 76290 29202 76302
rect 34750 76354 34802 76366
rect 34750 76290 34802 76302
rect 8990 76242 9042 76254
rect 8990 76178 9042 76190
rect 28254 76242 28306 76254
rect 28254 76178 28306 76190
rect 29038 76242 29090 76254
rect 29038 76178 29090 76190
rect 29934 76242 29986 76254
rect 34526 76242 34578 76254
rect 34178 76190 34190 76242
rect 34242 76190 34254 76242
rect 29934 76178 29986 76190
rect 34526 76178 34578 76190
rect 1344 76074 38640 76108
rect 1344 76022 4478 76074
rect 4530 76022 4582 76074
rect 4634 76022 4686 76074
rect 4738 76022 35198 76074
rect 35250 76022 35302 76074
rect 35354 76022 35406 76074
rect 35458 76022 38640 76074
rect 1344 75988 38640 76022
rect 19518 75906 19570 75918
rect 34078 75906 34130 75918
rect 32498 75854 32510 75906
rect 32562 75903 32574 75906
rect 33282 75903 33294 75906
rect 32562 75857 33294 75903
rect 32562 75854 32574 75857
rect 33282 75854 33294 75857
rect 33346 75854 33358 75906
rect 19518 75842 19570 75854
rect 34078 75842 34130 75854
rect 6862 75794 6914 75806
rect 11006 75794 11058 75806
rect 7634 75742 7646 75794
rect 7698 75742 7710 75794
rect 9762 75742 9774 75794
rect 9826 75742 9838 75794
rect 6862 75730 6914 75742
rect 11006 75730 11058 75742
rect 20750 75794 20802 75806
rect 29262 75794 29314 75806
rect 31054 75794 31106 75806
rect 22642 75742 22654 75794
rect 22706 75742 22718 75794
rect 26114 75742 26126 75794
rect 26178 75742 26190 75794
rect 30034 75742 30046 75794
rect 30098 75742 30110 75794
rect 20750 75730 20802 75742
rect 29262 75730 29314 75742
rect 31054 75730 31106 75742
rect 32958 75794 33010 75806
rect 32958 75730 33010 75742
rect 35534 75794 35586 75806
rect 35534 75730 35586 75742
rect 37102 75794 37154 75806
rect 37102 75730 37154 75742
rect 5966 75682 6018 75694
rect 5966 75618 6018 75630
rect 6302 75682 6354 75694
rect 6302 75618 6354 75630
rect 6526 75682 6578 75694
rect 14590 75682 14642 75694
rect 10434 75630 10446 75682
rect 10498 75630 10510 75682
rect 6526 75618 6578 75630
rect 14590 75618 14642 75630
rect 15934 75682 15986 75694
rect 30158 75682 30210 75694
rect 31278 75682 31330 75694
rect 16258 75630 16270 75682
rect 16322 75630 16334 75682
rect 21634 75630 21646 75682
rect 21698 75630 21710 75682
rect 24770 75630 24782 75682
rect 24834 75630 24846 75682
rect 30594 75630 30606 75682
rect 30658 75630 30670 75682
rect 15934 75618 15986 75630
rect 30158 75618 30210 75630
rect 31278 75618 31330 75630
rect 31838 75682 31890 75694
rect 31838 75618 31890 75630
rect 31950 75682 32002 75694
rect 31950 75618 32002 75630
rect 34414 75682 34466 75694
rect 34414 75618 34466 75630
rect 34526 75682 34578 75694
rect 34526 75618 34578 75630
rect 35198 75682 35250 75694
rect 35198 75618 35250 75630
rect 35310 75682 35362 75694
rect 35310 75618 35362 75630
rect 36094 75682 36146 75694
rect 36094 75618 36146 75630
rect 36206 75682 36258 75694
rect 36206 75618 36258 75630
rect 6078 75570 6130 75582
rect 6078 75506 6130 75518
rect 30942 75570 30994 75582
rect 30942 75506 30994 75518
rect 31502 75570 31554 75582
rect 31502 75506 31554 75518
rect 32174 75570 32226 75582
rect 32174 75506 32226 75518
rect 32398 75570 32450 75582
rect 32398 75506 32450 75518
rect 33518 75570 33570 75582
rect 33518 75506 33570 75518
rect 33966 75570 34018 75582
rect 34974 75570 35026 75582
rect 34626 75518 34638 75570
rect 34690 75518 34702 75570
rect 33966 75506 34018 75518
rect 34974 75506 35026 75518
rect 35646 75570 35698 75582
rect 35646 75506 35698 75518
rect 36990 75570 37042 75582
rect 36990 75506 37042 75518
rect 37214 75570 37266 75582
rect 37214 75506 37266 75518
rect 7310 75458 7362 75470
rect 7310 75394 7362 75406
rect 15038 75458 15090 75470
rect 15038 75394 15090 75406
rect 30046 75458 30098 75470
rect 30046 75394 30098 75406
rect 30382 75458 30434 75470
rect 30382 75394 30434 75406
rect 33742 75458 33794 75470
rect 33742 75394 33794 75406
rect 35870 75458 35922 75470
rect 35870 75394 35922 75406
rect 37438 75458 37490 75470
rect 37438 75394 37490 75406
rect 1344 75290 38640 75324
rect 1344 75238 19838 75290
rect 19890 75238 19942 75290
rect 19994 75238 20046 75290
rect 20098 75238 38640 75290
rect 1344 75204 38640 75238
rect 17726 75122 17778 75134
rect 17726 75058 17778 75070
rect 24558 75122 24610 75134
rect 31726 75122 31778 75134
rect 25218 75070 25230 75122
rect 25282 75070 25294 75122
rect 27458 75070 27470 75122
rect 27522 75070 27534 75122
rect 24558 75058 24610 75070
rect 31726 75058 31778 75070
rect 32510 75122 32562 75134
rect 32510 75058 32562 75070
rect 33070 75122 33122 75134
rect 33070 75058 33122 75070
rect 33742 75122 33794 75134
rect 33742 75058 33794 75070
rect 33966 75122 34018 75134
rect 33966 75058 34018 75070
rect 35310 75122 35362 75134
rect 36766 75122 36818 75134
rect 36306 75070 36318 75122
rect 36370 75070 36382 75122
rect 35310 75058 35362 75070
rect 36766 75058 36818 75070
rect 8766 75010 8818 75022
rect 8766 74946 8818 74958
rect 23774 75010 23826 75022
rect 23774 74946 23826 74958
rect 24446 75010 24498 75022
rect 33406 75010 33458 75022
rect 26450 74958 26462 75010
rect 26514 74958 26526 75010
rect 27122 74958 27134 75010
rect 27186 74958 27198 75010
rect 29026 74958 29038 75010
rect 29090 74958 29102 75010
rect 24446 74946 24498 74958
rect 33406 74946 33458 74958
rect 34078 75010 34130 75022
rect 34078 74946 34130 74958
rect 35422 75010 35474 75022
rect 35422 74946 35474 74958
rect 36654 75010 36706 75022
rect 36654 74946 36706 74958
rect 37214 75010 37266 75022
rect 37214 74946 37266 74958
rect 7758 74898 7810 74910
rect 7186 74846 7198 74898
rect 7250 74846 7262 74898
rect 7758 74834 7810 74846
rect 7870 74898 7922 74910
rect 7870 74834 7922 74846
rect 8318 74898 8370 74910
rect 17950 74898 18002 74910
rect 11330 74846 11342 74898
rect 11394 74846 11406 74898
rect 8318 74834 8370 74846
rect 17950 74834 18002 74846
rect 18174 74898 18226 74910
rect 18174 74834 18226 74846
rect 18510 74898 18562 74910
rect 22430 74898 22482 74910
rect 19058 74846 19070 74898
rect 19122 74846 19134 74898
rect 18510 74834 18562 74846
rect 22430 74834 22482 74846
rect 22878 74898 22930 74910
rect 22878 74834 22930 74846
rect 22990 74898 23042 74910
rect 22990 74834 23042 74846
rect 23102 74898 23154 74910
rect 23102 74834 23154 74846
rect 23326 74898 23378 74910
rect 23326 74834 23378 74846
rect 23886 74898 23938 74910
rect 23886 74834 23938 74846
rect 24782 74898 24834 74910
rect 24782 74834 24834 74846
rect 25790 74898 25842 74910
rect 30494 74898 30546 74910
rect 34750 74898 34802 74910
rect 26786 74846 26798 74898
rect 26850 74846 26862 74898
rect 27570 74846 27582 74898
rect 27634 74846 27646 74898
rect 28466 74846 28478 74898
rect 28530 74846 28542 74898
rect 29138 74846 29150 74898
rect 29202 74846 29214 74898
rect 30146 74846 30158 74898
rect 30210 74846 30222 74898
rect 30594 74846 30606 74898
rect 30658 74846 30670 74898
rect 25790 74834 25842 74846
rect 30494 74834 30546 74846
rect 34750 74834 34802 74846
rect 34974 74898 35026 74910
rect 34974 74834 35026 74846
rect 36878 74898 36930 74910
rect 36878 74834 36930 74846
rect 38222 74898 38274 74910
rect 38222 74834 38274 74846
rect 8094 74786 8146 74798
rect 4386 74734 4398 74786
rect 4450 74734 4462 74786
rect 6514 74734 6526 74786
rect 6578 74734 6590 74786
rect 8094 74722 8146 74734
rect 11006 74786 11058 74798
rect 18062 74786 18114 74798
rect 23550 74786 23602 74798
rect 35758 74786 35810 74798
rect 13682 74734 13694 74786
rect 13746 74734 13758 74786
rect 19730 74734 19742 74786
rect 19794 74734 19806 74786
rect 21858 74734 21870 74786
rect 21922 74734 21934 74786
rect 29250 74734 29262 74786
rect 29314 74734 29326 74786
rect 11006 74722 11058 74734
rect 18062 74722 18114 74734
rect 23550 74722 23602 74734
rect 35758 74722 35810 74734
rect 37662 74786 37714 74798
rect 37662 74722 37714 74734
rect 25566 74674 25618 74686
rect 35982 74674 36034 74686
rect 34402 74622 34414 74674
rect 34466 74622 34478 74674
rect 25566 74610 25618 74622
rect 35982 74610 36034 74622
rect 1344 74506 38640 74540
rect 1344 74454 4478 74506
rect 4530 74454 4582 74506
rect 4634 74454 4686 74506
rect 4738 74454 35198 74506
rect 35250 74454 35302 74506
rect 35354 74454 35406 74506
rect 35458 74454 38640 74506
rect 1344 74420 38640 74454
rect 27806 74338 27858 74350
rect 35758 74338 35810 74350
rect 7186 74286 7198 74338
rect 7250 74335 7262 74338
rect 7746 74335 7758 74338
rect 7250 74289 7758 74335
rect 7250 74286 7262 74289
rect 7746 74286 7758 74289
rect 7810 74286 7822 74338
rect 18834 74286 18846 74338
rect 18898 74335 18910 74338
rect 19618 74335 19630 74338
rect 18898 74289 19630 74335
rect 18898 74286 18910 74289
rect 19618 74286 19630 74289
rect 19682 74286 19694 74338
rect 29698 74286 29710 74338
rect 29762 74335 29774 74338
rect 30146 74335 30158 74338
rect 29762 74289 30158 74335
rect 29762 74286 29774 74289
rect 30146 74286 30158 74289
rect 30210 74286 30222 74338
rect 27806 74274 27858 74286
rect 35758 74274 35810 74286
rect 36206 74338 36258 74350
rect 36206 74274 36258 74286
rect 7758 74226 7810 74238
rect 2146 74174 2158 74226
rect 2210 74174 2222 74226
rect 4274 74174 4286 74226
rect 4338 74174 4350 74226
rect 7758 74162 7810 74174
rect 8430 74226 8482 74238
rect 8430 74162 8482 74174
rect 19070 74226 19122 74238
rect 19070 74162 19122 74174
rect 19966 74226 20018 74238
rect 19966 74162 20018 74174
rect 21422 74226 21474 74238
rect 29822 74226 29874 74238
rect 23650 74174 23662 74226
rect 23714 74174 23726 74226
rect 21422 74162 21474 74174
rect 29822 74162 29874 74174
rect 30270 74226 30322 74238
rect 30270 74162 30322 74174
rect 30718 74226 30770 74238
rect 30718 74162 30770 74174
rect 38334 74226 38386 74238
rect 38334 74162 38386 74174
rect 5742 74114 5794 74126
rect 5058 74062 5070 74114
rect 5122 74062 5134 74114
rect 5742 74050 5794 74062
rect 6078 74114 6130 74126
rect 6078 74050 6130 74062
rect 6638 74114 6690 74126
rect 6638 74050 6690 74062
rect 6974 74114 7026 74126
rect 6974 74050 7026 74062
rect 7310 74114 7362 74126
rect 19854 74114 19906 74126
rect 14354 74062 14366 74114
rect 14418 74062 14430 74114
rect 7310 74050 7362 74062
rect 19854 74050 19906 74062
rect 20078 74114 20130 74126
rect 20078 74050 20130 74062
rect 20526 74114 20578 74126
rect 28142 74114 28194 74126
rect 26114 74062 26126 74114
rect 26178 74062 26190 74114
rect 20526 74050 20578 74062
rect 28142 74050 28194 74062
rect 28366 74114 28418 74126
rect 28366 74050 28418 74062
rect 33742 74114 33794 74126
rect 33742 74050 33794 74062
rect 33966 74114 34018 74126
rect 33966 74050 34018 74062
rect 34974 74114 35026 74126
rect 34974 74050 35026 74062
rect 35310 74114 35362 74126
rect 35310 74050 35362 74062
rect 35646 74114 35698 74126
rect 35646 74050 35698 74062
rect 36318 74114 36370 74126
rect 36318 74050 36370 74062
rect 5854 74002 5906 74014
rect 5854 73938 5906 73950
rect 6750 74002 6802 74014
rect 29262 74002 29314 74014
rect 15810 73950 15822 74002
rect 15874 73950 15886 74002
rect 6750 73938 6802 73950
rect 29262 73938 29314 73950
rect 29374 74002 29426 74014
rect 29374 73938 29426 73950
rect 33518 74002 33570 74014
rect 33518 73938 33570 73950
rect 35198 74002 35250 74014
rect 35198 73938 35250 73950
rect 19518 73890 19570 73902
rect 19518 73826 19570 73838
rect 29038 73890 29090 73902
rect 29038 73826 29090 73838
rect 33854 73890 33906 73902
rect 33854 73826 33906 73838
rect 35758 73890 35810 73902
rect 35758 73826 35810 73838
rect 1344 73722 38640 73756
rect 1344 73670 19838 73722
rect 19890 73670 19942 73722
rect 19994 73670 20046 73722
rect 20098 73670 38640 73722
rect 1344 73636 38640 73670
rect 5294 73554 5346 73566
rect 5294 73490 5346 73502
rect 6190 73554 6242 73566
rect 6190 73490 6242 73502
rect 17502 73554 17554 73566
rect 17502 73490 17554 73502
rect 17838 73554 17890 73566
rect 17838 73490 17890 73502
rect 17950 73554 18002 73566
rect 17950 73490 18002 73502
rect 18846 73554 18898 73566
rect 18846 73490 18898 73502
rect 26238 73554 26290 73566
rect 30494 73554 30546 73566
rect 27234 73502 27246 73554
rect 27298 73502 27310 73554
rect 28690 73502 28702 73554
rect 28754 73502 28766 73554
rect 26238 73490 26290 73502
rect 30494 73490 30546 73502
rect 31502 73554 31554 73566
rect 31502 73490 31554 73502
rect 29822 73442 29874 73454
rect 16034 73390 16046 73442
rect 16098 73390 16110 73442
rect 23090 73390 23102 73442
rect 23154 73390 23166 73442
rect 29822 73378 29874 73390
rect 31054 73442 31106 73454
rect 31054 73378 31106 73390
rect 17726 73330 17778 73342
rect 28366 73330 28418 73342
rect 16818 73278 16830 73330
rect 16882 73278 16894 73330
rect 19394 73278 19406 73330
rect 19458 73278 19470 73330
rect 26114 73278 26126 73330
rect 26178 73278 26190 73330
rect 26898 73278 26910 73330
rect 26962 73278 26974 73330
rect 17726 73266 17778 73278
rect 28366 73266 28418 73278
rect 29038 73330 29090 73342
rect 29038 73266 29090 73278
rect 29598 73330 29650 73342
rect 30146 73278 30158 73330
rect 30210 73278 30222 73330
rect 29598 73266 29650 73278
rect 18398 73218 18450 73230
rect 29262 73218 29314 73230
rect 13906 73166 13918 73218
rect 13970 73166 13982 73218
rect 26226 73166 26238 73218
rect 26290 73166 26302 73218
rect 18398 73154 18450 73166
rect 29262 73154 29314 73166
rect 29710 73218 29762 73230
rect 29710 73154 29762 73166
rect 30606 73218 30658 73230
rect 30606 73154 30658 73166
rect 1344 72938 38640 72972
rect 1344 72886 4478 72938
rect 4530 72886 4582 72938
rect 4634 72886 4686 72938
rect 4738 72886 35198 72938
rect 35250 72886 35302 72938
rect 35354 72886 35406 72938
rect 35458 72886 38640 72938
rect 1344 72852 38640 72886
rect 28254 72770 28306 72782
rect 28254 72706 28306 72718
rect 22206 72658 22258 72670
rect 31950 72658 32002 72670
rect 15138 72606 15150 72658
rect 15202 72606 15214 72658
rect 29810 72606 29822 72658
rect 29874 72606 29886 72658
rect 35074 72606 35086 72658
rect 35138 72606 35150 72658
rect 22206 72594 22258 72606
rect 31950 72594 32002 72606
rect 20414 72546 20466 72558
rect 31278 72546 31330 72558
rect 11778 72494 11790 72546
rect 11842 72494 11854 72546
rect 13682 72494 13694 72546
rect 13746 72494 13758 72546
rect 19954 72494 19966 72546
rect 20018 72494 20030 72546
rect 27794 72494 27806 72546
rect 27858 72494 27870 72546
rect 29362 72494 29374 72546
rect 29426 72494 29438 72546
rect 20414 72482 20466 72494
rect 31278 72482 31330 72494
rect 28254 72434 28306 72446
rect 24994 72382 25006 72434
rect 25058 72382 25070 72434
rect 28254 72370 28306 72382
rect 28366 72434 28418 72446
rect 29250 72382 29262 72434
rect 29314 72382 29326 72434
rect 28366 72370 28418 72382
rect 11566 72322 11618 72334
rect 11566 72258 11618 72270
rect 13470 72322 13522 72334
rect 13470 72258 13522 72270
rect 33630 72322 33682 72334
rect 33630 72258 33682 72270
rect 34078 72322 34130 72334
rect 34078 72258 34130 72270
rect 34638 72322 34690 72334
rect 34638 72258 34690 72270
rect 35646 72322 35698 72334
rect 35646 72258 35698 72270
rect 36094 72322 36146 72334
rect 36094 72258 36146 72270
rect 1344 72154 38640 72188
rect 1344 72102 19838 72154
rect 19890 72102 19942 72154
rect 19994 72102 20046 72154
rect 20098 72102 38640 72154
rect 1344 72068 38640 72102
rect 26126 71986 26178 71998
rect 26126 71922 26178 71934
rect 26238 71986 26290 71998
rect 26238 71922 26290 71934
rect 32398 71986 32450 71998
rect 32398 71922 32450 71934
rect 36766 71986 36818 71998
rect 36766 71922 36818 71934
rect 8542 71874 8594 71886
rect 33294 71874 33346 71886
rect 34862 71874 34914 71886
rect 22530 71822 22542 71874
rect 22594 71822 22606 71874
rect 29922 71822 29934 71874
rect 29986 71822 29998 71874
rect 34402 71822 34414 71874
rect 34466 71822 34478 71874
rect 8542 71810 8594 71822
rect 33294 71810 33346 71822
rect 34862 71810 34914 71822
rect 35982 71874 36034 71886
rect 35982 71810 36034 71822
rect 8878 71762 8930 71774
rect 14478 71762 14530 71774
rect 11106 71710 11118 71762
rect 11170 71710 11182 71762
rect 8878 71698 8930 71710
rect 14478 71698 14530 71710
rect 17502 71762 17554 71774
rect 25566 71762 25618 71774
rect 18834 71710 18846 71762
rect 18898 71710 18910 71762
rect 21858 71710 21870 71762
rect 21922 71710 21934 71762
rect 17502 71698 17554 71710
rect 25566 71698 25618 71710
rect 26014 71762 26066 71774
rect 34974 71762 35026 71774
rect 27794 71710 27806 71762
rect 27858 71710 27870 71762
rect 34178 71710 34190 71762
rect 34242 71710 34254 71762
rect 26014 71698 26066 71710
rect 34974 71698 35026 71710
rect 36094 71762 36146 71774
rect 36306 71710 36318 71762
rect 36370 71710 36382 71762
rect 36094 71698 36146 71710
rect 9998 71650 10050 71662
rect 25790 71650 25842 71662
rect 37214 71650 37266 71662
rect 11778 71598 11790 71650
rect 11842 71598 11854 71650
rect 13906 71598 13918 71650
rect 13970 71598 13982 71650
rect 21074 71598 21086 71650
rect 21138 71598 21150 71650
rect 24658 71598 24670 71650
rect 24722 71598 24734 71650
rect 33954 71598 33966 71650
rect 34018 71598 34030 71650
rect 9998 71586 10050 71598
rect 25790 71586 25842 71598
rect 37214 71586 37266 71598
rect 37662 71650 37714 71662
rect 37662 71586 37714 71598
rect 33406 71538 33458 71550
rect 33406 71474 33458 71486
rect 34862 71538 34914 71550
rect 35522 71486 35534 71538
rect 35586 71486 35598 71538
rect 34862 71474 34914 71486
rect 1344 71370 38640 71404
rect 1344 71318 4478 71370
rect 4530 71318 4582 71370
rect 4634 71318 4686 71370
rect 4738 71318 35198 71370
rect 35250 71318 35302 71370
rect 35354 71318 35406 71370
rect 35458 71318 38640 71370
rect 1344 71284 38640 71318
rect 13806 71202 13858 71214
rect 13458 71150 13470 71202
rect 13522 71150 13534 71202
rect 13806 71138 13858 71150
rect 14478 71090 14530 71102
rect 18286 71090 18338 71102
rect 25006 71090 25058 71102
rect 37214 71090 37266 71102
rect 7522 71038 7534 71090
rect 7586 71038 7598 71090
rect 9650 71038 9662 71090
rect 9714 71038 9726 71090
rect 10770 71038 10782 71090
rect 10834 71038 10846 71090
rect 12898 71038 12910 71090
rect 12962 71038 12974 71090
rect 17826 71038 17838 71090
rect 17890 71038 17902 71090
rect 22418 71038 22430 71090
rect 22482 71038 22494 71090
rect 30146 71038 30158 71090
rect 30210 71038 30222 71090
rect 32498 71038 32510 71090
rect 32562 71038 32574 71090
rect 14478 71026 14530 71038
rect 18286 71026 18338 71038
rect 25006 71026 25058 71038
rect 37214 71026 37266 71038
rect 14030 70978 14082 70990
rect 25230 70978 25282 70990
rect 6738 70926 6750 70978
rect 6802 70926 6814 70978
rect 9986 70926 9998 70978
rect 10050 70926 10062 70978
rect 15026 70926 15038 70978
rect 15090 70926 15102 70978
rect 23874 70926 23886 70978
rect 23938 70926 23950 70978
rect 14030 70914 14082 70926
rect 25230 70914 25282 70926
rect 25566 70978 25618 70990
rect 29374 70978 29426 70990
rect 26786 70926 26798 70978
rect 26850 70926 26862 70978
rect 27346 70926 27358 70978
rect 27410 70926 27422 70978
rect 31714 70926 31726 70978
rect 31778 70926 31790 70978
rect 32722 70926 32734 70978
rect 32786 70926 32798 70978
rect 33730 70926 33742 70978
rect 33794 70926 33806 70978
rect 35298 70926 35310 70978
rect 35362 70926 35374 70978
rect 25566 70914 25618 70926
rect 29374 70914 29426 70926
rect 5630 70866 5682 70878
rect 25790 70866 25842 70878
rect 15698 70814 15710 70866
rect 15762 70814 15774 70866
rect 27682 70814 27694 70866
rect 27746 70814 27758 70866
rect 28018 70814 28030 70866
rect 28082 70814 28094 70866
rect 31042 70814 31054 70866
rect 31106 70814 31118 70866
rect 32610 70814 32622 70866
rect 32674 70814 32686 70866
rect 35410 70814 35422 70866
rect 35474 70814 35486 70866
rect 38210 70814 38222 70866
rect 38274 70814 38286 70866
rect 5630 70802 5682 70814
rect 25790 70802 25842 70814
rect 5966 70754 6018 70766
rect 5966 70690 6018 70702
rect 14590 70754 14642 70766
rect 14590 70690 14642 70702
rect 18398 70754 18450 70766
rect 18398 70690 18450 70702
rect 18846 70754 18898 70766
rect 18846 70690 18898 70702
rect 24334 70754 24386 70766
rect 24334 70690 24386 70702
rect 25454 70754 25506 70766
rect 26450 70702 26462 70754
rect 26514 70702 26526 70754
rect 27906 70702 27918 70754
rect 27970 70702 27982 70754
rect 36082 70702 36094 70754
rect 36146 70702 36158 70754
rect 25454 70690 25506 70702
rect 1344 70586 38640 70620
rect 1344 70534 19838 70586
rect 19890 70534 19942 70586
rect 19994 70534 20046 70586
rect 20098 70534 38640 70586
rect 1344 70500 38640 70534
rect 15262 70418 15314 70430
rect 11554 70366 11566 70418
rect 11618 70366 11630 70418
rect 15262 70354 15314 70366
rect 15934 70418 15986 70430
rect 15934 70354 15986 70366
rect 25342 70418 25394 70430
rect 25342 70354 25394 70366
rect 26238 70418 26290 70430
rect 26238 70354 26290 70366
rect 26462 70418 26514 70430
rect 26462 70354 26514 70366
rect 27470 70418 27522 70430
rect 27470 70354 27522 70366
rect 28142 70418 28194 70430
rect 28142 70354 28194 70366
rect 33630 70418 33682 70430
rect 33630 70354 33682 70366
rect 34078 70418 34130 70430
rect 34078 70354 34130 70366
rect 15710 70306 15762 70318
rect 6178 70254 6190 70306
rect 6242 70254 6254 70306
rect 10658 70254 10670 70306
rect 10722 70254 10734 70306
rect 12674 70254 12686 70306
rect 12738 70254 12750 70306
rect 15710 70242 15762 70254
rect 18398 70306 18450 70318
rect 18398 70242 18450 70254
rect 26686 70306 26738 70318
rect 26686 70242 26738 70254
rect 28254 70306 28306 70318
rect 30606 70306 30658 70318
rect 28914 70254 28926 70306
rect 28978 70254 28990 70306
rect 28254 70242 28306 70254
rect 30606 70242 30658 70254
rect 30830 70306 30882 70318
rect 30830 70242 30882 70254
rect 34302 70306 34354 70318
rect 34302 70242 34354 70254
rect 15598 70194 15650 70206
rect 22318 70194 22370 70206
rect 5506 70142 5518 70194
rect 5570 70142 5582 70194
rect 11890 70142 11902 70194
rect 11954 70142 11966 70194
rect 18946 70142 18958 70194
rect 19010 70142 19022 70194
rect 15598 70130 15650 70142
rect 22318 70130 22370 70142
rect 26126 70194 26178 70206
rect 26126 70130 26178 70142
rect 26798 70194 26850 70206
rect 26798 70130 26850 70142
rect 27246 70194 27298 70206
rect 27246 70130 27298 70142
rect 27582 70194 27634 70206
rect 27582 70130 27634 70142
rect 27918 70194 27970 70206
rect 30382 70194 30434 70206
rect 31838 70194 31890 70206
rect 33070 70194 33122 70206
rect 29138 70142 29150 70194
rect 29202 70142 29214 70194
rect 31154 70142 31166 70194
rect 31218 70142 31230 70194
rect 32162 70142 32174 70194
rect 32226 70142 32238 70194
rect 27918 70130 27970 70142
rect 30382 70130 30434 70142
rect 31838 70130 31890 70142
rect 33070 70130 33122 70142
rect 33294 70194 33346 70206
rect 33294 70130 33346 70142
rect 33518 70194 33570 70206
rect 33518 70130 33570 70142
rect 33742 70194 33794 70206
rect 33742 70130 33794 70142
rect 34414 70194 34466 70206
rect 34850 70142 34862 70194
rect 34914 70142 34926 70194
rect 36978 70142 36990 70194
rect 37042 70142 37054 70194
rect 34414 70130 34466 70142
rect 8766 70082 8818 70094
rect 8306 70030 8318 70082
rect 8370 70030 8382 70082
rect 8766 70018 8818 70030
rect 9886 70082 9938 70094
rect 9886 70018 9938 70030
rect 10110 70082 10162 70094
rect 10110 70018 10162 70030
rect 10334 70082 10386 70094
rect 10334 70018 10386 70030
rect 11006 70082 11058 70094
rect 16270 70082 16322 70094
rect 14802 70030 14814 70082
rect 14866 70030 14878 70082
rect 11006 70018 11058 70030
rect 16270 70018 16322 70030
rect 17838 70082 17890 70094
rect 17838 70018 17890 70030
rect 18174 70082 18226 70094
rect 25902 70082 25954 70094
rect 18498 70030 18510 70082
rect 18562 70030 18574 70082
rect 19618 70030 19630 70082
rect 19682 70030 19694 70082
rect 21746 70030 21758 70082
rect 21810 70030 21822 70082
rect 18174 70018 18226 70030
rect 25902 70018 25954 70030
rect 28478 70082 28530 70094
rect 28478 70018 28530 70030
rect 29486 70082 29538 70094
rect 37314 70030 37326 70082
rect 37378 70030 37390 70082
rect 29486 70018 29538 70030
rect 11230 69970 11282 69982
rect 11230 69906 11282 69918
rect 28702 69970 28754 69982
rect 28702 69906 28754 69918
rect 29710 69970 29762 69982
rect 32174 69970 32226 69982
rect 30034 69918 30046 69970
rect 30098 69918 30110 69970
rect 35746 69918 35758 69970
rect 35810 69918 35822 69970
rect 29710 69906 29762 69918
rect 32174 69906 32226 69918
rect 1344 69802 38640 69836
rect 1344 69750 4478 69802
rect 4530 69750 4582 69802
rect 4634 69750 4686 69802
rect 4738 69750 35198 69802
rect 35250 69750 35302 69802
rect 35354 69750 35406 69802
rect 35458 69750 38640 69802
rect 1344 69716 38640 69750
rect 9102 69634 9154 69646
rect 5618 69582 5630 69634
rect 5682 69582 5694 69634
rect 6738 69582 6750 69634
rect 6802 69631 6814 69634
rect 7074 69631 7086 69634
rect 6802 69585 7086 69631
rect 6802 69582 6814 69585
rect 7074 69582 7086 69585
rect 7138 69582 7150 69634
rect 9102 69570 9154 69582
rect 26798 69634 26850 69646
rect 26798 69570 26850 69582
rect 32174 69634 32226 69646
rect 32174 69570 32226 69582
rect 9550 69522 9602 69534
rect 5058 69470 5070 69522
rect 5122 69470 5134 69522
rect 9550 69458 9602 69470
rect 10670 69522 10722 69534
rect 10670 69458 10722 69470
rect 13582 69522 13634 69534
rect 13582 69458 13634 69470
rect 14030 69522 14082 69534
rect 14030 69458 14082 69470
rect 14478 69522 14530 69534
rect 18174 69522 18226 69534
rect 38222 69522 38274 69534
rect 17714 69470 17726 69522
rect 17778 69470 17790 69522
rect 28354 69470 28366 69522
rect 28418 69470 28430 69522
rect 31378 69470 31390 69522
rect 31442 69470 31454 69522
rect 32946 69470 32958 69522
rect 33010 69470 33022 69522
rect 35634 69470 35646 69522
rect 35698 69470 35710 69522
rect 14478 69458 14530 69470
rect 18174 69458 18226 69470
rect 38222 69458 38274 69470
rect 5966 69410 6018 69422
rect 2146 69358 2158 69410
rect 2210 69358 2222 69410
rect 5966 69346 6018 69358
rect 6190 69410 6242 69422
rect 6190 69346 6242 69358
rect 8766 69410 8818 69422
rect 8766 69346 8818 69358
rect 11230 69410 11282 69422
rect 26686 69410 26738 69422
rect 14802 69358 14814 69410
rect 14866 69358 14878 69410
rect 22082 69358 22094 69410
rect 22146 69358 22158 69410
rect 11230 69346 11282 69358
rect 26686 69346 26738 69358
rect 27358 69410 27410 69422
rect 29150 69410 29202 69422
rect 27682 69358 27694 69410
rect 27746 69358 27758 69410
rect 27358 69346 27410 69358
rect 29150 69346 29202 69358
rect 29598 69410 29650 69422
rect 30258 69358 30270 69410
rect 30322 69358 30334 69410
rect 31826 69358 31838 69410
rect 31890 69358 31902 69410
rect 32834 69358 32846 69410
rect 32898 69358 32910 69410
rect 34850 69358 34862 69410
rect 34914 69358 34926 69410
rect 35858 69358 35870 69410
rect 35922 69358 35934 69410
rect 36978 69358 36990 69410
rect 37042 69358 37054 69410
rect 29598 69346 29650 69358
rect 8542 69298 8594 69310
rect 2930 69246 2942 69298
rect 2994 69246 3006 69298
rect 8542 69234 8594 69246
rect 11566 69298 11618 69310
rect 29486 69298 29538 69310
rect 15586 69246 15598 69298
rect 15650 69246 15662 69298
rect 24434 69246 24446 69298
rect 24498 69246 24510 69298
rect 27906 69246 27918 69298
rect 27970 69246 27982 69298
rect 11566 69234 11618 69246
rect 29486 69234 29538 69246
rect 33406 69298 33458 69310
rect 37214 69298 37266 69310
rect 34514 69246 34526 69298
rect 34578 69246 34590 69298
rect 33406 69234 33458 69246
rect 37214 69234 37266 69246
rect 37326 69298 37378 69310
rect 37326 69234 37378 69246
rect 6638 69186 6690 69198
rect 6638 69122 6690 69134
rect 7086 69186 7138 69198
rect 7086 69122 7138 69134
rect 9998 69186 10050 69198
rect 9998 69122 10050 69134
rect 18062 69186 18114 69198
rect 18062 69122 18114 69134
rect 29374 69186 29426 69198
rect 29374 69122 29426 69134
rect 32062 69186 32114 69198
rect 37762 69134 37774 69186
rect 37826 69134 37838 69186
rect 32062 69122 32114 69134
rect 1344 69018 38640 69052
rect 1344 68966 19838 69018
rect 19890 68966 19942 69018
rect 19994 68966 20046 69018
rect 20098 68966 38640 69018
rect 1344 68932 38640 68966
rect 3502 68850 3554 68862
rect 3502 68786 3554 68798
rect 15822 68850 15874 68862
rect 15822 68786 15874 68798
rect 16270 68850 16322 68862
rect 16270 68786 16322 68798
rect 28254 68850 28306 68862
rect 28254 68786 28306 68798
rect 28478 68850 28530 68862
rect 28478 68786 28530 68798
rect 30942 68850 30994 68862
rect 30942 68786 30994 68798
rect 33182 68850 33234 68862
rect 33182 68786 33234 68798
rect 16382 68738 16434 68750
rect 16382 68674 16434 68686
rect 20750 68738 20802 68750
rect 20750 68674 20802 68686
rect 21198 68738 21250 68750
rect 21198 68674 21250 68686
rect 33070 68738 33122 68750
rect 33070 68674 33122 68686
rect 3838 68626 3890 68638
rect 28590 68626 28642 68638
rect 4498 68574 4510 68626
rect 4562 68574 4574 68626
rect 6066 68574 6078 68626
rect 6130 68574 6142 68626
rect 17490 68574 17502 68626
rect 17554 68574 17566 68626
rect 31602 68574 31614 68626
rect 31666 68574 31678 68626
rect 32610 68574 32622 68626
rect 32674 68574 32686 68626
rect 33954 68574 33966 68626
rect 34018 68574 34030 68626
rect 36082 68574 36094 68626
rect 36146 68574 36158 68626
rect 36754 68574 36766 68626
rect 36818 68574 36830 68626
rect 3838 68562 3890 68574
rect 28590 68562 28642 68574
rect 9550 68514 9602 68526
rect 6850 68462 6862 68514
rect 6914 68462 6926 68514
rect 8978 68462 8990 68514
rect 9042 68462 9054 68514
rect 9550 68450 9602 68462
rect 10110 68514 10162 68526
rect 10110 68450 10162 68462
rect 10558 68514 10610 68526
rect 10558 68450 10610 68462
rect 15374 68514 15426 68526
rect 29038 68514 29090 68526
rect 29486 68514 29538 68526
rect 18162 68462 18174 68514
rect 18226 68462 18238 68514
rect 20290 68462 20302 68514
rect 20354 68462 20366 68514
rect 29362 68462 29374 68514
rect 29426 68462 29438 68514
rect 15374 68450 15426 68462
rect 29038 68450 29090 68462
rect 5294 68402 5346 68414
rect 5294 68338 5346 68350
rect 9886 68402 9938 68414
rect 9886 68338 9938 68350
rect 16158 68402 16210 68414
rect 16158 68338 16210 68350
rect 21086 68402 21138 68414
rect 29377 68399 29423 68462
rect 29486 68450 29538 68462
rect 30046 68514 30098 68526
rect 30046 68450 30098 68462
rect 30382 68514 30434 68526
rect 31938 68462 31950 68514
rect 32002 68462 32014 68514
rect 34962 68462 34974 68514
rect 35026 68462 35038 68514
rect 37538 68462 37550 68514
rect 37602 68462 37614 68514
rect 30382 68450 30434 68462
rect 30370 68399 30382 68402
rect 29377 68353 30382 68399
rect 30370 68350 30382 68353
rect 30434 68350 30446 68402
rect 31826 68350 31838 68402
rect 31890 68350 31902 68402
rect 35186 68350 35198 68402
rect 35250 68350 35262 68402
rect 21086 68338 21138 68350
rect 1344 68234 38640 68268
rect 1344 68182 4478 68234
rect 4530 68182 4582 68234
rect 4634 68182 4686 68234
rect 4738 68182 35198 68234
rect 35250 68182 35302 68234
rect 35354 68182 35406 68234
rect 35458 68182 38640 68234
rect 1344 68148 38640 68182
rect 17950 68066 18002 68078
rect 8866 68014 8878 68066
rect 8930 68063 8942 68066
rect 9202 68063 9214 68066
rect 8930 68017 9214 68063
rect 8930 68014 8942 68017
rect 9202 68014 9214 68017
rect 9266 68014 9278 68066
rect 17950 68002 18002 68014
rect 31950 68066 32002 68078
rect 31950 68002 32002 68014
rect 33070 68066 33122 68078
rect 33070 68002 33122 68014
rect 34414 68066 34466 68078
rect 34414 68002 34466 68014
rect 34750 68066 34802 68078
rect 34750 68002 34802 68014
rect 36878 68066 36930 68078
rect 36878 68002 36930 68014
rect 9214 67954 9266 67966
rect 9214 67890 9266 67902
rect 18622 67954 18674 67966
rect 18622 67890 18674 67902
rect 19742 67954 19794 67966
rect 19742 67890 19794 67902
rect 20190 67954 20242 67966
rect 29598 67954 29650 67966
rect 37326 67954 37378 67966
rect 24098 67902 24110 67954
rect 24162 67902 24174 67954
rect 31714 67902 31726 67954
rect 31778 67902 31790 67954
rect 20190 67890 20242 67902
rect 29598 67890 29650 67902
rect 37326 67890 37378 67902
rect 20526 67842 20578 67854
rect 27470 67842 27522 67854
rect 27010 67790 27022 67842
rect 27074 67790 27086 67842
rect 20526 67778 20578 67790
rect 27470 67778 27522 67790
rect 31278 67842 31330 67854
rect 37550 67842 37602 67854
rect 33618 67790 33630 67842
rect 33682 67790 33694 67842
rect 35522 67790 35534 67842
rect 35586 67790 35598 67842
rect 36082 67790 36094 67842
rect 36146 67790 36158 67842
rect 31278 67778 31330 67790
rect 37550 67778 37602 67790
rect 37774 67842 37826 67854
rect 37774 67778 37826 67790
rect 3166 67730 3218 67742
rect 3166 67666 3218 67678
rect 7870 67730 7922 67742
rect 7870 67666 7922 67678
rect 8206 67730 8258 67742
rect 8206 67666 8258 67678
rect 16830 67730 16882 67742
rect 16830 67666 16882 67678
rect 17614 67730 17666 67742
rect 17614 67666 17666 67678
rect 17838 67730 17890 67742
rect 17838 67666 17890 67678
rect 20638 67730 20690 67742
rect 20638 67666 20690 67678
rect 23102 67730 23154 67742
rect 30382 67730 30434 67742
rect 26226 67678 26238 67730
rect 26290 67678 26302 67730
rect 23102 67666 23154 67678
rect 30382 67666 30434 67678
rect 30718 67730 30770 67742
rect 30718 67666 30770 67678
rect 31726 67730 31778 67742
rect 31726 67666 31778 67678
rect 33182 67730 33234 67742
rect 33842 67678 33854 67730
rect 33906 67678 33918 67730
rect 35298 67678 35310 67730
rect 35362 67678 35374 67730
rect 33182 67666 33234 67678
rect 2830 67618 2882 67630
rect 2830 67554 2882 67566
rect 5742 67618 5794 67630
rect 5742 67554 5794 67566
rect 17390 67618 17442 67630
rect 17390 67554 17442 67566
rect 19406 67618 19458 67630
rect 19406 67554 19458 67566
rect 19630 67618 19682 67630
rect 19630 67554 19682 67566
rect 20862 67618 20914 67630
rect 20862 67554 20914 67566
rect 21534 67618 21586 67630
rect 36082 67566 36094 67618
rect 36146 67566 36158 67618
rect 21534 67554 21586 67566
rect 1344 67450 38640 67484
rect 1344 67398 19838 67450
rect 19890 67398 19942 67450
rect 19994 67398 20046 67450
rect 20098 67398 38640 67450
rect 1344 67364 38640 67398
rect 35074 67230 35086 67282
rect 35138 67230 35150 67282
rect 29262 67170 29314 67182
rect 2482 67118 2494 67170
rect 2546 67118 2558 67170
rect 11106 67118 11118 67170
rect 11170 67118 11182 67170
rect 20738 67118 20750 67170
rect 20802 67118 20814 67170
rect 29262 67106 29314 67118
rect 30494 67170 30546 67182
rect 30494 67106 30546 67118
rect 33406 67170 33458 67182
rect 34178 67118 34190 67170
rect 34242 67118 34254 67170
rect 37426 67118 37438 67170
rect 37490 67118 37502 67170
rect 33406 67106 33458 67118
rect 8766 67058 8818 67070
rect 18734 67058 18786 67070
rect 29150 67058 29202 67070
rect 1810 67006 1822 67058
rect 1874 67006 1886 67058
rect 15026 67006 15038 67058
rect 15090 67006 15102 67058
rect 17602 67006 17614 67058
rect 17666 67006 17678 67058
rect 17938 67006 17950 67058
rect 18002 67006 18014 67058
rect 19282 67006 19294 67058
rect 19346 67006 19358 67058
rect 20066 67006 20078 67058
rect 20130 67006 20142 67058
rect 29474 67006 29486 67058
rect 29538 67006 29550 67058
rect 33618 67006 33630 67058
rect 33682 67006 33694 67058
rect 34290 67006 34302 67058
rect 34354 67006 34366 67058
rect 35970 67006 35982 67058
rect 36034 67006 36046 67058
rect 37874 67006 37886 67058
rect 37938 67006 37950 67058
rect 8766 66994 8818 67006
rect 18734 66994 18786 67006
rect 29150 66994 29202 67006
rect 5070 66946 5122 66958
rect 4610 66894 4622 66946
rect 4674 66894 4686 66946
rect 5070 66882 5122 66894
rect 8430 66946 8482 66958
rect 8430 66882 8482 66894
rect 8990 66946 9042 66958
rect 8990 66882 9042 66894
rect 15486 66946 15538 66958
rect 15486 66882 15538 66894
rect 16046 66946 16098 66958
rect 16046 66882 16098 66894
rect 16494 66946 16546 66958
rect 16494 66882 16546 66894
rect 16942 66946 16994 66958
rect 23438 66946 23490 66958
rect 18162 66894 18174 66946
rect 18226 66894 18238 66946
rect 22866 66894 22878 66946
rect 22930 66894 22942 66946
rect 16942 66882 16994 66894
rect 23438 66882 23490 66894
rect 23886 66946 23938 66958
rect 23886 66882 23938 66894
rect 24334 66946 24386 66958
rect 24334 66882 24386 66894
rect 24782 66946 24834 66958
rect 24782 66882 24834 66894
rect 30046 66946 30098 66958
rect 30046 66882 30098 66894
rect 30942 66946 30994 66958
rect 30942 66882 30994 66894
rect 31390 66946 31442 66958
rect 31390 66882 31442 66894
rect 15250 66782 15262 66834
rect 15314 66831 15326 66834
rect 16482 66831 16494 66834
rect 15314 66785 16494 66831
rect 15314 66782 15326 66785
rect 16482 66782 16494 66785
rect 16546 66782 16558 66834
rect 19058 66782 19070 66834
rect 19122 66782 19134 66834
rect 23986 66782 23998 66834
rect 24050 66831 24062 66834
rect 24322 66831 24334 66834
rect 24050 66785 24334 66831
rect 24050 66782 24062 66785
rect 24322 66782 24334 66785
rect 24386 66831 24398 66834
rect 24770 66831 24782 66834
rect 24386 66785 24782 66831
rect 24386 66782 24398 66785
rect 24770 66782 24782 66785
rect 24834 66782 24846 66834
rect 1344 66666 38640 66700
rect 1344 66614 4478 66666
rect 4530 66614 4582 66666
rect 4634 66614 4686 66666
rect 4738 66614 35198 66666
rect 35250 66614 35302 66666
rect 35354 66614 35406 66666
rect 35458 66614 38640 66666
rect 1344 66580 38640 66614
rect 29262 66498 29314 66510
rect 3378 66446 3390 66498
rect 3442 66446 3454 66498
rect 17378 66446 17390 66498
rect 17442 66446 17454 66498
rect 19170 66446 19182 66498
rect 19234 66446 19246 66498
rect 29262 66434 29314 66446
rect 30046 66498 30098 66510
rect 30046 66434 30098 66446
rect 30382 66498 30434 66510
rect 30382 66434 30434 66446
rect 32958 66498 33010 66510
rect 32958 66434 33010 66446
rect 5070 66386 5122 66398
rect 9998 66386 10050 66398
rect 8642 66334 8654 66386
rect 8706 66334 8718 66386
rect 5070 66322 5122 66334
rect 9998 66322 10050 66334
rect 10894 66386 10946 66398
rect 10894 66322 10946 66334
rect 14814 66386 14866 66398
rect 14814 66322 14866 66334
rect 15598 66386 15650 66398
rect 21422 66386 21474 66398
rect 26014 66386 26066 66398
rect 31166 66386 31218 66398
rect 16594 66334 16606 66386
rect 16658 66334 16670 66386
rect 18722 66334 18734 66386
rect 18786 66334 18798 66386
rect 24882 66334 24894 66386
rect 24946 66334 24958 66386
rect 29698 66334 29710 66386
rect 29762 66334 29774 66386
rect 15598 66322 15650 66334
rect 21422 66322 21474 66334
rect 26014 66322 26066 66334
rect 31166 66322 31218 66334
rect 34638 66386 34690 66398
rect 34638 66322 34690 66334
rect 3726 66274 3778 66286
rect 3726 66210 3778 66222
rect 3950 66274 4002 66286
rect 9102 66274 9154 66286
rect 4498 66222 4510 66274
rect 4562 66222 4574 66274
rect 5842 66222 5854 66274
rect 5906 66222 5918 66274
rect 3950 66210 4002 66222
rect 9102 66210 9154 66222
rect 9326 66274 9378 66286
rect 9326 66210 9378 66222
rect 10222 66274 10274 66286
rect 10222 66210 10274 66222
rect 11118 66274 11170 66286
rect 18174 66274 18226 66286
rect 20638 66274 20690 66286
rect 29486 66274 29538 66286
rect 33294 66274 33346 66286
rect 37326 66274 37378 66286
rect 16482 66222 16494 66274
rect 16546 66222 16558 66274
rect 17714 66222 17726 66274
rect 17778 66222 17790 66274
rect 17938 66222 17950 66274
rect 18002 66222 18014 66274
rect 18946 66222 18958 66274
rect 19010 66222 19022 66274
rect 19394 66222 19406 66274
rect 19458 66222 19470 66274
rect 20402 66222 20414 66274
rect 20466 66222 20478 66274
rect 22082 66222 22094 66274
rect 22146 66222 22158 66274
rect 30370 66222 30382 66274
rect 30434 66222 30446 66274
rect 34850 66222 34862 66274
rect 34914 66222 34926 66274
rect 11118 66210 11170 66222
rect 18174 66210 18226 66222
rect 20638 66210 20690 66222
rect 29486 66210 29538 66222
rect 33294 66210 33346 66222
rect 37326 66210 37378 66222
rect 14254 66162 14306 66174
rect 25230 66162 25282 66174
rect 6514 66110 6526 66162
rect 6578 66110 6590 66162
rect 22754 66110 22766 66162
rect 22818 66110 22830 66162
rect 14254 66098 14306 66110
rect 25230 66098 25282 66110
rect 25566 66162 25618 66174
rect 25566 66098 25618 66110
rect 29822 66162 29874 66174
rect 29822 66098 29874 66110
rect 30718 66162 30770 66174
rect 30718 66098 30770 66110
rect 31838 66162 31890 66174
rect 31838 66098 31890 66110
rect 33518 66162 33570 66174
rect 33518 66098 33570 66110
rect 35422 66162 35474 66174
rect 35422 66098 35474 66110
rect 37550 66162 37602 66174
rect 37550 66098 37602 66110
rect 4286 66050 4338 66062
rect 11902 66050 11954 66062
rect 9650 65998 9662 66050
rect 9714 65998 9726 66050
rect 10546 65998 10558 66050
rect 10610 65998 10622 66050
rect 11442 65998 11454 66050
rect 11506 65998 11518 66050
rect 4286 65986 4338 65998
rect 11902 65986 11954 65998
rect 14142 66050 14194 66062
rect 14142 65986 14194 65998
rect 36318 66050 36370 66062
rect 36978 65998 36990 66050
rect 37042 65998 37054 66050
rect 36318 65986 36370 65998
rect 1344 65882 38640 65916
rect 1344 65830 19838 65882
rect 19890 65830 19942 65882
rect 19994 65830 20046 65882
rect 20098 65830 38640 65882
rect 1344 65796 38640 65830
rect 9886 65714 9938 65726
rect 9886 65650 9938 65662
rect 10782 65714 10834 65726
rect 10782 65650 10834 65662
rect 22654 65714 22706 65726
rect 33294 65714 33346 65726
rect 25778 65662 25790 65714
rect 25842 65662 25854 65714
rect 22654 65650 22706 65662
rect 33294 65650 33346 65662
rect 7086 65602 7138 65614
rect 20526 65602 20578 65614
rect 32398 65602 32450 65614
rect 3602 65550 3614 65602
rect 3666 65550 3678 65602
rect 16258 65550 16270 65602
rect 16322 65550 16334 65602
rect 17490 65550 17502 65602
rect 17554 65550 17566 65602
rect 30930 65550 30942 65602
rect 30994 65550 31006 65602
rect 33842 65550 33854 65602
rect 33906 65550 33918 65602
rect 7086 65538 7138 65550
rect 20526 65538 20578 65550
rect 32398 65538 32450 65550
rect 7422 65490 7474 65502
rect 19070 65490 19122 65502
rect 22318 65490 22370 65502
rect 2930 65438 2942 65490
rect 2994 65438 3006 65490
rect 11778 65438 11790 65490
rect 11842 65438 11854 65490
rect 15026 65438 15038 65490
rect 15090 65438 15102 65490
rect 15586 65438 15598 65490
rect 15650 65438 15662 65490
rect 21186 65438 21198 65490
rect 21250 65438 21262 65490
rect 7422 65426 7474 65438
rect 19070 65426 19122 65438
rect 22318 65426 22370 65438
rect 22990 65490 23042 65502
rect 22990 65426 23042 65438
rect 23214 65490 23266 65502
rect 23214 65426 23266 65438
rect 23438 65490 23490 65502
rect 23438 65426 23490 65438
rect 23886 65490 23938 65502
rect 23886 65426 23938 65438
rect 23998 65490 24050 65502
rect 23998 65426 24050 65438
rect 25230 65490 25282 65502
rect 32174 65490 32226 65502
rect 28802 65438 28814 65490
rect 28866 65438 28878 65490
rect 30034 65438 30046 65490
rect 30098 65438 30110 65490
rect 30594 65438 30606 65490
rect 30658 65438 30670 65490
rect 25230 65426 25282 65438
rect 32174 65426 32226 65438
rect 32510 65490 32562 65502
rect 32510 65426 32562 65438
rect 33406 65490 33458 65502
rect 34178 65438 34190 65490
rect 34242 65438 34254 65490
rect 35186 65438 35198 65490
rect 35250 65438 35262 65490
rect 35858 65438 35870 65490
rect 35922 65438 35934 65490
rect 37426 65438 37438 65490
rect 37490 65438 37502 65490
rect 33406 65426 33458 65438
rect 6190 65378 6242 65390
rect 5730 65326 5742 65378
rect 5794 65326 5806 65378
rect 6190 65314 6242 65326
rect 8878 65378 8930 65390
rect 16046 65378 16098 65390
rect 12450 65326 12462 65378
rect 12514 65326 12526 65378
rect 14578 65326 14590 65378
rect 14642 65326 14654 65378
rect 8878 65314 8930 65326
rect 16046 65314 16098 65326
rect 16718 65378 16770 65390
rect 16718 65314 16770 65326
rect 19182 65378 19234 65390
rect 19182 65314 19234 65326
rect 21870 65378 21922 65390
rect 21870 65314 21922 65326
rect 24222 65378 24274 65390
rect 24222 65314 24274 65326
rect 24670 65378 24722 65390
rect 24670 65314 24722 65326
rect 26238 65378 26290 65390
rect 26238 65314 26290 65326
rect 26686 65378 26738 65390
rect 26686 65314 26738 65326
rect 28590 65378 28642 65390
rect 28590 65314 28642 65326
rect 31614 65378 31666 65390
rect 31614 65314 31666 65326
rect 33518 65378 33570 65390
rect 34514 65326 34526 65378
rect 34578 65326 34590 65378
rect 35970 65326 35982 65378
rect 36034 65326 36046 65378
rect 37762 65326 37774 65378
rect 37826 65326 37838 65378
rect 33518 65314 33570 65326
rect 21758 65266 21810 65278
rect 21758 65202 21810 65214
rect 25454 65266 25506 65278
rect 25454 65202 25506 65214
rect 1344 65098 38640 65132
rect 1344 65046 4478 65098
rect 4530 65046 4582 65098
rect 4634 65046 4686 65098
rect 4738 65046 35198 65098
rect 35250 65046 35302 65098
rect 35354 65046 35406 65098
rect 35458 65046 38640 65098
rect 1344 65012 38640 65046
rect 13470 64930 13522 64942
rect 3826 64878 3838 64930
rect 3890 64878 3902 64930
rect 7858 64878 7870 64930
rect 7922 64878 7934 64930
rect 13470 64866 13522 64878
rect 15038 64930 15090 64942
rect 26350 64930 26402 64942
rect 29598 64930 29650 64942
rect 22978 64878 22990 64930
rect 23042 64878 23054 64930
rect 28578 64878 28590 64930
rect 28642 64878 28654 64930
rect 15038 64866 15090 64878
rect 26350 64866 26402 64878
rect 29598 64866 29650 64878
rect 34974 64930 35026 64942
rect 35522 64878 35534 64930
rect 35586 64878 35598 64930
rect 34974 64866 35026 64878
rect 4174 64818 4226 64830
rect 4174 64754 4226 64766
rect 4398 64818 4450 64830
rect 4398 64754 4450 64766
rect 12462 64818 12514 64830
rect 12462 64754 12514 64766
rect 13022 64818 13074 64830
rect 13022 64754 13074 64766
rect 13582 64818 13634 64830
rect 13582 64754 13634 64766
rect 22094 64818 22146 64830
rect 22094 64754 22146 64766
rect 25118 64818 25170 64830
rect 25118 64754 25170 64766
rect 25454 64818 25506 64830
rect 25454 64754 25506 64766
rect 28030 64818 28082 64830
rect 33618 64766 33630 64818
rect 33682 64766 33694 64818
rect 36306 64766 36318 64818
rect 36370 64766 36382 64818
rect 36978 64766 36990 64818
rect 37042 64766 37054 64818
rect 28030 64754 28082 64766
rect 8206 64706 8258 64718
rect 8206 64642 8258 64654
rect 8430 64706 8482 64718
rect 14366 64706 14418 64718
rect 18622 64706 18674 64718
rect 23326 64706 23378 64718
rect 13794 64654 13806 64706
rect 13858 64654 13870 64706
rect 15026 64654 15038 64706
rect 15090 64654 15102 64706
rect 15474 64654 15486 64706
rect 15538 64654 15550 64706
rect 16034 64654 16046 64706
rect 16098 64654 16110 64706
rect 20738 64654 20750 64706
rect 20802 64654 20814 64706
rect 21298 64654 21310 64706
rect 21362 64654 21374 64706
rect 8430 64642 8482 64654
rect 14366 64642 14418 64654
rect 18622 64642 18674 64654
rect 23326 64642 23378 64654
rect 23550 64706 23602 64718
rect 23550 64642 23602 64654
rect 24110 64706 24162 64718
rect 24110 64642 24162 64654
rect 24334 64706 24386 64718
rect 24334 64642 24386 64654
rect 24894 64706 24946 64718
rect 24894 64642 24946 64654
rect 25678 64706 25730 64718
rect 25678 64642 25730 64654
rect 28254 64706 28306 64718
rect 37886 64706 37938 64718
rect 31154 64654 31166 64706
rect 31218 64654 31230 64706
rect 32610 64654 32622 64706
rect 32674 64654 32686 64706
rect 33394 64654 33406 64706
rect 33458 64654 33470 64706
rect 34066 64654 34078 64706
rect 34130 64654 34142 64706
rect 34626 64654 34638 64706
rect 34690 64654 34702 64706
rect 35858 64654 35870 64706
rect 35922 64654 35934 64706
rect 36082 64654 36094 64706
rect 36146 64654 36158 64706
rect 37090 64654 37102 64706
rect 37154 64654 37166 64706
rect 28254 64642 28306 64654
rect 37886 64642 37938 64654
rect 4846 64594 4898 64606
rect 19518 64594 19570 64606
rect 16146 64542 16158 64594
rect 16210 64542 16222 64594
rect 16930 64542 16942 64594
rect 16994 64542 17006 64594
rect 4846 64530 4898 64542
rect 19518 64530 19570 64542
rect 21646 64594 21698 64606
rect 21646 64530 21698 64542
rect 22542 64594 22594 64606
rect 26462 64594 26514 64606
rect 24658 64542 24670 64594
rect 24722 64542 24734 64594
rect 22542 64530 22594 64542
rect 26462 64530 26514 64542
rect 27806 64594 27858 64606
rect 27806 64530 27858 64542
rect 29262 64594 29314 64606
rect 34414 64594 34466 64606
rect 33058 64542 33070 64594
rect 33122 64542 33134 64594
rect 29262 64530 29314 64542
rect 34414 64530 34466 64542
rect 34862 64594 34914 64606
rect 38222 64594 38274 64606
rect 37314 64542 37326 64594
rect 37378 64542 37390 64594
rect 34862 64530 34914 64542
rect 38222 64530 38274 64542
rect 7534 64482 7586 64494
rect 7534 64418 7586 64430
rect 14030 64482 14082 64494
rect 14030 64418 14082 64430
rect 14254 64482 14306 64494
rect 21534 64482 21586 64494
rect 26910 64482 26962 64494
rect 18498 64430 18510 64482
rect 18562 64430 18574 64482
rect 26002 64430 26014 64482
rect 26066 64430 26078 64482
rect 14254 64418 14306 64430
rect 21534 64418 21586 64430
rect 26910 64418 26962 64430
rect 29486 64482 29538 64494
rect 29486 64418 29538 64430
rect 30046 64482 30098 64494
rect 30046 64418 30098 64430
rect 32062 64482 32114 64494
rect 32062 64418 32114 64430
rect 32174 64482 32226 64494
rect 32174 64418 32226 64430
rect 32286 64482 32338 64494
rect 32286 64418 32338 64430
rect 38110 64482 38162 64494
rect 38110 64418 38162 64430
rect 1344 64314 38640 64348
rect 1344 64262 19838 64314
rect 19890 64262 19942 64314
rect 19994 64262 20046 64314
rect 20098 64262 38640 64314
rect 1344 64228 38640 64262
rect 16830 64146 16882 64158
rect 25342 64146 25394 64158
rect 23202 64094 23214 64146
rect 23266 64094 23278 64146
rect 16830 64082 16882 64094
rect 25342 64082 25394 64094
rect 26238 64146 26290 64158
rect 26238 64082 26290 64094
rect 28702 64146 28754 64158
rect 28702 64082 28754 64094
rect 32062 64146 32114 64158
rect 32062 64082 32114 64094
rect 14590 64034 14642 64046
rect 19966 64034 20018 64046
rect 27134 64034 27186 64046
rect 12114 63982 12126 64034
rect 12178 63982 12190 64034
rect 16370 63982 16382 64034
rect 16434 63982 16446 64034
rect 17490 63982 17502 64034
rect 17554 63982 17566 64034
rect 21858 63982 21870 64034
rect 21922 63982 21934 64034
rect 14590 63970 14642 63982
rect 19966 63970 20018 63982
rect 27134 63970 27186 63982
rect 29150 64034 29202 64046
rect 29150 63970 29202 63982
rect 29262 64034 29314 64046
rect 29262 63970 29314 63982
rect 30382 64034 30434 64046
rect 31950 64034 32002 64046
rect 30930 63982 30942 64034
rect 30994 63982 31006 64034
rect 30382 63970 30434 63982
rect 31950 63970 32002 63982
rect 32286 64034 32338 64046
rect 32286 63970 32338 63982
rect 32510 64034 32562 64046
rect 33506 63982 33518 64034
rect 33570 63982 33582 64034
rect 34626 63982 34638 64034
rect 34690 63982 34702 64034
rect 36082 63982 36094 64034
rect 36146 63982 36158 64034
rect 37426 63982 37438 64034
rect 37490 63982 37502 64034
rect 32510 63970 32562 63982
rect 23550 63922 23602 63934
rect 11442 63870 11454 63922
rect 11506 63870 11518 63922
rect 15138 63870 15150 63922
rect 15202 63870 15214 63922
rect 15698 63870 15710 63922
rect 15762 63870 15774 63922
rect 16258 63870 16270 63922
rect 16322 63870 16334 63922
rect 17378 63870 17390 63922
rect 17442 63870 17454 63922
rect 21186 63870 21198 63922
rect 21250 63870 21262 63922
rect 22978 63870 22990 63922
rect 23042 63870 23054 63922
rect 23550 63858 23602 63870
rect 23774 63922 23826 63934
rect 23774 63858 23826 63870
rect 24222 63922 24274 63934
rect 24222 63858 24274 63870
rect 24334 63922 24386 63934
rect 24334 63858 24386 63870
rect 24558 63922 24610 63934
rect 24558 63858 24610 63870
rect 25790 63922 25842 63934
rect 25790 63858 25842 63870
rect 27806 63922 27858 63934
rect 27806 63858 27858 63870
rect 28590 63922 28642 63934
rect 28590 63858 28642 63870
rect 28926 63922 28978 63934
rect 28926 63858 28978 63870
rect 29486 63922 29538 63934
rect 29922 63870 29934 63922
rect 29986 63870 29998 63922
rect 30818 63870 30830 63922
rect 30882 63870 30894 63922
rect 33842 63870 33854 63922
rect 33906 63870 33918 63922
rect 35074 63870 35086 63922
rect 35138 63870 35150 63922
rect 36306 63870 36318 63922
rect 36370 63870 36382 63922
rect 38210 63870 38222 63922
rect 38274 63870 38286 63922
rect 29486 63858 29538 63870
rect 26686 63810 26738 63822
rect 14242 63758 14254 63810
rect 14306 63758 14318 63810
rect 19618 63758 19630 63810
rect 19682 63758 19694 63810
rect 26686 63746 26738 63758
rect 28254 63810 28306 63822
rect 31266 63758 31278 63810
rect 31330 63758 31342 63810
rect 28254 63746 28306 63758
rect 14702 63698 14754 63710
rect 14702 63634 14754 63646
rect 1344 63530 38640 63564
rect 1344 63478 4478 63530
rect 4530 63478 4582 63530
rect 4634 63478 4686 63530
rect 4738 63478 35198 63530
rect 35250 63478 35302 63530
rect 35354 63478 35406 63530
rect 35458 63478 38640 63530
rect 1344 63444 38640 63478
rect 14018 63310 14030 63362
rect 14082 63310 14094 63362
rect 15138 63310 15150 63362
rect 15202 63310 15214 63362
rect 30706 63310 30718 63362
rect 30770 63310 30782 63362
rect 33394 63310 33406 63362
rect 33458 63310 33470 63362
rect 37538 63310 37550 63362
rect 37602 63310 37614 63362
rect 13470 63250 13522 63262
rect 11890 63198 11902 63250
rect 11954 63198 11966 63250
rect 18610 63198 18622 63250
rect 18674 63198 18686 63250
rect 20738 63198 20750 63250
rect 20802 63198 20814 63250
rect 27346 63198 27358 63250
rect 27410 63198 27422 63250
rect 35970 63198 35982 63250
rect 36034 63198 36046 63250
rect 13470 63186 13522 63198
rect 13694 63138 13746 63150
rect 21422 63138 21474 63150
rect 8978 63086 8990 63138
rect 9042 63086 9054 63138
rect 15026 63086 15038 63138
rect 15090 63086 15102 63138
rect 15474 63086 15486 63138
rect 15538 63086 15550 63138
rect 16034 63086 16046 63138
rect 16098 63086 16110 63138
rect 17938 63086 17950 63138
rect 18002 63086 18014 63138
rect 13694 63074 13746 63086
rect 21422 63074 21474 63086
rect 23102 63138 23154 63150
rect 27806 63138 27858 63150
rect 30606 63138 30658 63150
rect 24546 63086 24558 63138
rect 24610 63086 24622 63138
rect 29922 63086 29934 63138
rect 29986 63086 29998 63138
rect 30818 63086 30830 63138
rect 30882 63086 30894 63138
rect 32162 63086 32174 63138
rect 32226 63086 32238 63138
rect 33506 63086 33518 63138
rect 33570 63086 33582 63138
rect 33842 63086 33854 63138
rect 33906 63086 33918 63138
rect 35522 63086 35534 63138
rect 35586 63086 35598 63138
rect 36082 63086 36094 63138
rect 36146 63086 36158 63138
rect 37538 63086 37550 63138
rect 37602 63086 37614 63138
rect 37874 63086 37886 63138
rect 37938 63086 37950 63138
rect 23102 63074 23154 63086
rect 27806 63074 27858 63086
rect 30606 63074 30658 63086
rect 6414 63026 6466 63038
rect 14478 63026 14530 63038
rect 16606 63026 16658 63038
rect 9762 62974 9774 63026
rect 9826 62974 9838 63026
rect 16146 62974 16158 63026
rect 16210 62974 16222 63026
rect 6414 62962 6466 62974
rect 14478 62962 14530 62974
rect 16606 62962 16658 62974
rect 17278 63026 17330 63038
rect 17278 62962 17330 62974
rect 21870 63026 21922 63038
rect 29262 63026 29314 63038
rect 25218 62974 25230 63026
rect 25282 62974 25294 63026
rect 21870 62962 21922 62974
rect 29262 62962 29314 62974
rect 29598 63026 29650 63038
rect 29598 62962 29650 62974
rect 35198 63026 35250 63038
rect 36418 62974 36430 63026
rect 36482 62974 36494 63026
rect 35198 62962 35250 62974
rect 6750 62914 6802 62926
rect 6750 62850 6802 62862
rect 12350 62914 12402 62926
rect 12350 62850 12402 62862
rect 16494 62914 16546 62926
rect 16494 62850 16546 62862
rect 16830 62914 16882 62926
rect 16830 62850 16882 62862
rect 17054 62914 17106 62926
rect 17054 62850 17106 62862
rect 21422 62914 21474 62926
rect 21422 62850 21474 62862
rect 1344 62746 38640 62780
rect 1344 62694 19838 62746
rect 19890 62694 19942 62746
rect 19994 62694 20046 62746
rect 20098 62694 38640 62746
rect 1344 62660 38640 62694
rect 9662 62578 9714 62590
rect 9662 62514 9714 62526
rect 9998 62578 10050 62590
rect 9998 62514 10050 62526
rect 14254 62578 14306 62590
rect 14254 62514 14306 62526
rect 14702 62578 14754 62590
rect 14702 62514 14754 62526
rect 16830 62578 16882 62590
rect 16830 62514 16882 62526
rect 18174 62578 18226 62590
rect 18174 62514 18226 62526
rect 18622 62578 18674 62590
rect 18622 62514 18674 62526
rect 19070 62578 19122 62590
rect 19070 62514 19122 62526
rect 23102 62578 23154 62590
rect 30494 62578 30546 62590
rect 29810 62526 29822 62578
rect 29874 62526 29886 62578
rect 23102 62514 23154 62526
rect 30494 62514 30546 62526
rect 37998 62578 38050 62590
rect 37998 62514 38050 62526
rect 25902 62466 25954 62478
rect 32622 62466 32674 62478
rect 6514 62414 6526 62466
rect 6578 62414 6590 62466
rect 20066 62414 20078 62466
rect 20130 62414 20142 62466
rect 21186 62414 21198 62466
rect 21250 62414 21262 62466
rect 31714 62414 31726 62466
rect 31778 62414 31790 62466
rect 32274 62414 32286 62466
rect 32338 62414 32350 62466
rect 25902 62402 25954 62414
rect 32622 62402 32674 62414
rect 10334 62354 10386 62366
rect 29486 62354 29538 62366
rect 1698 62302 1710 62354
rect 1762 62302 1774 62354
rect 5730 62302 5742 62354
rect 5794 62302 5806 62354
rect 15362 62302 15374 62354
rect 15426 62302 15438 62354
rect 16482 62302 16494 62354
rect 16546 62302 16558 62354
rect 19394 62302 19406 62354
rect 19458 62302 19470 62354
rect 21074 62302 21086 62354
rect 21138 62302 21150 62354
rect 22978 62302 22990 62354
rect 23042 62302 23054 62354
rect 25666 62302 25678 62354
rect 25730 62302 25742 62354
rect 10334 62290 10386 62302
rect 29486 62290 29538 62302
rect 32510 62354 32562 62366
rect 33618 62302 33630 62354
rect 33682 62302 33694 62354
rect 34738 62302 34750 62354
rect 34802 62302 34814 62354
rect 35074 62302 35086 62354
rect 35138 62302 35150 62354
rect 36418 62302 36430 62354
rect 36482 62302 36494 62354
rect 36642 62302 36654 62354
rect 36706 62302 36718 62354
rect 32510 62290 32562 62302
rect 5070 62242 5122 62254
rect 17726 62242 17778 62254
rect 2482 62190 2494 62242
rect 2546 62190 2558 62242
rect 4610 62190 4622 62242
rect 4674 62190 4686 62242
rect 8642 62190 8654 62242
rect 8706 62190 8718 62242
rect 15810 62190 15822 62242
rect 15874 62190 15886 62242
rect 5070 62178 5122 62190
rect 17726 62178 17778 62190
rect 29038 62242 29090 62254
rect 29038 62178 29090 62190
rect 29262 62242 29314 62254
rect 29262 62178 29314 62190
rect 31054 62242 31106 62254
rect 31054 62178 31106 62190
rect 38110 62242 38162 62254
rect 38110 62178 38162 62190
rect 16270 62130 16322 62142
rect 16270 62066 16322 62078
rect 19518 62130 19570 62142
rect 34402 62078 34414 62130
rect 34466 62078 34478 62130
rect 19518 62066 19570 62078
rect 1344 61962 38640 61996
rect 1344 61910 4478 61962
rect 4530 61910 4582 61962
rect 4634 61910 4686 61962
rect 4738 61910 35198 61962
rect 35250 61910 35302 61962
rect 35354 61910 35406 61962
rect 35458 61910 38640 61962
rect 1344 61876 38640 61910
rect 6190 61794 6242 61806
rect 6190 61730 6242 61742
rect 14030 61794 14082 61806
rect 16146 61742 16158 61794
rect 16210 61791 16222 61794
rect 16706 61791 16718 61794
rect 16210 61745 16718 61791
rect 16210 61742 16222 61745
rect 16706 61742 16718 61745
rect 16770 61742 16782 61794
rect 27570 61742 27582 61794
rect 27634 61791 27646 61794
rect 27794 61791 27806 61794
rect 27634 61745 27806 61791
rect 27634 61742 27646 61745
rect 27794 61742 27806 61745
rect 27858 61742 27870 61794
rect 29698 61742 29710 61794
rect 29762 61742 29774 61794
rect 14030 61730 14082 61742
rect 5966 61682 6018 61694
rect 5966 61618 6018 61630
rect 6526 61682 6578 61694
rect 6526 61618 6578 61630
rect 9998 61682 10050 61694
rect 9998 61618 10050 61630
rect 16158 61682 16210 61694
rect 16158 61618 16210 61630
rect 17726 61682 17778 61694
rect 17726 61618 17778 61630
rect 20750 61682 20802 61694
rect 20750 61618 20802 61630
rect 21422 61682 21474 61694
rect 27806 61682 27858 61694
rect 24434 61630 24446 61682
rect 24498 61630 24510 61682
rect 26562 61630 26574 61682
rect 26626 61630 26638 61682
rect 29362 61630 29374 61682
rect 29426 61630 29438 61682
rect 35746 61630 35758 61682
rect 35810 61630 35822 61682
rect 37762 61630 37774 61682
rect 37826 61630 37838 61682
rect 21422 61618 21474 61630
rect 27806 61618 27858 61630
rect 15150 61570 15202 61582
rect 15150 61506 15202 61518
rect 20190 61570 20242 61582
rect 36990 61570 37042 61582
rect 21746 61518 21758 61570
rect 21810 61518 21822 61570
rect 27346 61518 27358 61570
rect 27410 61518 27422 61570
rect 29474 61518 29486 61570
rect 29538 61518 29550 61570
rect 30482 61518 30494 61570
rect 30546 61518 30558 61570
rect 31826 61518 31838 61570
rect 31890 61518 31902 61570
rect 32274 61518 32286 61570
rect 32338 61518 32350 61570
rect 33170 61518 33182 61570
rect 33234 61518 33246 61570
rect 33618 61518 33630 61570
rect 33682 61518 33694 61570
rect 34402 61518 34414 61570
rect 34466 61518 34478 61570
rect 35410 61518 35422 61570
rect 35474 61518 35486 61570
rect 20190 61506 20242 61518
rect 36990 61506 37042 61518
rect 2830 61458 2882 61470
rect 2830 61394 2882 61406
rect 3166 61458 3218 61470
rect 3166 61394 3218 61406
rect 6750 61458 6802 61470
rect 6750 61394 6802 61406
rect 13918 61458 13970 61470
rect 13918 61394 13970 61406
rect 14590 61458 14642 61470
rect 14590 61394 14642 61406
rect 14702 61458 14754 61470
rect 14702 61394 14754 61406
rect 17054 61458 17106 61470
rect 30942 61458 30994 61470
rect 37214 61458 37266 61470
rect 20290 61406 20302 61458
rect 20354 61455 20366 61458
rect 20514 61455 20526 61458
rect 20354 61409 20526 61455
rect 20354 61406 20366 61409
rect 20514 61406 20526 61409
rect 20578 61406 20590 61458
rect 23090 61406 23102 61458
rect 23154 61406 23166 61458
rect 31714 61406 31726 61458
rect 31778 61406 31790 61458
rect 33282 61406 33294 61458
rect 33346 61406 33358 61458
rect 36194 61406 36206 61458
rect 36258 61406 36270 61458
rect 17054 61394 17106 61406
rect 30942 61394 30994 61406
rect 37214 61394 37266 61406
rect 37438 61458 37490 61470
rect 37438 61394 37490 61406
rect 4174 61346 4226 61358
rect 4174 61282 4226 61294
rect 7646 61346 7698 61358
rect 7646 61282 7698 61294
rect 8094 61346 8146 61358
rect 8094 61282 8146 61294
rect 9102 61346 9154 61358
rect 9102 61282 9154 61294
rect 14366 61346 14418 61358
rect 14366 61282 14418 61294
rect 16606 61346 16658 61358
rect 16606 61282 16658 61294
rect 20078 61346 20130 61358
rect 20078 61282 20130 61294
rect 23886 61346 23938 61358
rect 23886 61282 23938 61294
rect 28590 61346 28642 61358
rect 31938 61294 31950 61346
rect 32002 61294 32014 61346
rect 28590 61282 28642 61294
rect 1344 61178 38640 61212
rect 1344 61126 19838 61178
rect 19890 61126 19942 61178
rect 19994 61126 20046 61178
rect 20098 61126 38640 61178
rect 1344 61092 38640 61126
rect 7982 61010 8034 61022
rect 18958 61010 19010 61022
rect 3378 60958 3390 61010
rect 3442 60958 3454 61010
rect 10322 60958 10334 61010
rect 10386 60958 10398 61010
rect 7982 60946 8034 60958
rect 18958 60946 19010 60958
rect 23214 61010 23266 61022
rect 23214 60946 23266 60958
rect 23662 61010 23714 61022
rect 23662 60946 23714 60958
rect 25342 61010 25394 61022
rect 25342 60946 25394 60958
rect 32286 61010 32338 61022
rect 32286 60946 32338 60958
rect 32398 61010 32450 61022
rect 32398 60946 32450 60958
rect 6862 60898 6914 60910
rect 9550 60898 9602 60910
rect 5730 60846 5742 60898
rect 5794 60846 5806 60898
rect 7410 60846 7422 60898
rect 7474 60846 7486 60898
rect 6862 60834 6914 60846
rect 9550 60834 9602 60846
rect 19406 60898 19458 60910
rect 19406 60834 19458 60846
rect 19518 60898 19570 60910
rect 28254 60898 28306 60910
rect 21410 60846 21422 60898
rect 21474 60846 21486 60898
rect 19518 60834 19570 60846
rect 4286 60786 4338 60798
rect 9886 60786 9938 60798
rect 6178 60734 6190 60786
rect 6242 60734 6254 60786
rect 6962 60734 6974 60786
rect 7026 60734 7038 60786
rect 4286 60722 4338 60734
rect 9886 60722 9938 60734
rect 10670 60786 10722 60798
rect 10670 60722 10722 60734
rect 19182 60786 19234 60798
rect 19182 60722 19234 60734
rect 21198 60786 21250 60798
rect 21198 60722 21250 60734
rect 3950 60674 4002 60686
rect 3950 60610 4002 60622
rect 5294 60674 5346 60686
rect 10894 60674 10946 60686
rect 6290 60622 6302 60674
rect 6354 60622 6366 60674
rect 5294 60610 5346 60622
rect 10894 60610 10946 60622
rect 11454 60674 11506 60686
rect 11454 60610 11506 60622
rect 20302 60674 20354 60686
rect 20302 60610 20354 60622
rect 20750 60674 20802 60686
rect 20750 60610 20802 60622
rect 3726 60562 3778 60574
rect 3726 60498 3778 60510
rect 4510 60562 4562 60574
rect 4834 60510 4846 60562
rect 4898 60510 4910 60562
rect 11106 60510 11118 60562
rect 11170 60559 11182 60562
rect 11442 60559 11454 60562
rect 11170 60513 11454 60559
rect 11170 60510 11182 60513
rect 11442 60510 11454 60513
rect 11506 60510 11518 60562
rect 20290 60510 20302 60562
rect 20354 60559 20366 60562
rect 20514 60559 20526 60562
rect 20354 60513 20526 60559
rect 20354 60510 20366 60513
rect 20514 60510 20526 60513
rect 20578 60559 20590 60562
rect 21425 60559 21471 60846
rect 28254 60834 28306 60846
rect 28366 60898 28418 60910
rect 28366 60834 28418 60846
rect 32510 60898 32562 60910
rect 33730 60846 33742 60898
rect 33794 60846 33806 60898
rect 34850 60846 34862 60898
rect 34914 60846 34926 60898
rect 32510 60834 32562 60846
rect 22766 60786 22818 60798
rect 27470 60786 27522 60798
rect 25554 60734 25566 60786
rect 25618 60734 25630 60786
rect 22766 60722 22818 60734
rect 27470 60722 27522 60734
rect 27918 60786 27970 60798
rect 29138 60734 29150 60786
rect 29202 60734 29214 60786
rect 29586 60734 29598 60786
rect 29650 60734 29662 60786
rect 30482 60734 30494 60786
rect 30546 60734 30558 60786
rect 30818 60734 30830 60786
rect 30882 60734 30894 60786
rect 33058 60734 33070 60786
rect 33122 60734 33134 60786
rect 34178 60734 34190 60786
rect 34242 60734 34254 60786
rect 35298 60734 35310 60786
rect 35362 60734 35374 60786
rect 36418 60734 36430 60786
rect 36482 60734 36494 60786
rect 37650 60734 37662 60786
rect 37714 60734 37726 60786
rect 27918 60722 27970 60734
rect 21646 60674 21698 60686
rect 31490 60622 31502 60674
rect 31554 60622 31566 60674
rect 33506 60622 33518 60674
rect 33570 60622 33582 60674
rect 35970 60622 35982 60674
rect 36034 60622 36046 60674
rect 21646 60610 21698 60622
rect 20578 60513 21471 60559
rect 28366 60562 28418 60574
rect 20578 60510 20590 60513
rect 4510 60498 4562 60510
rect 28366 60498 28418 60510
rect 28814 60562 28866 60574
rect 28814 60498 28866 60510
rect 29150 60562 29202 60574
rect 29150 60498 29202 60510
rect 1344 60394 38640 60428
rect 1344 60342 4478 60394
rect 4530 60342 4582 60394
rect 4634 60342 4686 60394
rect 4738 60342 35198 60394
rect 35250 60342 35302 60394
rect 35354 60342 35406 60394
rect 35458 60342 38640 60394
rect 1344 60308 38640 60342
rect 25342 60226 25394 60238
rect 19058 60174 19070 60226
rect 19122 60174 19134 60226
rect 24658 60174 24670 60226
rect 24722 60223 24734 60226
rect 24994 60223 25006 60226
rect 24722 60177 25006 60223
rect 24722 60174 24734 60177
rect 24994 60174 25006 60177
rect 25058 60174 25070 60226
rect 25342 60162 25394 60174
rect 29598 60226 29650 60238
rect 29598 60162 29650 60174
rect 33070 60226 33122 60238
rect 37538 60174 37550 60226
rect 37602 60174 37614 60226
rect 33070 60162 33122 60174
rect 6974 60114 7026 60126
rect 12462 60114 12514 60126
rect 24222 60114 24274 60126
rect 4610 60062 4622 60114
rect 4674 60062 4686 60114
rect 9090 60062 9102 60114
rect 9154 60062 9166 60114
rect 14242 60062 14254 60114
rect 14306 60062 14318 60114
rect 16370 60062 16382 60114
rect 16434 60062 16446 60114
rect 18722 60062 18734 60114
rect 18786 60062 18798 60114
rect 21634 60062 21646 60114
rect 21698 60062 21710 60114
rect 22418 60062 22430 60114
rect 22482 60062 22494 60114
rect 6974 60050 7026 60062
rect 12462 60050 12514 60062
rect 24222 60050 24274 60062
rect 24670 60114 24722 60126
rect 34638 60114 34690 60126
rect 32050 60062 32062 60114
rect 32114 60062 32126 60114
rect 24670 60050 24722 60062
rect 34638 60050 34690 60062
rect 37662 60114 37714 60126
rect 37662 60050 37714 60062
rect 20638 60002 20690 60014
rect 23886 60002 23938 60014
rect 1810 59950 1822 60002
rect 1874 59950 1886 60002
rect 5842 59950 5854 60002
rect 5906 59950 5918 60002
rect 7746 59950 7758 60002
rect 7810 59950 7822 60002
rect 8418 59950 8430 60002
rect 8482 59950 8494 60002
rect 12002 59950 12014 60002
rect 12066 59950 12078 60002
rect 13458 59950 13470 60002
rect 13522 59950 13534 60002
rect 18946 59950 18958 60002
rect 19010 59950 19022 60002
rect 19394 59950 19406 60002
rect 19458 59950 19470 60002
rect 20402 59950 20414 60002
rect 20466 59950 20478 60002
rect 21970 59950 21982 60002
rect 22034 59950 22046 60002
rect 23650 59950 23662 60002
rect 23714 59950 23726 60002
rect 20638 59938 20690 59950
rect 23886 59938 23938 59950
rect 25678 60002 25730 60014
rect 25678 59938 25730 59950
rect 26350 60002 26402 60014
rect 29586 59950 29598 60002
rect 29650 59950 29662 60002
rect 29922 59950 29934 60002
rect 29986 59950 29998 60002
rect 31266 59950 31278 60002
rect 31330 59950 31342 60002
rect 34850 59950 34862 60002
rect 34914 59950 34926 60002
rect 37874 59950 37886 60002
rect 37938 59950 37950 60002
rect 26350 59938 26402 59950
rect 21310 59890 21362 59902
rect 2482 59838 2494 59890
rect 2546 59838 2558 59890
rect 8530 59838 8542 59890
rect 8594 59838 8606 59890
rect 11218 59838 11230 59890
rect 11282 59838 11294 59890
rect 21310 59826 21362 59838
rect 21534 59890 21586 59902
rect 25902 59890 25954 59902
rect 24098 59838 24110 59890
rect 24162 59838 24174 59890
rect 21534 59826 21586 59838
rect 25902 59826 25954 59838
rect 27694 59890 27746 59902
rect 27694 59826 27746 59838
rect 29262 59890 29314 59902
rect 32846 59890 32898 59902
rect 31826 59838 31838 59890
rect 31890 59838 31902 59890
rect 29262 59826 29314 59838
rect 32846 59826 32898 59838
rect 35870 59890 35922 59902
rect 35870 59826 35922 59838
rect 5070 59778 5122 59790
rect 5070 59714 5122 59726
rect 5630 59778 5682 59790
rect 5630 59714 5682 59726
rect 7534 59778 7586 59790
rect 16830 59778 16882 59790
rect 7634 59726 7646 59778
rect 7698 59726 7710 59778
rect 7534 59714 7586 59726
rect 16830 59714 16882 59726
rect 18174 59778 18226 59790
rect 18174 59714 18226 59726
rect 23214 59778 23266 59790
rect 23214 59714 23266 59726
rect 28254 59778 28306 59790
rect 28254 59714 28306 59726
rect 28702 59778 28754 59790
rect 36318 59778 36370 59790
rect 33394 59726 33406 59778
rect 33458 59726 33470 59778
rect 28702 59714 28754 59726
rect 36318 59714 36370 59726
rect 1344 59610 38640 59644
rect 1344 59558 19838 59610
rect 19890 59558 19942 59610
rect 19994 59558 20046 59610
rect 20098 59558 38640 59610
rect 1344 59524 38640 59558
rect 8990 59442 9042 59454
rect 14254 59442 14306 59454
rect 10098 59390 10110 59442
rect 10162 59390 10174 59442
rect 8990 59378 9042 59390
rect 14254 59378 14306 59390
rect 18734 59442 18786 59454
rect 18734 59378 18786 59390
rect 25454 59442 25506 59454
rect 25454 59378 25506 59390
rect 29822 59442 29874 59454
rect 29822 59378 29874 59390
rect 37662 59442 37714 59454
rect 37662 59378 37714 59390
rect 37886 59442 37938 59454
rect 37886 59378 37938 59390
rect 9550 59330 9602 59342
rect 4610 59278 4622 59330
rect 4674 59278 4686 59330
rect 9550 59266 9602 59278
rect 15486 59330 15538 59342
rect 15486 59266 15538 59278
rect 17502 59330 17554 59342
rect 17502 59266 17554 59278
rect 19518 59330 19570 59342
rect 19518 59266 19570 59278
rect 21534 59330 21586 59342
rect 30942 59330 30994 59342
rect 32398 59330 32450 59342
rect 37998 59330 38050 59342
rect 27906 59278 27918 59330
rect 27970 59278 27982 59330
rect 31602 59278 31614 59330
rect 31666 59278 31678 59330
rect 36306 59278 36318 59330
rect 36370 59278 36382 59330
rect 21534 59266 21586 59278
rect 30942 59266 30994 59278
rect 32398 59266 32450 59278
rect 37998 59266 38050 59278
rect 9774 59218 9826 59230
rect 14590 59218 14642 59230
rect 17390 59218 17442 59230
rect 3826 59166 3838 59218
rect 3890 59166 3902 59218
rect 10882 59166 10894 59218
rect 10946 59166 10958 59218
rect 15698 59166 15710 59218
rect 15762 59166 15774 59218
rect 9774 59154 9826 59166
rect 14590 59154 14642 59166
rect 17390 59154 17442 59166
rect 17614 59218 17666 59230
rect 17614 59154 17666 59166
rect 18062 59218 18114 59230
rect 24446 59218 24498 59230
rect 18946 59166 18958 59218
rect 19010 59166 19022 59218
rect 22754 59166 22766 59218
rect 22818 59166 22830 59218
rect 18062 59154 18114 59166
rect 24446 59154 24498 59166
rect 24670 59218 24722 59230
rect 27570 59166 27582 59218
rect 27634 59166 27646 59218
rect 29698 59166 29710 59218
rect 29762 59166 29774 59218
rect 30482 59166 30494 59218
rect 30546 59166 30558 59218
rect 31714 59166 31726 59218
rect 31778 59166 31790 59218
rect 33282 59166 33294 59218
rect 33346 59166 33358 59218
rect 35298 59166 35310 59218
rect 35362 59166 35374 59218
rect 36194 59166 36206 59218
rect 36258 59166 36270 59218
rect 36418 59166 36430 59218
rect 36482 59166 36494 59218
rect 37090 59166 37102 59218
rect 37154 59166 37166 59218
rect 24670 59154 24722 59166
rect 7198 59106 7250 59118
rect 6738 59054 6750 59106
rect 6802 59054 6814 59106
rect 7198 59042 7250 59054
rect 7646 59106 7698 59118
rect 7646 59042 7698 59054
rect 8542 59106 8594 59118
rect 16382 59106 16434 59118
rect 11666 59054 11678 59106
rect 11730 59054 11742 59106
rect 13794 59054 13806 59106
rect 13858 59054 13870 59106
rect 15138 59054 15150 59106
rect 15202 59054 15214 59106
rect 8542 59042 8594 59054
rect 16382 59042 16434 59054
rect 16830 59106 16882 59118
rect 23214 59106 23266 59118
rect 20962 59054 20974 59106
rect 21026 59054 21038 59106
rect 16830 59042 16882 59054
rect 23214 59042 23266 59054
rect 23774 59106 23826 59118
rect 23774 59042 23826 59054
rect 27358 59106 27410 59118
rect 31266 59054 31278 59106
rect 31330 59054 31342 59106
rect 33506 59054 33518 59106
rect 33570 59054 33582 59106
rect 27358 59042 27410 59054
rect 14814 58994 14866 59006
rect 32510 58994 32562 59006
rect 6962 58942 6974 58994
rect 7026 58991 7038 58994
rect 7522 58991 7534 58994
rect 7026 58945 7534 58991
rect 7026 58942 7038 58945
rect 7522 58942 7534 58945
rect 7586 58942 7598 58994
rect 24098 58942 24110 58994
rect 24162 58942 24174 58994
rect 34178 58942 34190 58994
rect 34242 58942 34254 58994
rect 14814 58930 14866 58942
rect 32510 58930 32562 58942
rect 1344 58826 38640 58860
rect 1344 58774 4478 58826
rect 4530 58774 4582 58826
rect 4634 58774 4686 58826
rect 4738 58774 35198 58826
rect 35250 58774 35302 58826
rect 35354 58774 35406 58826
rect 35458 58774 38640 58826
rect 1344 58740 38640 58774
rect 29486 58658 29538 58670
rect 7970 58655 7982 58658
rect 7649 58609 7982 58655
rect 7298 58494 7310 58546
rect 7362 58494 7374 58546
rect 4846 58434 4898 58446
rect 6862 58434 6914 58446
rect 4386 58382 4398 58434
rect 4450 58382 4462 58434
rect 5058 58382 5070 58434
rect 5122 58382 5134 58434
rect 4846 58370 4898 58382
rect 6862 58370 6914 58382
rect 7198 58434 7250 58446
rect 7198 58370 7250 58382
rect 7310 58322 7362 58334
rect 7522 58270 7534 58322
rect 7586 58319 7598 58322
rect 7649 58319 7695 58609
rect 7970 58606 7982 58609
rect 8034 58606 8046 58658
rect 27794 58606 27806 58658
rect 27858 58655 27870 58658
rect 28130 58655 28142 58658
rect 27858 58609 28142 58655
rect 27858 58606 27870 58609
rect 28130 58606 28142 58609
rect 28194 58655 28206 58658
rect 28466 58655 28478 58658
rect 28194 58609 28478 58655
rect 28194 58606 28206 58609
rect 28466 58606 28478 58609
rect 28530 58606 28542 58658
rect 29486 58594 29538 58606
rect 13582 58546 13634 58558
rect 28478 58546 28530 58558
rect 9090 58494 9102 58546
rect 9154 58494 9166 58546
rect 11218 58494 11230 58546
rect 11282 58494 11294 58546
rect 14690 58494 14702 58546
rect 14754 58494 14766 58546
rect 16818 58494 16830 58546
rect 16882 58494 16894 58546
rect 18610 58494 18622 58546
rect 18674 58494 18686 58546
rect 20738 58494 20750 58546
rect 20802 58494 20814 58546
rect 22082 58494 22094 58546
rect 22146 58494 22158 58546
rect 24210 58494 24222 58546
rect 24274 58494 24286 58546
rect 30258 58494 30270 58546
rect 30322 58494 30334 58546
rect 32722 58494 32734 58546
rect 32786 58494 32798 58546
rect 34850 58494 34862 58546
rect 34914 58494 34926 58546
rect 37426 58494 37438 58546
rect 37490 58494 37502 58546
rect 13582 58482 13634 58494
rect 28478 58482 28530 58494
rect 24670 58434 24722 58446
rect 8418 58382 8430 58434
rect 8482 58382 8494 58434
rect 14018 58382 14030 58434
rect 14082 58382 14094 58434
rect 17826 58382 17838 58434
rect 17890 58382 17902 58434
rect 21410 58382 21422 58434
rect 21474 58382 21486 58434
rect 24670 58370 24722 58382
rect 29374 58434 29426 58446
rect 33182 58434 33234 58446
rect 30594 58382 30606 58434
rect 30658 58382 30670 58434
rect 31714 58382 31726 58434
rect 31778 58382 31790 58434
rect 31938 58382 31950 58434
rect 32002 58382 32014 58434
rect 33842 58382 33854 58434
rect 33906 58382 33918 58434
rect 35522 58382 35534 58434
rect 35586 58382 35598 58434
rect 36978 58382 36990 58434
rect 37042 58382 37054 58434
rect 29374 58370 29426 58382
rect 33182 58370 33234 58382
rect 7586 58273 7695 58319
rect 17278 58322 17330 58334
rect 7586 58270 7598 58273
rect 7310 58258 7362 58270
rect 17278 58258 17330 58270
rect 27694 58322 27746 58334
rect 27694 58258 27746 58270
rect 29934 58322 29986 58334
rect 29934 58258 29986 58270
rect 30158 58322 30210 58334
rect 30158 58258 30210 58270
rect 33406 58322 33458 58334
rect 33406 58258 33458 58270
rect 33518 58322 33570 58334
rect 36194 58270 36206 58322
rect 36258 58270 36270 58322
rect 37090 58270 37102 58322
rect 37154 58270 37166 58322
rect 33518 58258 33570 58270
rect 4622 58210 4674 58222
rect 4622 58146 4674 58158
rect 4734 58210 4786 58222
rect 4734 58146 4786 58158
rect 5742 58210 5794 58222
rect 5742 58146 5794 58158
rect 6190 58210 6242 58222
rect 6190 58146 6242 58158
rect 6974 58210 7026 58222
rect 6974 58146 7026 58158
rect 7870 58210 7922 58222
rect 7870 58146 7922 58158
rect 11678 58210 11730 58222
rect 11678 58146 11730 58158
rect 28030 58210 28082 58222
rect 28030 58146 28082 58158
rect 29486 58210 29538 58222
rect 29486 58146 29538 58158
rect 1344 58042 38640 58076
rect 1344 57990 19838 58042
rect 19890 57990 19942 58042
rect 19994 57990 20046 58042
rect 20098 57990 38640 58042
rect 1344 57956 38640 57990
rect 7534 57874 7586 57886
rect 7534 57810 7586 57822
rect 10894 57874 10946 57886
rect 10894 57810 10946 57822
rect 12126 57874 12178 57886
rect 12126 57810 12178 57822
rect 16046 57874 16098 57886
rect 16046 57810 16098 57822
rect 16830 57874 16882 57886
rect 16830 57810 16882 57822
rect 17614 57874 17666 57886
rect 17614 57810 17666 57822
rect 17838 57874 17890 57886
rect 22318 57874 22370 57886
rect 18050 57822 18062 57874
rect 18114 57822 18126 57874
rect 17838 57810 17890 57822
rect 22318 57810 22370 57822
rect 31614 57874 31666 57886
rect 31614 57810 31666 57822
rect 32286 57874 32338 57886
rect 32286 57810 32338 57822
rect 37886 57874 37938 57886
rect 37886 57810 37938 57822
rect 5070 57762 5122 57774
rect 5070 57698 5122 57710
rect 7086 57762 7138 57774
rect 16158 57762 16210 57774
rect 14130 57710 14142 57762
rect 14194 57710 14206 57762
rect 7086 57698 7138 57710
rect 16158 57698 16210 57710
rect 17390 57762 17442 57774
rect 24222 57762 24274 57774
rect 19170 57710 19182 57762
rect 19234 57710 19246 57762
rect 20178 57710 20190 57762
rect 20242 57710 20254 57762
rect 17390 57698 17442 57710
rect 24222 57698 24274 57710
rect 24558 57762 24610 57774
rect 32510 57762 32562 57774
rect 27794 57710 27806 57762
rect 27858 57710 27870 57762
rect 24558 57698 24610 57710
rect 32510 57698 32562 57710
rect 34302 57762 34354 57774
rect 38222 57762 38274 57774
rect 36530 57710 36542 57762
rect 36594 57710 36606 57762
rect 34302 57698 34354 57710
rect 38222 57698 38274 57710
rect 12462 57650 12514 57662
rect 1810 57598 1822 57650
rect 1874 57598 1886 57650
rect 10658 57598 10670 57650
rect 10722 57598 10734 57650
rect 12462 57586 12514 57598
rect 18062 57650 18114 57662
rect 23214 57650 23266 57662
rect 34190 57650 34242 57662
rect 19954 57598 19966 57650
rect 20018 57598 20030 57650
rect 21858 57598 21870 57650
rect 21922 57598 21934 57650
rect 27906 57598 27918 57650
rect 27970 57598 27982 57650
rect 30594 57598 30606 57650
rect 30658 57598 30670 57650
rect 31042 57598 31054 57650
rect 31106 57598 31118 57650
rect 33842 57598 33854 57650
rect 33906 57598 33918 57650
rect 35522 57598 35534 57650
rect 35586 57598 35598 57650
rect 35858 57598 35870 57650
rect 35922 57598 35934 57650
rect 37202 57598 37214 57650
rect 37266 57598 37278 57650
rect 18062 57586 18114 57598
rect 23214 57586 23266 57598
rect 34190 57586 34242 57598
rect 6862 57538 6914 57550
rect 22766 57538 22818 57550
rect 2482 57486 2494 57538
rect 2546 57486 2558 57538
rect 4610 57486 4622 57538
rect 4674 57486 4686 57538
rect 15026 57486 15038 57538
rect 15090 57486 15102 57538
rect 20402 57486 20414 57538
rect 20466 57486 20478 57538
rect 6862 57474 6914 57486
rect 22766 57474 22818 57486
rect 27134 57538 27186 57550
rect 28802 57486 28814 57538
rect 28866 57486 28878 57538
rect 32162 57486 32174 57538
rect 32226 57486 32238 57538
rect 35746 57486 35758 57538
rect 35810 57486 35822 57538
rect 37090 57486 37102 57538
rect 37154 57486 37166 57538
rect 27134 57474 27186 57486
rect 6526 57426 6578 57438
rect 6526 57362 6578 57374
rect 1344 57258 38640 57292
rect 1344 57206 4478 57258
rect 4530 57206 4582 57258
rect 4634 57206 4686 57258
rect 4738 57206 35198 57258
rect 35250 57206 35302 57258
rect 35354 57206 35406 57258
rect 35458 57206 38640 57258
rect 1344 57172 38640 57206
rect 16942 56978 16994 56990
rect 16942 56914 16994 56926
rect 17950 56978 18002 56990
rect 31950 56978 32002 56990
rect 22082 56926 22094 56978
rect 22146 56926 22158 56978
rect 25330 56926 25342 56978
rect 25394 56926 25406 56978
rect 27458 56926 27470 56978
rect 27522 56926 27534 56978
rect 17950 56914 18002 56926
rect 31950 56914 32002 56926
rect 33518 56978 33570 56990
rect 35646 56978 35698 56990
rect 33842 56926 33854 56978
rect 33906 56926 33918 56978
rect 35186 56926 35198 56978
rect 35250 56926 35262 56978
rect 33518 56914 33570 56926
rect 35646 56914 35698 56926
rect 38334 56978 38386 56990
rect 38334 56914 38386 56926
rect 17166 56866 17218 56878
rect 3042 56814 3054 56866
rect 3106 56814 3118 56866
rect 6850 56814 6862 56866
rect 6914 56814 6926 56866
rect 17166 56802 17218 56814
rect 18286 56866 18338 56878
rect 18286 56802 18338 56814
rect 18510 56866 18562 56878
rect 18510 56802 18562 56814
rect 19294 56866 19346 56878
rect 30718 56866 30770 56878
rect 24882 56814 24894 56866
rect 24946 56814 24958 56866
rect 28130 56814 28142 56866
rect 28194 56814 28206 56866
rect 29138 56814 29150 56866
rect 29202 56814 29214 56866
rect 30146 56814 30158 56866
rect 30210 56814 30222 56866
rect 31266 56814 31278 56866
rect 31330 56814 31342 56866
rect 34962 56814 34974 56866
rect 35026 56814 35038 56866
rect 19294 56802 19346 56814
rect 30718 56802 30770 56814
rect 2830 56754 2882 56766
rect 2830 56690 2882 56702
rect 14590 56754 14642 56766
rect 14590 56690 14642 56702
rect 14702 56754 14754 56766
rect 24210 56702 24222 56754
rect 24274 56702 24286 56754
rect 30258 56702 30270 56754
rect 30322 56702 30334 56754
rect 30930 56702 30942 56754
rect 30994 56702 31006 56754
rect 14702 56690 14754 56702
rect 6638 56642 6690 56654
rect 6638 56578 6690 56590
rect 14142 56642 14194 56654
rect 14142 56578 14194 56590
rect 14366 56642 14418 56654
rect 14366 56578 14418 56590
rect 15598 56642 15650 56654
rect 15598 56578 15650 56590
rect 16606 56642 16658 56654
rect 17490 56590 17502 56642
rect 17554 56590 17566 56642
rect 18834 56590 18846 56642
rect 18898 56590 18910 56642
rect 16606 56578 16658 56590
rect 1344 56474 38640 56508
rect 1344 56422 19838 56474
rect 19890 56422 19942 56474
rect 19994 56422 20046 56474
rect 20098 56422 38640 56474
rect 1344 56388 38640 56422
rect 2830 56306 2882 56318
rect 23886 56306 23938 56318
rect 11218 56254 11230 56306
rect 11282 56254 11294 56306
rect 2830 56242 2882 56254
rect 23886 56242 23938 56254
rect 25342 56306 25394 56318
rect 25342 56242 25394 56254
rect 30942 56306 30994 56318
rect 30942 56242 30994 56254
rect 17502 56194 17554 56206
rect 17502 56130 17554 56142
rect 17838 56194 17890 56206
rect 17838 56130 17890 56142
rect 18510 56194 18562 56206
rect 18510 56130 18562 56142
rect 3166 56082 3218 56094
rect 3166 56018 3218 56030
rect 11566 56082 11618 56094
rect 11566 56018 11618 56030
rect 12238 56082 12290 56094
rect 23650 56030 23662 56082
rect 23714 56030 23726 56082
rect 26674 56030 26686 56082
rect 26738 56030 26750 56082
rect 12238 56018 12290 56030
rect 11790 55970 11842 55982
rect 30046 55970 30098 55982
rect 27458 55918 27470 55970
rect 27522 55918 27534 55970
rect 29586 55918 29598 55970
rect 29650 55918 29662 55970
rect 11790 55906 11842 55918
rect 30046 55906 30098 55918
rect 30494 55970 30546 55982
rect 30494 55906 30546 55918
rect 1344 55690 38640 55724
rect 1344 55638 4478 55690
rect 4530 55638 4582 55690
rect 4634 55638 4686 55690
rect 4738 55638 35198 55690
rect 35250 55638 35302 55690
rect 35354 55638 35406 55690
rect 35458 55638 38640 55690
rect 1344 55604 38640 55638
rect 27682 55470 27694 55522
rect 27746 55519 27758 55522
rect 28018 55519 28030 55522
rect 27746 55473 28030 55519
rect 27746 55470 27758 55473
rect 28018 55470 28030 55473
rect 28082 55470 28094 55522
rect 30370 55470 30382 55522
rect 30434 55470 30446 55522
rect 9774 55410 9826 55422
rect 3602 55358 3614 55410
rect 3666 55358 3678 55410
rect 6514 55358 6526 55410
rect 6578 55358 6590 55410
rect 8642 55358 8654 55410
rect 8706 55358 8718 55410
rect 9774 55346 9826 55358
rect 19742 55410 19794 55422
rect 19742 55346 19794 55358
rect 20638 55410 20690 55422
rect 20638 55346 20690 55358
rect 22094 55410 22146 55422
rect 22094 55346 22146 55358
rect 22542 55410 22594 55422
rect 32286 55410 32338 55422
rect 24210 55358 24222 55410
rect 24274 55358 24286 55410
rect 22542 55346 22594 55358
rect 32286 55346 32338 55358
rect 3950 55298 4002 55310
rect 3950 55234 4002 55246
rect 4174 55298 4226 55310
rect 25678 55298 25730 55310
rect 5730 55246 5742 55298
rect 5794 55246 5806 55298
rect 23314 55246 23326 55298
rect 23378 55246 23390 55298
rect 4174 55234 4226 55246
rect 25678 55234 25730 55246
rect 27918 55298 27970 55310
rect 27918 55234 27970 55246
rect 28142 55298 28194 55310
rect 28142 55234 28194 55246
rect 28478 55298 28530 55310
rect 28478 55234 28530 55246
rect 29150 55298 29202 55310
rect 29362 55246 29374 55298
rect 29426 55246 29438 55298
rect 31154 55246 31166 55298
rect 31218 55246 31230 55298
rect 35410 55246 35422 55298
rect 35474 55246 35486 55298
rect 29150 55234 29202 55246
rect 34862 55186 34914 55198
rect 24546 55134 24558 55186
rect 24610 55134 24622 55186
rect 34862 55122 34914 55134
rect 4622 55074 4674 55086
rect 4622 55010 4674 55022
rect 9326 55074 9378 55086
rect 9326 55010 9378 55022
rect 12238 55074 12290 55086
rect 12238 55010 12290 55022
rect 12686 55074 12738 55086
rect 12686 55010 12738 55022
rect 17950 55074 18002 55086
rect 17950 55010 18002 55022
rect 18510 55074 18562 55086
rect 18510 55010 18562 55022
rect 21422 55074 21474 55086
rect 21422 55010 21474 55022
rect 25566 55074 25618 55086
rect 25566 55010 25618 55022
rect 28366 55074 28418 55086
rect 28366 55010 28418 55022
rect 35758 55074 35810 55086
rect 35758 55010 35810 55022
rect 1344 54906 38640 54940
rect 1344 54854 19838 54906
rect 19890 54854 19942 54906
rect 19994 54854 20046 54906
rect 20098 54854 38640 54906
rect 1344 54820 38640 54854
rect 21870 54738 21922 54750
rect 30046 54738 30098 54750
rect 3602 54686 3614 54738
rect 3666 54686 3678 54738
rect 11666 54686 11678 54738
rect 11730 54686 11742 54738
rect 23874 54686 23886 54738
rect 23938 54686 23950 54738
rect 21870 54674 21922 54686
rect 30046 54674 30098 54686
rect 9550 54626 9602 54638
rect 21422 54626 21474 54638
rect 6850 54574 6862 54626
rect 6914 54574 6926 54626
rect 10434 54574 10446 54626
rect 10498 54574 10510 54626
rect 13010 54574 13022 54626
rect 13074 54574 13086 54626
rect 18162 54574 18174 54626
rect 18226 54574 18238 54626
rect 9550 54562 9602 54574
rect 21422 54562 21474 54574
rect 27918 54626 27970 54638
rect 27918 54562 27970 54574
rect 33182 54626 33234 54638
rect 33182 54562 33234 54574
rect 16830 54514 16882 54526
rect 28814 54514 28866 54526
rect 6178 54462 6190 54514
rect 6242 54462 6254 54514
rect 9762 54462 9774 54514
rect 9826 54462 9838 54514
rect 10882 54462 10894 54514
rect 10946 54462 10958 54514
rect 11218 54462 11230 54514
rect 11282 54462 11294 54514
rect 12338 54462 12350 54514
rect 12402 54462 12414 54514
rect 17378 54462 17390 54514
rect 17442 54462 17454 54514
rect 21186 54462 21198 54514
rect 21250 54462 21262 54514
rect 33394 54462 33406 54514
rect 33458 54462 33470 54514
rect 35298 54462 35310 54514
rect 35362 54462 35374 54514
rect 16830 54450 16882 54462
rect 28814 54450 28866 54462
rect 3950 54402 4002 54414
rect 3950 54338 4002 54350
rect 4174 54402 4226 54414
rect 4174 54338 4226 54350
rect 4622 54402 4674 54414
rect 15598 54402 15650 54414
rect 20750 54402 20802 54414
rect 8978 54350 8990 54402
rect 9042 54350 9054 54402
rect 10434 54350 10446 54402
rect 10498 54350 10510 54402
rect 15138 54350 15150 54402
rect 15202 54350 15214 54402
rect 20290 54350 20302 54402
rect 20354 54350 20366 54402
rect 4622 54338 4674 54350
rect 15598 54338 15650 54350
rect 20750 54338 20802 54350
rect 22430 54402 22482 54414
rect 22430 54338 22482 54350
rect 22878 54402 22930 54414
rect 22878 54338 22930 54350
rect 23438 54402 23490 54414
rect 23438 54338 23490 54350
rect 24446 54402 24498 54414
rect 24446 54338 24498 54350
rect 27022 54402 27074 54414
rect 27022 54338 27074 54350
rect 30158 54402 30210 54414
rect 36082 54350 36094 54402
rect 36146 54350 36158 54402
rect 38210 54350 38222 54402
rect 38274 54350 38286 54402
rect 30158 54338 30210 54350
rect 24222 54290 24274 54302
rect 24222 54226 24274 54238
rect 27358 54290 27410 54302
rect 27358 54226 27410 54238
rect 27694 54290 27746 54302
rect 27694 54226 27746 54238
rect 1344 54122 38640 54156
rect 1344 54070 4478 54122
rect 4530 54070 4582 54122
rect 4634 54070 4686 54122
rect 4738 54070 35198 54122
rect 35250 54070 35302 54122
rect 35354 54070 35406 54122
rect 35458 54070 38640 54122
rect 1344 54036 38640 54070
rect 8206 53954 8258 53966
rect 8206 53890 8258 53902
rect 8542 53954 8594 53966
rect 8542 53890 8594 53902
rect 21310 53954 21362 53966
rect 21310 53890 21362 53902
rect 21646 53954 21698 53966
rect 21646 53890 21698 53902
rect 4846 53842 4898 53854
rect 22878 53842 22930 53854
rect 10770 53790 10782 53842
rect 10834 53790 10846 53842
rect 12898 53790 12910 53842
rect 12962 53790 12974 53842
rect 17042 53790 17054 53842
rect 17106 53790 17118 53842
rect 32050 53790 32062 53842
rect 32114 53790 32126 53842
rect 33170 53790 33182 53842
rect 33234 53790 33246 53842
rect 35298 53790 35310 53842
rect 35362 53790 35374 53842
rect 4846 53778 4898 53790
rect 22878 53778 22930 53790
rect 8990 53730 9042 53742
rect 15822 53730 15874 53742
rect 10098 53678 10110 53730
rect 10162 53678 10174 53730
rect 8990 53666 9042 53678
rect 15822 53666 15874 53678
rect 16718 53730 16770 53742
rect 20402 53678 20414 53730
rect 20466 53678 20478 53730
rect 26786 53678 26798 53730
rect 26850 53678 26862 53730
rect 29138 53678 29150 53730
rect 29202 53678 29214 53730
rect 32386 53678 32398 53730
rect 32450 53678 32462 53730
rect 16718 53666 16770 53678
rect 3726 53618 3778 53630
rect 3726 53554 3778 53566
rect 7982 53618 8034 53630
rect 7982 53554 8034 53566
rect 13470 53618 13522 53630
rect 13470 53554 13522 53566
rect 13806 53618 13858 53630
rect 13806 53554 13858 53566
rect 17838 53618 17890 53630
rect 17838 53554 17890 53566
rect 19294 53618 19346 53630
rect 19294 53554 19346 53566
rect 21870 53618 21922 53630
rect 21870 53554 21922 53566
rect 22430 53618 22482 53630
rect 35982 53618 36034 53630
rect 29922 53566 29934 53618
rect 29986 53566 29998 53618
rect 22430 53554 22482 53566
rect 35982 53554 36034 53566
rect 36318 53618 36370 53630
rect 36318 53554 36370 53566
rect 36990 53618 37042 53630
rect 36990 53554 37042 53566
rect 3390 53506 3442 53518
rect 3390 53442 3442 53454
rect 5854 53506 5906 53518
rect 5854 53442 5906 53454
rect 14254 53506 14306 53518
rect 14254 53442 14306 53454
rect 16382 53506 16434 53518
rect 22094 53506 22146 53518
rect 20626 53454 20638 53506
rect 20690 53503 20702 53506
rect 20850 53503 20862 53506
rect 20690 53457 20862 53503
rect 20690 53454 20702 53457
rect 20850 53454 20862 53457
rect 20914 53454 20926 53506
rect 16382 53442 16434 53454
rect 22094 53442 22146 53454
rect 22318 53506 22370 53518
rect 22318 53442 22370 53454
rect 23438 53506 23490 53518
rect 23438 53442 23490 53454
rect 27022 53506 27074 53518
rect 27022 53442 27074 53454
rect 37326 53506 37378 53518
rect 37326 53442 37378 53454
rect 38222 53506 38274 53518
rect 38222 53442 38274 53454
rect 1344 53338 38640 53372
rect 1344 53286 19838 53338
rect 19890 53286 19942 53338
rect 19994 53286 20046 53338
rect 20098 53286 38640 53338
rect 1344 53252 38640 53286
rect 5406 53170 5458 53182
rect 7310 53170 7362 53182
rect 6290 53118 6302 53170
rect 6354 53118 6366 53170
rect 5406 53106 5458 53118
rect 7310 53106 7362 53118
rect 8654 53170 8706 53182
rect 8654 53106 8706 53118
rect 11454 53170 11506 53182
rect 16270 53170 16322 53182
rect 34974 53170 35026 53182
rect 12338 53118 12350 53170
rect 12402 53118 12414 53170
rect 18834 53118 18846 53170
rect 18898 53118 18910 53170
rect 22418 53118 22430 53170
rect 22482 53118 22494 53170
rect 33058 53118 33070 53170
rect 33122 53118 33134 53170
rect 11454 53106 11506 53118
rect 16270 53106 16322 53118
rect 34974 53106 35026 53118
rect 8206 53058 8258 53070
rect 16606 53058 16658 53070
rect 2482 53006 2494 53058
rect 2546 53006 2558 53058
rect 15138 53006 15150 53058
rect 15202 53006 15214 53058
rect 8206 52994 8258 53006
rect 16606 52994 16658 53006
rect 17502 53058 17554 53070
rect 17502 52994 17554 53006
rect 18510 53058 18562 53070
rect 18510 52994 18562 53006
rect 19406 53058 19458 53070
rect 31166 53058 31218 53070
rect 21522 53006 21534 53058
rect 21586 53006 21598 53058
rect 22082 53006 22094 53058
rect 22146 53006 22158 53058
rect 22642 53006 22654 53058
rect 22706 53006 22718 53058
rect 27346 53006 27358 53058
rect 27410 53006 27422 53058
rect 37426 53006 37438 53058
rect 37490 53006 37502 53058
rect 19406 52994 19458 53006
rect 31166 52994 31218 53006
rect 5182 52946 5234 52958
rect 6638 52946 6690 52958
rect 1810 52894 1822 52946
rect 1874 52894 1886 52946
rect 4946 52894 4958 52946
rect 5010 52894 5022 52946
rect 5618 52894 5630 52946
rect 5682 52894 5694 52946
rect 5182 52882 5234 52894
rect 6638 52882 6690 52894
rect 7982 52946 8034 52958
rect 7982 52882 8034 52894
rect 12014 52946 12066 52958
rect 19182 52946 19234 52958
rect 15810 52894 15822 52946
rect 15874 52894 15886 52946
rect 12014 52882 12066 52894
rect 19182 52882 19234 52894
rect 20078 52946 20130 52958
rect 21982 52946 22034 52958
rect 30830 52946 30882 52958
rect 20626 52894 20638 52946
rect 20690 52894 20702 52946
rect 21298 52894 21310 52946
rect 21362 52894 21374 52946
rect 28018 52894 28030 52946
rect 28082 52894 28094 52946
rect 20078 52882 20130 52894
rect 21982 52882 22034 52894
rect 30830 52882 30882 52894
rect 32286 52946 32338 52958
rect 38210 52894 38222 52946
rect 38274 52894 38286 52946
rect 32286 52882 32338 52894
rect 5294 52834 5346 52846
rect 4610 52782 4622 52834
rect 4674 52782 4686 52834
rect 5294 52770 5346 52782
rect 6862 52834 6914 52846
rect 6862 52770 6914 52782
rect 11790 52834 11842 52846
rect 23438 52834 23490 52846
rect 13010 52782 13022 52834
rect 13074 52782 13086 52834
rect 11790 52770 11842 52782
rect 23438 52770 23490 52782
rect 23886 52834 23938 52846
rect 28590 52834 28642 52846
rect 25218 52782 25230 52834
rect 25282 52782 25294 52834
rect 23886 52770 23938 52782
rect 28590 52770 28642 52782
rect 33630 52834 33682 52846
rect 33630 52770 33682 52782
rect 34078 52834 34130 52846
rect 35298 52782 35310 52834
rect 35362 52782 35374 52834
rect 34078 52770 34130 52782
rect 7646 52722 7698 52734
rect 7646 52658 7698 52670
rect 17390 52722 17442 52734
rect 17390 52658 17442 52670
rect 17726 52722 17778 52734
rect 33406 52722 33458 52734
rect 20402 52670 20414 52722
rect 20466 52670 20478 52722
rect 17726 52658 17778 52670
rect 33406 52658 33458 52670
rect 1344 52554 38640 52588
rect 1344 52502 4478 52554
rect 4530 52502 4582 52554
rect 4634 52502 4686 52554
rect 4738 52502 35198 52554
rect 35250 52502 35302 52554
rect 35354 52502 35406 52554
rect 35458 52502 38640 52554
rect 1344 52468 38640 52502
rect 35870 52386 35922 52398
rect 36978 52334 36990 52386
rect 37042 52334 37054 52386
rect 35870 52322 35922 52334
rect 12910 52274 12962 52286
rect 4834 52222 4846 52274
rect 4898 52222 4910 52274
rect 12910 52210 12962 52222
rect 14702 52274 14754 52286
rect 14702 52210 14754 52222
rect 16830 52274 16882 52286
rect 16830 52210 16882 52222
rect 17278 52274 17330 52286
rect 33854 52274 33906 52286
rect 19282 52222 19294 52274
rect 19346 52222 19358 52274
rect 22082 52222 22094 52274
rect 22146 52222 22158 52274
rect 24210 52222 24222 52274
rect 24274 52222 24286 52274
rect 31266 52222 31278 52274
rect 31330 52222 31342 52274
rect 33394 52222 33406 52274
rect 33458 52222 33470 52274
rect 17278 52210 17330 52222
rect 33854 52210 33906 52222
rect 6078 52162 6130 52174
rect 17726 52162 17778 52174
rect 20078 52162 20130 52174
rect 2034 52110 2046 52162
rect 2098 52110 2110 52162
rect 15586 52110 15598 52162
rect 15650 52110 15662 52162
rect 16258 52110 16270 52162
rect 16322 52110 16334 52162
rect 18386 52110 18398 52162
rect 18450 52110 18462 52162
rect 6078 52098 6130 52110
rect 17726 52098 17778 52110
rect 20078 52098 20130 52110
rect 20190 52162 20242 52174
rect 20190 52098 20242 52110
rect 20862 52162 20914 52174
rect 24670 52162 24722 52174
rect 21298 52110 21310 52162
rect 21362 52110 21374 52162
rect 20862 52098 20914 52110
rect 24670 52098 24722 52110
rect 25118 52162 25170 52174
rect 25118 52098 25170 52110
rect 29374 52162 29426 52174
rect 29374 52098 29426 52110
rect 29710 52162 29762 52174
rect 35310 52162 35362 52174
rect 30482 52110 30494 52162
rect 30546 52110 30558 52162
rect 29710 52098 29762 52110
rect 35310 52098 35362 52110
rect 35534 52162 35586 52174
rect 35534 52098 35586 52110
rect 36318 52162 36370 52174
rect 36318 52098 36370 52110
rect 37326 52162 37378 52174
rect 37326 52098 37378 52110
rect 37550 52162 37602 52174
rect 37550 52098 37602 52110
rect 38222 52162 38274 52174
rect 38222 52098 38274 52110
rect 16046 52050 16098 52062
rect 20302 52050 20354 52062
rect 2706 51998 2718 52050
rect 2770 51998 2782 52050
rect 18050 51998 18062 52050
rect 18114 51998 18126 52050
rect 16046 51986 16098 51998
rect 20302 51986 20354 51998
rect 20526 52050 20578 52062
rect 20526 51986 20578 51998
rect 14590 51938 14642 51950
rect 14590 51874 14642 51886
rect 15374 51938 15426 51950
rect 15374 51874 15426 51886
rect 15822 51938 15874 51950
rect 15822 51874 15874 51886
rect 15934 51938 15986 51950
rect 15934 51874 15986 51886
rect 29486 51938 29538 51950
rect 29486 51874 29538 51886
rect 30046 51938 30098 51950
rect 30046 51874 30098 51886
rect 1344 51770 38640 51804
rect 1344 51718 19838 51770
rect 19890 51718 19942 51770
rect 19994 51718 20046 51770
rect 20098 51718 38640 51770
rect 1344 51684 38640 51718
rect 3838 51602 3890 51614
rect 3838 51538 3890 51550
rect 5070 51602 5122 51614
rect 5070 51538 5122 51550
rect 16830 51602 16882 51614
rect 16830 51538 16882 51550
rect 17838 51602 17890 51614
rect 25342 51602 25394 51614
rect 24546 51550 24558 51602
rect 24610 51550 24622 51602
rect 17838 51538 17890 51550
rect 25342 51538 25394 51550
rect 25790 51602 25842 51614
rect 31166 51602 31218 51614
rect 30706 51550 30718 51602
rect 30770 51550 30782 51602
rect 25790 51538 25842 51550
rect 31166 51538 31218 51550
rect 36654 51602 36706 51614
rect 36654 51538 36706 51550
rect 3166 51490 3218 51502
rect 3166 51426 3218 51438
rect 3502 51490 3554 51502
rect 3502 51426 3554 51438
rect 18062 51490 18114 51502
rect 18062 51426 18114 51438
rect 19294 51490 19346 51502
rect 19294 51426 19346 51438
rect 21534 51490 21586 51502
rect 21534 51426 21586 51438
rect 23550 51490 23602 51502
rect 23550 51426 23602 51438
rect 4174 51378 4226 51390
rect 4174 51314 4226 51326
rect 16382 51378 16434 51390
rect 20638 51378 20690 51390
rect 22990 51378 23042 51390
rect 19170 51326 19182 51378
rect 19234 51326 19246 51378
rect 19954 51326 19966 51378
rect 20018 51326 20030 51378
rect 20402 51326 20414 51378
rect 20466 51326 20478 51378
rect 20850 51326 20862 51378
rect 20914 51326 20926 51378
rect 16382 51314 16434 51326
rect 20638 51314 20690 51326
rect 22990 51314 23042 51326
rect 30382 51378 30434 51390
rect 30382 51314 30434 51326
rect 10782 51266 10834 51278
rect 10782 51202 10834 51214
rect 15934 51266 15986 51278
rect 15934 51202 15986 51214
rect 30158 51266 30210 51278
rect 30158 51202 30210 51214
rect 18286 51154 18338 51166
rect 18610 51102 18622 51154
rect 18674 51102 18686 51154
rect 18286 51090 18338 51102
rect 1344 50986 38640 51020
rect 1344 50934 4478 50986
rect 4530 50934 4582 50986
rect 4634 50934 4686 50986
rect 4738 50934 35198 50986
rect 35250 50934 35302 50986
rect 35354 50934 35406 50986
rect 35458 50934 38640 50986
rect 1344 50900 38640 50934
rect 6302 50818 6354 50830
rect 6302 50754 6354 50766
rect 6638 50818 6690 50830
rect 6638 50754 6690 50766
rect 7310 50706 7362 50718
rect 11342 50706 11394 50718
rect 9426 50654 9438 50706
rect 9490 50654 9502 50706
rect 7310 50642 7362 50654
rect 11342 50642 11394 50654
rect 14702 50706 14754 50718
rect 14702 50642 14754 50654
rect 16606 50706 16658 50718
rect 16606 50642 16658 50654
rect 23438 50706 23490 50718
rect 27694 50706 27746 50718
rect 26786 50654 26798 50706
rect 26850 50654 26862 50706
rect 23438 50642 23490 50654
rect 27694 50642 27746 50654
rect 35198 50706 35250 50718
rect 35198 50642 35250 50654
rect 10894 50594 10946 50606
rect 9314 50542 9326 50594
rect 9378 50542 9390 50594
rect 9650 50542 9662 50594
rect 9714 50542 9726 50594
rect 10894 50530 10946 50542
rect 18622 50594 18674 50606
rect 27246 50594 27298 50606
rect 20738 50542 20750 50594
rect 20802 50542 20814 50594
rect 21746 50542 21758 50594
rect 21810 50542 21822 50594
rect 23986 50542 23998 50594
rect 24050 50542 24062 50594
rect 18622 50530 18674 50542
rect 27246 50530 27298 50542
rect 6862 50482 6914 50494
rect 15374 50482 15426 50494
rect 8866 50430 8878 50482
rect 8930 50430 8942 50482
rect 6862 50418 6914 50430
rect 15374 50418 15426 50430
rect 15598 50482 15650 50494
rect 15598 50418 15650 50430
rect 15710 50482 15762 50494
rect 15710 50418 15762 50430
rect 18062 50482 18114 50494
rect 18062 50418 18114 50430
rect 19518 50482 19570 50494
rect 21410 50430 21422 50482
rect 21474 50430 21486 50482
rect 24658 50430 24670 50482
rect 24722 50430 24734 50482
rect 19518 50418 19570 50430
rect 15934 50370 15986 50382
rect 34862 50370 34914 50382
rect 10098 50318 10110 50370
rect 10162 50318 10174 50370
rect 10546 50318 10558 50370
rect 10610 50318 10622 50370
rect 17042 50318 17054 50370
rect 17106 50318 17118 50370
rect 22418 50318 22430 50370
rect 22482 50318 22494 50370
rect 15934 50306 15986 50318
rect 34862 50306 34914 50318
rect 1344 50202 38640 50236
rect 1344 50150 19838 50202
rect 19890 50150 19942 50202
rect 19994 50150 20046 50202
rect 20098 50150 38640 50202
rect 1344 50116 38640 50150
rect 5070 50034 5122 50046
rect 5070 49970 5122 49982
rect 11118 50034 11170 50046
rect 19406 50034 19458 50046
rect 18050 49982 18062 50034
rect 18114 49982 18126 50034
rect 11118 49970 11170 49982
rect 19406 49970 19458 49982
rect 20526 50034 20578 50046
rect 20526 49970 20578 49982
rect 35646 50034 35698 50046
rect 35646 49970 35698 49982
rect 10222 49922 10274 49934
rect 20302 49922 20354 49934
rect 23326 49922 23378 49934
rect 2482 49870 2494 49922
rect 2546 49870 2558 49922
rect 16258 49870 16270 49922
rect 16322 49870 16334 49922
rect 18610 49870 18622 49922
rect 18674 49870 18686 49922
rect 20738 49870 20750 49922
rect 20802 49870 20814 49922
rect 10222 49858 10274 49870
rect 20302 49858 20354 49870
rect 23326 49858 23378 49870
rect 25566 49922 25618 49934
rect 25566 49858 25618 49870
rect 33630 49922 33682 49934
rect 33630 49858 33682 49870
rect 14814 49810 14866 49822
rect 16494 49810 16546 49822
rect 20190 49810 20242 49822
rect 25230 49810 25282 49822
rect 1810 49758 1822 49810
rect 1874 49758 1886 49810
rect 10434 49758 10446 49810
rect 10498 49758 10510 49810
rect 11666 49758 11678 49810
rect 11730 49758 11742 49810
rect 15250 49758 15262 49810
rect 15314 49758 15326 49810
rect 15922 49758 15934 49810
rect 15986 49758 15998 49810
rect 17490 49758 17502 49810
rect 17554 49758 17566 49810
rect 22306 49758 22318 49810
rect 22370 49758 22382 49810
rect 24546 49758 24558 49810
rect 24610 49758 24622 49810
rect 14814 49746 14866 49758
rect 16494 49746 16546 49758
rect 20190 49746 20242 49758
rect 25230 49746 25282 49758
rect 26126 49810 26178 49822
rect 33966 49810 34018 49822
rect 26898 49758 26910 49810
rect 26962 49758 26974 49810
rect 26126 49746 26178 49758
rect 33966 49746 34018 49758
rect 34974 49810 35026 49822
rect 34974 49746 35026 49758
rect 8206 49698 8258 49710
rect 19854 49698 19906 49710
rect 25902 49698 25954 49710
rect 30270 49698 30322 49710
rect 4610 49646 4622 49698
rect 4674 49646 4686 49698
rect 12338 49646 12350 49698
rect 12402 49646 12414 49698
rect 14466 49646 14478 49698
rect 14530 49646 14542 49698
rect 19170 49646 19182 49698
rect 19234 49646 19246 49698
rect 22978 49646 22990 49698
rect 23042 49646 23054 49698
rect 27682 49646 27694 49698
rect 27746 49646 27758 49698
rect 29810 49646 29822 49698
rect 29874 49646 29886 49698
rect 8206 49634 8258 49646
rect 7970 49534 7982 49586
rect 8034 49583 8046 49586
rect 8194 49583 8206 49586
rect 8034 49537 8206 49583
rect 8034 49534 8046 49537
rect 8194 49534 8206 49537
rect 8258 49534 8270 49586
rect 19185 49583 19231 49646
rect 19854 49634 19906 49646
rect 25902 49634 25954 49646
rect 30270 49634 30322 49646
rect 30718 49698 30770 49710
rect 30718 49634 30770 49646
rect 34638 49698 34690 49710
rect 34638 49634 34690 49646
rect 35198 49698 35250 49710
rect 35198 49634 35250 49646
rect 26462 49586 26514 49598
rect 19842 49583 19854 49586
rect 19185 49537 19854 49583
rect 19842 49534 19854 49537
rect 19906 49534 19918 49586
rect 26462 49522 26514 49534
rect 1344 49418 38640 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 38640 49418
rect 1344 49332 38640 49366
rect 13470 49250 13522 49262
rect 13470 49186 13522 49198
rect 21422 49250 21474 49262
rect 21422 49186 21474 49198
rect 7982 49138 8034 49150
rect 11678 49138 11730 49150
rect 8306 49086 8318 49138
rect 8370 49086 8382 49138
rect 10434 49086 10446 49138
rect 10498 49086 10510 49138
rect 7982 49074 8034 49086
rect 11678 49074 11730 49086
rect 12462 49138 12514 49150
rect 12462 49074 12514 49086
rect 13582 49138 13634 49150
rect 13582 49074 13634 49086
rect 15262 49138 15314 49150
rect 29710 49138 29762 49150
rect 31166 49138 31218 49150
rect 16146 49086 16158 49138
rect 16210 49086 16222 49138
rect 24882 49086 24894 49138
rect 24946 49086 24958 49138
rect 27010 49086 27022 49138
rect 27074 49086 27086 49138
rect 30482 49086 30494 49138
rect 30546 49086 30558 49138
rect 31714 49086 31726 49138
rect 31778 49086 31790 49138
rect 33842 49086 33854 49138
rect 33906 49086 33918 49138
rect 15262 49074 15314 49086
rect 29710 49074 29762 49086
rect 31166 49074 31218 49086
rect 7758 49026 7810 49038
rect 14478 49026 14530 49038
rect 11218 48974 11230 49026
rect 11282 48974 11294 49026
rect 13794 48974 13806 49026
rect 13858 48974 13870 49026
rect 7758 48962 7810 48974
rect 14478 48962 14530 48974
rect 16046 49026 16098 49038
rect 16046 48962 16098 48974
rect 18622 49026 18674 49038
rect 30270 49026 30322 49038
rect 35310 49026 35362 49038
rect 20738 48974 20750 49026
rect 20802 48974 20814 49026
rect 22642 48974 22654 49026
rect 22706 48974 22718 49026
rect 22866 48974 22878 49026
rect 22930 48974 22942 49026
rect 27682 48974 27694 49026
rect 27746 48974 27758 49026
rect 30034 48974 30046 49026
rect 30098 48974 30110 49026
rect 34626 48974 34638 49026
rect 34690 48974 34702 49026
rect 35746 48974 35758 49026
rect 35810 48974 35822 49026
rect 37090 48974 37102 49026
rect 37154 48974 37166 49026
rect 18622 48962 18674 48974
rect 30270 48962 30322 48974
rect 35310 48962 35362 48974
rect 7086 48914 7138 48926
rect 14142 48914 14194 48926
rect 7410 48862 7422 48914
rect 7474 48862 7486 48914
rect 7086 48850 7138 48862
rect 14142 48850 14194 48862
rect 15598 48914 15650 48926
rect 15598 48850 15650 48862
rect 17614 48914 17666 48926
rect 17614 48850 17666 48862
rect 20190 48914 20242 48926
rect 30606 48914 30658 48926
rect 22082 48862 22094 48914
rect 22146 48862 22158 48914
rect 23090 48862 23102 48914
rect 23154 48862 23166 48914
rect 20190 48850 20242 48862
rect 30606 48850 30658 48862
rect 6750 48802 6802 48814
rect 6750 48738 6802 48750
rect 13022 48802 13074 48814
rect 13022 48738 13074 48750
rect 14254 48802 14306 48814
rect 14254 48738 14306 48750
rect 14926 48802 14978 48814
rect 14926 48738 14978 48750
rect 15822 48802 15874 48814
rect 15822 48738 15874 48750
rect 16158 48802 16210 48814
rect 28254 48802 28306 48814
rect 17042 48750 17054 48802
rect 17106 48750 17118 48802
rect 16158 48738 16210 48750
rect 28254 48738 28306 48750
rect 29262 48802 29314 48814
rect 29262 48738 29314 48750
rect 30494 48802 30546 48814
rect 30494 48738 30546 48750
rect 35198 48802 35250 48814
rect 35198 48738 35250 48750
rect 35422 48802 35474 48814
rect 35422 48738 35474 48750
rect 35534 48802 35586 48814
rect 35534 48738 35586 48750
rect 36206 48802 36258 48814
rect 36206 48738 36258 48750
rect 37326 48802 37378 48814
rect 37326 48738 37378 48750
rect 38222 48802 38274 48814
rect 38222 48738 38274 48750
rect 1344 48634 38640 48668
rect 1344 48582 19838 48634
rect 19890 48582 19942 48634
rect 19994 48582 20046 48634
rect 20098 48582 38640 48634
rect 1344 48548 38640 48582
rect 9662 48466 9714 48478
rect 9662 48402 9714 48414
rect 10222 48466 10274 48478
rect 10222 48402 10274 48414
rect 10334 48466 10386 48478
rect 10334 48402 10386 48414
rect 10446 48466 10498 48478
rect 13918 48466 13970 48478
rect 24670 48466 24722 48478
rect 11330 48414 11342 48466
rect 11394 48414 11406 48466
rect 19394 48414 19406 48466
rect 19458 48414 19470 48466
rect 24210 48414 24222 48466
rect 24274 48414 24286 48466
rect 10446 48402 10498 48414
rect 13918 48402 13970 48414
rect 24670 48402 24722 48414
rect 25342 48466 25394 48478
rect 25342 48402 25394 48414
rect 27134 48466 27186 48478
rect 27134 48402 27186 48414
rect 28030 48466 28082 48478
rect 28030 48402 28082 48414
rect 33854 48466 33906 48478
rect 33854 48402 33906 48414
rect 34190 48466 34242 48478
rect 34190 48402 34242 48414
rect 34750 48466 34802 48478
rect 34750 48402 34802 48414
rect 3726 48354 3778 48366
rect 11902 48354 11954 48366
rect 6738 48302 6750 48354
rect 6802 48302 6814 48354
rect 3726 48290 3778 48302
rect 11902 48290 11954 48302
rect 14590 48354 14642 48366
rect 14590 48290 14642 48302
rect 17950 48354 18002 48366
rect 26798 48354 26850 48366
rect 21074 48302 21086 48354
rect 21138 48302 21150 48354
rect 22978 48302 22990 48354
rect 23042 48302 23054 48354
rect 17950 48290 18002 48302
rect 26798 48290 26850 48302
rect 33630 48354 33682 48366
rect 37426 48302 37438 48354
rect 37490 48302 37502 48354
rect 33630 48290 33682 48302
rect 4062 48242 4114 48254
rect 16158 48242 16210 48254
rect 21870 48242 21922 48254
rect 23886 48242 23938 48254
rect 4722 48190 4734 48242
rect 4786 48190 4798 48242
rect 5954 48190 5966 48242
rect 6018 48190 6030 48242
rect 9986 48190 9998 48242
rect 10050 48190 10062 48242
rect 10658 48190 10670 48242
rect 10722 48190 10734 48242
rect 15362 48190 15374 48242
rect 15426 48190 15438 48242
rect 16370 48190 16382 48242
rect 16434 48190 16446 48242
rect 17378 48190 17390 48242
rect 17442 48190 17454 48242
rect 21186 48190 21198 48242
rect 21250 48190 21262 48242
rect 22642 48190 22654 48242
rect 22706 48190 22718 48242
rect 4062 48178 4114 48190
rect 16158 48178 16210 48190
rect 21870 48178 21922 48190
rect 23886 48178 23938 48190
rect 25678 48242 25730 48254
rect 34078 48242 34130 48254
rect 28466 48190 28478 48242
rect 28530 48190 28542 48242
rect 38098 48190 38110 48242
rect 38162 48190 38174 48242
rect 25678 48178 25730 48190
rect 34078 48178 34130 48190
rect 5294 48130 5346 48142
rect 12350 48130 12402 48142
rect 8866 48078 8878 48130
rect 8930 48078 8942 48130
rect 5294 48066 5346 48078
rect 12350 48066 12402 48078
rect 12798 48130 12850 48142
rect 12798 48066 12850 48078
rect 14366 48130 14418 48142
rect 23662 48130 23714 48142
rect 15810 48078 15822 48130
rect 15874 48078 15886 48130
rect 16482 48078 16494 48130
rect 16546 48078 16558 48130
rect 22194 48078 22206 48130
rect 22258 48078 22270 48130
rect 23090 48078 23102 48130
rect 23154 48078 23166 48130
rect 14366 48066 14418 48078
rect 23662 48066 23714 48078
rect 26126 48130 26178 48142
rect 26126 48066 26178 48078
rect 27582 48130 27634 48142
rect 32286 48130 32338 48142
rect 29250 48078 29262 48130
rect 29314 48078 29326 48130
rect 31378 48078 31390 48130
rect 31442 48078 31454 48130
rect 27582 48066 27634 48078
rect 32286 48066 32338 48078
rect 33182 48130 33234 48142
rect 33182 48066 33234 48078
rect 33966 48130 34018 48142
rect 35298 48078 35310 48130
rect 35362 48078 35374 48130
rect 33966 48066 34018 48078
rect 5070 48018 5122 48030
rect 5070 47954 5122 47966
rect 11678 48018 11730 48030
rect 11678 47954 11730 47966
rect 14702 48018 14754 48030
rect 32062 48018 32114 48030
rect 21634 47966 21646 48018
rect 21698 47966 21710 48018
rect 31714 47966 31726 48018
rect 31778 47966 31790 48018
rect 14702 47954 14754 47966
rect 32062 47954 32114 47966
rect 1344 47850 38640 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 38640 47850
rect 1344 47764 38640 47798
rect 14242 47630 14254 47682
rect 14306 47679 14318 47682
rect 14690 47679 14702 47682
rect 14306 47633 14702 47679
rect 14306 47630 14318 47633
rect 14690 47630 14702 47633
rect 14754 47630 14766 47682
rect 14366 47570 14418 47582
rect 2930 47518 2942 47570
rect 2994 47518 3006 47570
rect 5058 47518 5070 47570
rect 5122 47518 5134 47570
rect 8978 47518 8990 47570
rect 9042 47518 9054 47570
rect 12898 47518 12910 47570
rect 12962 47518 12974 47570
rect 14366 47506 14418 47518
rect 14814 47570 14866 47582
rect 27470 47570 27522 47582
rect 37550 47570 37602 47582
rect 15474 47518 15486 47570
rect 15538 47518 15550 47570
rect 24770 47518 24782 47570
rect 24834 47518 24846 47570
rect 34738 47518 34750 47570
rect 34802 47518 34814 47570
rect 14814 47506 14866 47518
rect 27470 47506 27522 47518
rect 37550 47506 37602 47518
rect 9438 47458 9490 47470
rect 30830 47458 30882 47470
rect 35534 47458 35586 47470
rect 37326 47458 37378 47470
rect 2258 47406 2270 47458
rect 2322 47406 2334 47458
rect 6066 47406 6078 47458
rect 6130 47406 6142 47458
rect 10098 47406 10110 47458
rect 10162 47406 10174 47458
rect 15698 47406 15710 47458
rect 15762 47406 15774 47458
rect 16482 47406 16494 47458
rect 16546 47406 16558 47458
rect 18498 47406 18510 47458
rect 18562 47406 18574 47458
rect 21858 47406 21870 47458
rect 21922 47406 21934 47458
rect 29698 47406 29710 47458
rect 29762 47406 29774 47458
rect 31266 47406 31278 47458
rect 31330 47406 31342 47458
rect 31826 47406 31838 47458
rect 31890 47406 31902 47458
rect 35074 47406 35086 47458
rect 35138 47406 35150 47458
rect 35746 47406 35758 47458
rect 35810 47406 35822 47458
rect 36194 47406 36206 47458
rect 36258 47406 36270 47458
rect 9438 47394 9490 47406
rect 30830 47394 30882 47406
rect 35534 47394 35586 47406
rect 37326 47394 37378 47406
rect 15038 47346 15090 47358
rect 6850 47294 6862 47346
rect 6914 47294 6926 47346
rect 10770 47294 10782 47346
rect 10834 47294 10846 47346
rect 15038 47282 15090 47294
rect 15486 47346 15538 47358
rect 15486 47282 15538 47294
rect 17054 47346 17106 47358
rect 17054 47282 17106 47294
rect 19070 47346 19122 47358
rect 19070 47282 19122 47294
rect 29486 47346 29538 47358
rect 29486 47282 29538 47294
rect 31502 47346 31554 47358
rect 32610 47294 32622 47346
rect 32674 47294 32686 47346
rect 36978 47294 36990 47346
rect 37042 47294 37054 47346
rect 31502 47282 31554 47294
rect 5742 47234 5794 47246
rect 5742 47170 5794 47182
rect 13582 47234 13634 47246
rect 13582 47170 13634 47182
rect 15262 47234 15314 47246
rect 15262 47170 15314 47182
rect 16270 47234 16322 47246
rect 20750 47234 20802 47246
rect 20066 47182 20078 47234
rect 20130 47182 20142 47234
rect 16270 47170 16322 47182
rect 20750 47170 20802 47182
rect 27022 47234 27074 47246
rect 27022 47170 27074 47182
rect 27918 47234 27970 47246
rect 27918 47170 27970 47182
rect 28366 47234 28418 47246
rect 28366 47170 28418 47182
rect 35310 47234 35362 47246
rect 35310 47170 35362 47182
rect 35422 47234 35474 47246
rect 35422 47170 35474 47182
rect 36430 47234 36482 47246
rect 36430 47170 36482 47182
rect 37998 47234 38050 47246
rect 37998 47170 38050 47182
rect 1344 47066 38640 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 38640 47066
rect 1344 46980 38640 47014
rect 7422 46898 7474 46910
rect 11230 46898 11282 46910
rect 10770 46846 10782 46898
rect 10834 46895 10846 46898
rect 10994 46895 11006 46898
rect 10834 46849 11006 46895
rect 10834 46846 10846 46849
rect 10994 46846 11006 46849
rect 11058 46846 11070 46898
rect 7422 46834 7474 46846
rect 11230 46834 11282 46846
rect 13806 46898 13858 46910
rect 13806 46834 13858 46846
rect 14254 46898 14306 46910
rect 14254 46834 14306 46846
rect 17838 46898 17890 46910
rect 17838 46834 17890 46846
rect 24222 46898 24274 46910
rect 27246 46898 27298 46910
rect 33406 46898 33458 46910
rect 26226 46846 26238 46898
rect 26290 46846 26302 46898
rect 29586 46846 29598 46898
rect 29650 46846 29662 46898
rect 24222 46834 24274 46846
rect 27246 46834 27298 46846
rect 33406 46834 33458 46846
rect 34638 46898 34690 46910
rect 34638 46834 34690 46846
rect 35086 46898 35138 46910
rect 35086 46834 35138 46846
rect 14142 46786 14194 46798
rect 25230 46786 25282 46798
rect 19394 46734 19406 46786
rect 19458 46734 19470 46786
rect 19954 46734 19966 46786
rect 20018 46734 20030 46786
rect 23650 46734 23662 46786
rect 23714 46734 23726 46786
rect 37426 46734 37438 46786
rect 37490 46734 37502 46786
rect 14142 46722 14194 46734
rect 25230 46722 25282 46734
rect 7758 46674 7810 46686
rect 24670 46674 24722 46686
rect 11442 46622 11454 46674
rect 11506 46622 11518 46674
rect 19506 46622 19518 46674
rect 19570 46622 19582 46674
rect 21522 46622 21534 46674
rect 21586 46622 21598 46674
rect 21970 46622 21982 46674
rect 22034 46622 22046 46674
rect 7758 46610 7810 46622
rect 24670 46610 24722 46622
rect 25454 46674 25506 46686
rect 25454 46610 25506 46622
rect 25678 46674 25730 46686
rect 25678 46610 25730 46622
rect 25790 46674 25842 46686
rect 25790 46610 25842 46622
rect 27694 46674 27746 46686
rect 27694 46610 27746 46622
rect 28590 46674 28642 46686
rect 38098 46622 38110 46674
rect 38162 46622 38174 46674
rect 28590 46610 28642 46622
rect 5294 46562 5346 46574
rect 5294 46498 5346 46510
rect 9662 46562 9714 46574
rect 9662 46498 9714 46510
rect 15038 46562 15090 46574
rect 15038 46498 15090 46510
rect 15598 46562 15650 46574
rect 15598 46498 15650 46510
rect 15934 46562 15986 46574
rect 15934 46498 15986 46510
rect 16494 46562 16546 46574
rect 16494 46498 16546 46510
rect 16830 46562 16882 46574
rect 25566 46562 25618 46574
rect 22306 46510 22318 46562
rect 22370 46510 22382 46562
rect 16830 46498 16882 46510
rect 25566 46498 25618 46510
rect 26798 46562 26850 46574
rect 26798 46498 26850 46510
rect 28142 46562 28194 46574
rect 28142 46498 28194 46510
rect 29038 46562 29090 46574
rect 29038 46498 29090 46510
rect 30158 46562 30210 46574
rect 30158 46498 30210 46510
rect 30606 46562 30658 46574
rect 35298 46510 35310 46562
rect 35362 46510 35374 46562
rect 30606 46498 30658 46510
rect 14254 46450 14306 46462
rect 26574 46450 26626 46462
rect 16034 46398 16046 46450
rect 16098 46447 16110 46450
rect 16706 46447 16718 46450
rect 16098 46401 16718 46447
rect 16098 46398 16110 46401
rect 16706 46398 16718 46401
rect 16770 46398 16782 46450
rect 18274 46398 18286 46450
rect 18338 46398 18350 46450
rect 14254 46386 14306 46398
rect 26574 46386 26626 46398
rect 29934 46450 29986 46462
rect 29934 46386 29986 46398
rect 1344 46282 38640 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 38640 46282
rect 1344 46196 38640 46230
rect 13470 46114 13522 46126
rect 37538 46062 37550 46114
rect 37602 46062 37614 46114
rect 13470 46050 13522 46062
rect 4622 46002 4674 46014
rect 4622 45938 4674 45950
rect 14030 46002 14082 46014
rect 30606 46002 30658 46014
rect 21746 45950 21758 46002
rect 21810 45950 21822 46002
rect 14030 45938 14082 45950
rect 30606 45938 30658 45950
rect 31054 46002 31106 46014
rect 31054 45938 31106 45950
rect 36990 46002 37042 46014
rect 36990 45938 37042 45950
rect 3950 45890 4002 45902
rect 3950 45826 4002 45838
rect 4174 45890 4226 45902
rect 4174 45826 4226 45838
rect 12910 45890 12962 45902
rect 12910 45826 12962 45838
rect 13806 45890 13858 45902
rect 13806 45826 13858 45838
rect 15934 45890 15986 45902
rect 15934 45826 15986 45838
rect 16382 45890 16434 45902
rect 16382 45826 16434 45838
rect 18398 45890 18450 45902
rect 26238 45890 26290 45902
rect 20514 45838 20526 45890
rect 20578 45838 20590 45890
rect 21522 45838 21534 45890
rect 21586 45838 21598 45890
rect 24098 45838 24110 45890
rect 24162 45838 24174 45890
rect 18398 45826 18450 45838
rect 26238 45826 26290 45838
rect 28478 45890 28530 45902
rect 28478 45826 28530 45838
rect 37214 45890 37266 45902
rect 37214 45826 37266 45838
rect 16158 45778 16210 45790
rect 19854 45778 19906 45790
rect 23550 45778 23602 45790
rect 16818 45726 16830 45778
rect 16882 45726 16894 45778
rect 22754 45726 22766 45778
rect 22818 45726 22830 45778
rect 16158 45714 16210 45726
rect 19854 45714 19906 45726
rect 23550 45714 23602 45726
rect 23662 45778 23714 45790
rect 23662 45714 23714 45726
rect 23886 45778 23938 45790
rect 26798 45778 26850 45790
rect 24210 45726 24222 45778
rect 24274 45726 24286 45778
rect 23886 45714 23938 45726
rect 26798 45714 26850 45726
rect 28366 45778 28418 45790
rect 28366 45714 28418 45726
rect 14814 45666 14866 45678
rect 3602 45614 3614 45666
rect 3666 45614 3678 45666
rect 14814 45602 14866 45614
rect 15150 45666 15202 45678
rect 28142 45666 28194 45678
rect 15586 45614 15598 45666
rect 15650 45614 15662 45666
rect 16930 45614 16942 45666
rect 16994 45614 17006 45666
rect 27794 45614 27806 45666
rect 27858 45614 27870 45666
rect 15150 45602 15202 45614
rect 28142 45602 28194 45614
rect 29262 45666 29314 45678
rect 29262 45602 29314 45614
rect 29710 45666 29762 45678
rect 29710 45602 29762 45614
rect 30158 45666 30210 45678
rect 30158 45602 30210 45614
rect 34974 45666 35026 45678
rect 34974 45602 35026 45614
rect 36430 45666 36482 45678
rect 36430 45602 36482 45614
rect 38222 45666 38274 45678
rect 38222 45602 38274 45614
rect 1344 45498 38640 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 38640 45498
rect 1344 45412 38640 45446
rect 14366 45330 14418 45342
rect 7970 45278 7982 45330
rect 8034 45278 8046 45330
rect 11330 45278 11342 45330
rect 11394 45278 11406 45330
rect 14366 45266 14418 45278
rect 17502 45330 17554 45342
rect 25330 45278 25342 45330
rect 25394 45278 25406 45330
rect 17502 45266 17554 45278
rect 17950 45218 18002 45230
rect 17950 45154 18002 45166
rect 23214 45218 23266 45230
rect 25554 45166 25566 45218
rect 25618 45166 25630 45218
rect 26002 45166 26014 45218
rect 26066 45166 26078 45218
rect 23214 45154 23266 45166
rect 27134 45162 27186 45174
rect 28242 45166 28254 45218
rect 28306 45166 28318 45218
rect 14030 45106 14082 45118
rect 17502 45106 17554 45118
rect 1810 45054 1822 45106
rect 1874 45054 1886 45106
rect 15362 45054 15374 45106
rect 15426 45054 15438 45106
rect 14030 45042 14082 45054
rect 17502 45042 17554 45054
rect 19182 45106 19234 45118
rect 23438 45106 23490 45118
rect 20514 45054 20526 45106
rect 20578 45054 20590 45106
rect 19182 45042 19234 45054
rect 23438 45042 23490 45054
rect 23662 45106 23714 45118
rect 23662 45042 23714 45054
rect 23774 45106 23826 45118
rect 26574 45106 26626 45118
rect 26338 45054 26350 45106
rect 26402 45054 26414 45106
rect 26898 45054 26910 45106
rect 26962 45054 26974 45106
rect 27134 45098 27186 45110
rect 27570 45054 27582 45106
rect 27634 45054 27646 45106
rect 23774 45042 23826 45054
rect 26574 45042 26626 45054
rect 5070 44994 5122 45006
rect 2482 44942 2494 44994
rect 2546 44942 2558 44994
rect 4610 44942 4622 44994
rect 4674 44942 4686 44994
rect 5070 44930 5122 44942
rect 7646 44994 7698 45006
rect 7646 44930 7698 44942
rect 8542 44994 8594 45006
rect 8542 44930 8594 44942
rect 11006 44994 11058 45006
rect 11006 44930 11058 44942
rect 11678 44994 11730 45006
rect 11678 44930 11730 44942
rect 11902 44994 11954 45006
rect 11902 44930 11954 44942
rect 12462 44994 12514 45006
rect 12462 44930 12514 44942
rect 14814 44994 14866 45006
rect 30830 44994 30882 45006
rect 15250 44942 15262 44994
rect 15314 44942 15326 44994
rect 16818 44942 16830 44994
rect 16882 44942 16894 44994
rect 30370 44942 30382 44994
rect 30434 44942 30446 44994
rect 14814 44930 14866 44942
rect 30830 44930 30882 44942
rect 31278 44994 31330 45006
rect 31278 44930 31330 44942
rect 31726 44994 31778 45006
rect 31726 44930 31778 44942
rect 8318 44882 8370 44894
rect 8318 44818 8370 44830
rect 21310 44882 21362 44894
rect 27246 44882 27298 44894
rect 24210 44830 24222 44882
rect 24274 44830 24286 44882
rect 21310 44818 21362 44830
rect 27246 44818 27298 44830
rect 1344 44714 38640 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 38640 44714
rect 1344 44628 38640 44662
rect 14478 44434 14530 44446
rect 14478 44370 14530 44382
rect 20302 44434 20354 44446
rect 20302 44370 20354 44382
rect 20750 44434 20802 44446
rect 20750 44370 20802 44382
rect 22542 44434 22594 44446
rect 22542 44370 22594 44382
rect 28478 44434 28530 44446
rect 28478 44370 28530 44382
rect 29710 44434 29762 44446
rect 29710 44370 29762 44382
rect 31950 44434 32002 44446
rect 31950 44370 32002 44382
rect 2270 44322 2322 44334
rect 2270 44258 2322 44270
rect 3278 44322 3330 44334
rect 3950 44322 4002 44334
rect 3602 44270 3614 44322
rect 3666 44270 3678 44322
rect 3278 44258 3330 44270
rect 3950 44258 4002 44270
rect 4174 44322 4226 44334
rect 18062 44322 18114 44334
rect 24670 44322 24722 44334
rect 27134 44322 27186 44334
rect 15922 44270 15934 44322
rect 15986 44270 15998 44322
rect 21298 44270 21310 44322
rect 21362 44270 21374 44322
rect 26786 44270 26798 44322
rect 26850 44270 26862 44322
rect 4174 44258 4226 44270
rect 18062 44258 18114 44270
rect 24670 44258 24722 44270
rect 27134 44258 27186 44270
rect 27358 44322 27410 44334
rect 27358 44258 27410 44270
rect 27582 44322 27634 44334
rect 27582 44258 27634 44270
rect 30270 44322 30322 44334
rect 30270 44258 30322 44270
rect 30494 44322 30546 44334
rect 30494 44258 30546 44270
rect 32398 44322 32450 44334
rect 32398 44258 32450 44270
rect 2942 44210 2994 44222
rect 2942 44146 2994 44158
rect 6638 44210 6690 44222
rect 6638 44146 6690 44158
rect 17054 44210 17106 44222
rect 17054 44146 17106 44158
rect 18510 44210 18562 44222
rect 23662 44210 23714 44222
rect 21522 44158 21534 44210
rect 21586 44158 21598 44210
rect 22194 44158 22206 44210
rect 22258 44158 22270 44210
rect 18510 44146 18562 44158
rect 23662 44146 23714 44158
rect 25006 44210 25058 44222
rect 25006 44146 25058 44158
rect 25678 44210 25730 44222
rect 25678 44146 25730 44158
rect 29262 44210 29314 44222
rect 29262 44146 29314 44158
rect 30606 44210 30658 44222
rect 30606 44146 30658 44158
rect 31166 44210 31218 44222
rect 31166 44146 31218 44158
rect 2606 44098 2658 44110
rect 2606 44034 2658 44046
rect 4622 44098 4674 44110
rect 4622 44034 4674 44046
rect 6974 44098 7026 44110
rect 6974 44034 7026 44046
rect 15150 44098 15202 44110
rect 15150 44034 15202 44046
rect 15598 44098 15650 44110
rect 15598 44034 15650 44046
rect 18174 44098 18226 44110
rect 30382 44098 30434 44110
rect 27906 44046 27918 44098
rect 27970 44046 27982 44098
rect 18174 44034 18226 44046
rect 30382 44034 30434 44046
rect 30718 44098 30770 44110
rect 30718 44034 30770 44046
rect 31502 44098 31554 44110
rect 31502 44034 31554 44046
rect 32846 44098 32898 44110
rect 32846 44034 32898 44046
rect 1344 43930 38640 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 38640 43930
rect 1344 43844 38640 43878
rect 24670 43762 24722 43774
rect 19282 43710 19294 43762
rect 19346 43710 19358 43762
rect 24670 43698 24722 43710
rect 16382 43650 16434 43662
rect 2930 43598 2942 43650
rect 2994 43598 3006 43650
rect 16382 43586 16434 43598
rect 17614 43650 17666 43662
rect 20414 43650 20466 43662
rect 23662 43650 23714 43662
rect 17826 43598 17838 43650
rect 17890 43598 17902 43650
rect 23426 43598 23438 43650
rect 23490 43598 23502 43650
rect 17614 43586 17666 43598
rect 20414 43586 20466 43598
rect 23662 43586 23714 43598
rect 23774 43650 23826 43662
rect 23774 43586 23826 43598
rect 29038 43650 29090 43662
rect 31714 43598 31726 43650
rect 31778 43598 31790 43650
rect 29038 43586 29090 43598
rect 5518 43538 5570 43550
rect 16718 43538 16770 43550
rect 2146 43486 2158 43538
rect 2210 43486 2222 43538
rect 6178 43486 6190 43538
rect 6242 43486 6254 43538
rect 11442 43486 11454 43538
rect 11506 43486 11518 43538
rect 15138 43486 15150 43538
rect 15202 43486 15214 43538
rect 16146 43486 16158 43538
rect 16210 43486 16222 43538
rect 5518 43474 5570 43486
rect 16718 43474 16770 43486
rect 16942 43538 16994 43550
rect 16942 43474 16994 43486
rect 19518 43538 19570 43550
rect 21982 43538 22034 43550
rect 24334 43538 24386 43550
rect 19842 43486 19854 43538
rect 19906 43486 19918 43538
rect 22530 43486 22542 43538
rect 22594 43486 22606 43538
rect 23202 43486 23214 43538
rect 23266 43486 23278 43538
rect 23986 43486 23998 43538
rect 24050 43486 24062 43538
rect 28354 43486 28366 43538
rect 28418 43486 28430 43538
rect 32386 43486 32398 43538
rect 32450 43486 32462 43538
rect 19518 43474 19570 43486
rect 21982 43474 22034 43486
rect 24334 43474 24386 43486
rect 9662 43426 9714 43438
rect 5058 43374 5070 43426
rect 5122 43374 5134 43426
rect 6850 43374 6862 43426
rect 6914 43374 6926 43426
rect 8978 43374 8990 43426
rect 9042 43374 9054 43426
rect 9662 43362 9714 43374
rect 10110 43426 10162 43438
rect 33182 43426 33234 43438
rect 12114 43374 12126 43426
rect 12178 43374 12190 43426
rect 14242 43374 14254 43426
rect 14306 43374 14318 43426
rect 25554 43374 25566 43426
rect 25618 43374 25630 43426
rect 27682 43374 27694 43426
rect 27746 43374 27758 43426
rect 29586 43374 29598 43426
rect 29650 43374 29662 43426
rect 10110 43362 10162 43374
rect 33182 43362 33234 43374
rect 34638 43426 34690 43438
rect 34638 43362 34690 43374
rect 21870 43314 21922 43326
rect 15362 43262 15374 43314
rect 15426 43262 15438 43314
rect 15810 43262 15822 43314
rect 15874 43262 15886 43314
rect 21870 43250 21922 43262
rect 34526 43314 34578 43326
rect 34526 43250 34578 43262
rect 1344 43146 38640 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 38640 43146
rect 1344 43060 38640 43094
rect 30942 42978 30994 42990
rect 6178 42926 6190 42978
rect 6242 42926 6254 42978
rect 30034 42926 30046 42978
rect 30098 42926 30110 42978
rect 30942 42914 30994 42926
rect 5630 42866 5682 42878
rect 16270 42866 16322 42878
rect 7298 42814 7310 42866
rect 7362 42814 7374 42866
rect 9426 42814 9438 42866
rect 9490 42814 9502 42866
rect 5630 42802 5682 42814
rect 16270 42802 16322 42814
rect 20750 42866 20802 42878
rect 29486 42866 29538 42878
rect 27122 42814 27134 42866
rect 27186 42814 27198 42866
rect 27906 42814 27918 42866
rect 27970 42814 27982 42866
rect 20750 42802 20802 42814
rect 5070 42754 5122 42766
rect 5070 42690 5122 42702
rect 5854 42754 5906 42766
rect 10222 42754 10274 42766
rect 6626 42702 6638 42754
rect 6690 42702 6702 42754
rect 5854 42690 5906 42702
rect 10222 42690 10274 42702
rect 10334 42754 10386 42766
rect 21310 42754 21362 42766
rect 21522 42758 21534 42810
rect 21586 42758 21598 42810
rect 29486 42802 29538 42814
rect 31390 42866 31442 42878
rect 31390 42802 31442 42814
rect 32286 42866 32338 42878
rect 36430 42866 36482 42878
rect 33058 42814 33070 42866
rect 33122 42814 33134 42866
rect 32286 42802 32338 42814
rect 36430 42802 36482 42814
rect 38222 42866 38274 42878
rect 38222 42802 38274 42814
rect 12562 42702 12574 42754
rect 12626 42702 12638 42754
rect 15138 42702 15150 42754
rect 15202 42702 15214 42754
rect 18050 42702 18062 42754
rect 18114 42702 18126 42754
rect 20290 42702 20302 42754
rect 20354 42702 20366 42754
rect 10334 42690 10386 42702
rect 21310 42690 21362 42702
rect 21758 42754 21810 42766
rect 21758 42690 21810 42702
rect 24222 42754 24274 42766
rect 29710 42754 29762 42766
rect 26338 42702 26350 42754
rect 26402 42702 26414 42754
rect 27010 42702 27022 42754
rect 27074 42702 27086 42754
rect 28130 42702 28142 42754
rect 28194 42702 28206 42754
rect 24222 42690 24274 42702
rect 29710 42690 29762 42702
rect 30606 42754 30658 42766
rect 35858 42702 35870 42754
rect 35922 42702 35934 42754
rect 30606 42690 30658 42702
rect 9774 42642 9826 42654
rect 9774 42578 9826 42590
rect 9998 42642 10050 42654
rect 9998 42578 10050 42590
rect 11342 42642 11394 42654
rect 11342 42578 11394 42590
rect 12350 42642 12402 42654
rect 17614 42642 17666 42654
rect 15362 42590 15374 42642
rect 15426 42590 15438 42642
rect 15922 42590 15934 42642
rect 15986 42590 15998 42642
rect 12350 42578 12402 42590
rect 17614 42578 17666 42590
rect 19070 42642 19122 42654
rect 25790 42642 25842 42654
rect 30382 42642 30434 42654
rect 36990 42642 37042 42654
rect 22530 42590 22542 42642
rect 22594 42590 22606 42642
rect 26786 42590 26798 42642
rect 26850 42590 26862 42642
rect 35186 42590 35198 42642
rect 35250 42590 35262 42642
rect 19070 42578 19122 42590
rect 25790 42578 25842 42590
rect 30382 42578 30434 42590
rect 36990 42578 37042 42590
rect 10110 42530 10162 42542
rect 10110 42466 10162 42478
rect 11006 42530 11058 42542
rect 11006 42466 11058 42478
rect 14366 42530 14418 42542
rect 14366 42466 14418 42478
rect 14814 42530 14866 42542
rect 31838 42530 31890 42542
rect 16706 42478 16718 42530
rect 16770 42478 16782 42530
rect 22082 42478 22094 42530
rect 22146 42478 22158 42530
rect 26226 42478 26238 42530
rect 26290 42478 26302 42530
rect 14814 42466 14866 42478
rect 31838 42466 31890 42478
rect 32734 42530 32786 42542
rect 32734 42466 32786 42478
rect 37326 42530 37378 42542
rect 37326 42466 37378 42478
rect 1344 42362 38640 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 38640 42362
rect 1344 42276 38640 42310
rect 15486 42194 15538 42206
rect 12562 42142 12574 42194
rect 12626 42142 12638 42194
rect 15486 42130 15538 42142
rect 16382 42194 16434 42206
rect 16382 42130 16434 42142
rect 16830 42194 16882 42206
rect 25454 42194 25506 42206
rect 18946 42142 18958 42194
rect 19010 42142 19022 42194
rect 16830 42130 16882 42142
rect 25454 42130 25506 42142
rect 25678 42194 25730 42206
rect 25678 42130 25730 42142
rect 26462 42194 26514 42206
rect 26462 42130 26514 42142
rect 26686 42194 26738 42206
rect 26686 42130 26738 42142
rect 27358 42194 27410 42206
rect 27358 42130 27410 42142
rect 34862 42194 34914 42206
rect 34862 42130 34914 42142
rect 5630 42082 5682 42094
rect 5630 42018 5682 42030
rect 5854 42082 5906 42094
rect 5854 42018 5906 42030
rect 9550 42082 9602 42094
rect 9550 42018 9602 42030
rect 10894 42082 10946 42094
rect 10894 42018 10946 42030
rect 15934 42082 15986 42094
rect 20638 42082 20690 42094
rect 17490 42030 17502 42082
rect 17554 42030 17566 42082
rect 15934 42018 15986 42030
rect 20638 42018 20690 42030
rect 23326 42082 23378 42094
rect 31278 42082 31330 42094
rect 29474 42030 29486 42082
rect 29538 42030 29550 42082
rect 29922 42030 29934 42082
rect 29986 42030 29998 42082
rect 37426 42030 37438 42082
rect 37490 42030 37502 42082
rect 23326 42018 23378 42030
rect 31278 42018 31330 42030
rect 6078 41970 6130 41982
rect 8094 41970 8146 41982
rect 6290 41918 6302 41970
rect 6354 41918 6366 41970
rect 6078 41906 6130 41918
rect 8094 41906 8146 41918
rect 10558 41970 10610 41982
rect 10558 41906 10610 41918
rect 13134 41970 13186 41982
rect 13134 41906 13186 41918
rect 19182 41970 19234 41982
rect 21646 41970 21698 41982
rect 19506 41918 19518 41970
rect 19570 41918 19582 41970
rect 19182 41906 19234 41918
rect 21646 41906 21698 41918
rect 21870 41970 21922 41982
rect 21870 41906 21922 41918
rect 22094 41970 22146 41982
rect 22094 41906 22146 41918
rect 23550 41970 23602 41982
rect 26798 41970 26850 41982
rect 25218 41918 25230 41970
rect 25282 41918 25294 41970
rect 26226 41918 26238 41970
rect 26290 41918 26302 41970
rect 23550 41906 23602 41918
rect 26798 41906 26850 41918
rect 27022 41970 27074 41982
rect 27022 41906 27074 41918
rect 28926 41970 28978 41982
rect 28926 41906 28978 41918
rect 30494 41970 30546 41982
rect 34626 41918 34638 41970
rect 34690 41918 34702 41970
rect 38210 41918 38222 41970
rect 38274 41918 38286 41970
rect 30494 41906 30546 41918
rect 7198 41858 7250 41870
rect 6178 41806 6190 41858
rect 6242 41806 6254 41858
rect 7198 41794 7250 41806
rect 7646 41858 7698 41870
rect 7646 41794 7698 41806
rect 9774 41858 9826 41870
rect 9774 41794 9826 41806
rect 10110 41858 10162 41870
rect 10110 41794 10162 41806
rect 11342 41858 11394 41870
rect 11342 41794 11394 41806
rect 12350 41858 12402 41870
rect 12350 41794 12402 41806
rect 12910 41858 12962 41870
rect 12910 41794 12962 41806
rect 15038 41858 15090 41870
rect 15038 41794 15090 41806
rect 22990 41858 23042 41870
rect 22990 41794 23042 41806
rect 24446 41858 24498 41870
rect 27806 41858 27858 41870
rect 25442 41806 25454 41858
rect 25506 41806 25518 41858
rect 24446 41794 24498 41806
rect 27806 41794 27858 41806
rect 28254 41858 28306 41870
rect 28254 41794 28306 41806
rect 28814 41858 28866 41870
rect 28814 41794 28866 41806
rect 30942 41858 30994 41870
rect 30942 41794 30994 41806
rect 32286 41858 32338 41870
rect 35298 41806 35310 41858
rect 35362 41806 35374 41858
rect 32286 41794 32338 41806
rect 6974 41746 7026 41758
rect 31502 41746 31554 41758
rect 6626 41694 6638 41746
rect 6690 41694 6702 41746
rect 22418 41694 22430 41746
rect 22482 41694 22494 41746
rect 23874 41694 23886 41746
rect 23938 41694 23950 41746
rect 6974 41682 7026 41694
rect 31502 41682 31554 41694
rect 31838 41746 31890 41758
rect 31838 41682 31890 41694
rect 1344 41578 38640 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 38640 41578
rect 1344 41492 38640 41526
rect 22654 41410 22706 41422
rect 34974 41410 35026 41422
rect 29026 41358 29038 41410
rect 29090 41407 29102 41410
rect 29474 41407 29486 41410
rect 29090 41361 29486 41407
rect 29090 41358 29102 41361
rect 29474 41358 29486 41361
rect 29538 41358 29550 41410
rect 29698 41358 29710 41410
rect 29762 41407 29774 41410
rect 30146 41407 30158 41410
rect 29762 41361 30158 41407
rect 29762 41358 29774 41361
rect 30146 41358 30158 41361
rect 30210 41407 30222 41410
rect 30594 41407 30606 41410
rect 30210 41361 30606 41407
rect 30210 41358 30222 41361
rect 30594 41358 30606 41361
rect 30658 41358 30670 41410
rect 22654 41346 22706 41358
rect 34974 41346 35026 41358
rect 36430 41410 36482 41422
rect 36430 41346 36482 41358
rect 37438 41410 37490 41422
rect 37438 41346 37490 41358
rect 7198 41298 7250 41310
rect 22878 41298 22930 41310
rect 10770 41246 10782 41298
rect 10834 41246 10846 41298
rect 12898 41246 12910 41298
rect 12962 41246 12974 41298
rect 21410 41246 21422 41298
rect 21474 41246 21486 41298
rect 7198 41234 7250 41246
rect 22878 41234 22930 41246
rect 23326 41298 23378 41310
rect 27134 41298 27186 41310
rect 25106 41246 25118 41298
rect 25170 41246 25182 41298
rect 25890 41246 25902 41298
rect 25954 41246 25966 41298
rect 23326 41234 23378 41246
rect 27134 41234 27186 41246
rect 27470 41298 27522 41310
rect 27470 41234 27522 41246
rect 28366 41298 28418 41310
rect 28366 41234 28418 41246
rect 29262 41298 29314 41310
rect 29262 41234 29314 41246
rect 29710 41298 29762 41310
rect 29710 41234 29762 41246
rect 30158 41298 30210 41310
rect 30158 41234 30210 41246
rect 30606 41298 30658 41310
rect 30606 41234 30658 41246
rect 35310 41298 35362 41310
rect 35310 41234 35362 41246
rect 36094 41298 36146 41310
rect 36094 41234 36146 41246
rect 37102 41298 37154 41310
rect 37102 41234 37154 41246
rect 14814 41186 14866 41198
rect 21534 41186 21586 41198
rect 25454 41186 25506 41198
rect 38222 41186 38274 41198
rect 6514 41134 6526 41186
rect 6578 41134 6590 41186
rect 9986 41134 9998 41186
rect 10050 41134 10062 41186
rect 15026 41134 15038 41186
rect 15090 41134 15102 41186
rect 18498 41134 18510 41186
rect 18562 41134 18574 41186
rect 20738 41134 20750 41186
rect 20802 41134 20814 41186
rect 21298 41134 21310 41186
rect 21362 41134 21374 41186
rect 24770 41134 24782 41186
rect 24834 41134 24846 41186
rect 25666 41134 25678 41186
rect 25730 41134 25742 41186
rect 31490 41134 31502 41186
rect 31554 41134 31566 41186
rect 14814 41122 14866 41134
rect 21534 41122 21586 41134
rect 25454 41122 25506 41134
rect 38222 41122 38274 41134
rect 6750 41074 6802 41086
rect 6750 41010 6802 41022
rect 15598 41084 15650 41096
rect 15598 41020 15650 41032
rect 17502 41074 17554 41086
rect 17502 41010 17554 41022
rect 20078 41074 20130 41086
rect 20078 41010 20130 41022
rect 21982 41074 22034 41086
rect 21982 41010 22034 41022
rect 23774 41074 23826 41086
rect 23774 41010 23826 41022
rect 26574 41074 26626 41086
rect 26574 41010 26626 41022
rect 35534 41074 35586 41086
rect 35534 41010 35586 41022
rect 35870 41074 35922 41086
rect 35870 41010 35922 41022
rect 13582 40962 13634 40974
rect 13582 40898 13634 40910
rect 16494 40962 16546 40974
rect 21758 40962 21810 40974
rect 27918 40962 27970 40974
rect 17042 40910 17054 40962
rect 17106 40910 17118 40962
rect 22306 40910 22318 40962
rect 22370 40910 22382 40962
rect 16494 40898 16546 40910
rect 21758 40898 21810 40910
rect 27918 40898 27970 40910
rect 31726 40962 31778 40974
rect 31726 40898 31778 40910
rect 1344 40794 38640 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 38640 40794
rect 1344 40708 38640 40742
rect 6974 40626 7026 40638
rect 6974 40562 7026 40574
rect 13246 40626 13298 40638
rect 13246 40562 13298 40574
rect 16382 40626 16434 40638
rect 16382 40562 16434 40574
rect 16942 40626 16994 40638
rect 16942 40562 16994 40574
rect 17502 40626 17554 40638
rect 17502 40562 17554 40574
rect 22094 40626 22146 40638
rect 22094 40562 22146 40574
rect 22878 40626 22930 40638
rect 22878 40562 22930 40574
rect 23886 40626 23938 40638
rect 23886 40562 23938 40574
rect 24222 40626 24274 40638
rect 24222 40562 24274 40574
rect 24670 40626 24722 40638
rect 24670 40562 24722 40574
rect 25902 40626 25954 40638
rect 25902 40562 25954 40574
rect 26238 40626 26290 40638
rect 27582 40626 27634 40638
rect 26562 40574 26574 40626
rect 26626 40574 26638 40626
rect 26238 40562 26290 40574
rect 27582 40562 27634 40574
rect 28478 40626 28530 40638
rect 35310 40626 35362 40638
rect 29474 40574 29486 40626
rect 29538 40574 29550 40626
rect 30482 40574 30494 40626
rect 30546 40574 30558 40626
rect 28478 40562 28530 40574
rect 35310 40562 35362 40574
rect 35758 40626 35810 40638
rect 35758 40562 35810 40574
rect 38334 40626 38386 40638
rect 38334 40562 38386 40574
rect 4958 40514 5010 40526
rect 4958 40450 5010 40462
rect 5854 40514 5906 40526
rect 15150 40514 15202 40526
rect 13570 40462 13582 40514
rect 13634 40462 13646 40514
rect 14354 40462 14366 40514
rect 14418 40462 14430 40514
rect 5854 40450 5906 40462
rect 15150 40450 15202 40462
rect 17950 40514 18002 40526
rect 17950 40450 18002 40462
rect 20414 40514 20466 40526
rect 20414 40450 20466 40462
rect 20862 40514 20914 40526
rect 20862 40450 20914 40462
rect 21198 40514 21250 40526
rect 29586 40462 29598 40514
rect 29650 40462 29662 40514
rect 21198 40450 21250 40462
rect 4286 40402 4338 40414
rect 3938 40350 3950 40402
rect 4002 40350 4014 40402
rect 4286 40338 4338 40350
rect 4510 40402 4562 40414
rect 5630 40402 5682 40414
rect 5394 40350 5406 40402
rect 5458 40350 5470 40402
rect 4510 40338 4562 40350
rect 5630 40338 5682 40350
rect 5966 40402 6018 40414
rect 5966 40338 6018 40350
rect 6526 40402 6578 40414
rect 19182 40402 19234 40414
rect 9986 40350 9998 40402
rect 10050 40350 10062 40402
rect 17378 40350 17390 40402
rect 17442 40350 17454 40402
rect 29138 40350 29150 40402
rect 29202 40350 29214 40402
rect 30258 40350 30270 40402
rect 30322 40350 30334 40402
rect 6526 40338 6578 40350
rect 19182 40338 19234 40350
rect 5742 40290 5794 40302
rect 15374 40290 15426 40302
rect 10658 40238 10670 40290
rect 10722 40238 10734 40290
rect 12786 40238 12798 40290
rect 12850 40238 12862 40290
rect 5742 40226 5794 40238
rect 15374 40226 15426 40238
rect 22542 40290 22594 40302
rect 22542 40226 22594 40238
rect 23438 40290 23490 40302
rect 23438 40226 23490 40238
rect 25342 40290 25394 40302
rect 25342 40226 25394 40238
rect 27134 40290 27186 40302
rect 27134 40226 27186 40238
rect 28030 40290 28082 40302
rect 28030 40226 28082 40238
rect 37774 40290 37826 40302
rect 37774 40226 37826 40238
rect 15710 40178 15762 40190
rect 26910 40178 26962 40190
rect 23762 40126 23774 40178
rect 23826 40175 23838 40178
rect 24770 40175 24782 40178
rect 23826 40129 24782 40175
rect 23826 40126 23838 40129
rect 24770 40126 24782 40129
rect 24834 40126 24846 40178
rect 25330 40126 25342 40178
rect 25394 40175 25406 40178
rect 25778 40175 25790 40178
rect 25394 40129 25790 40175
rect 25394 40126 25406 40129
rect 25778 40126 25790 40129
rect 25842 40126 25854 40178
rect 15710 40114 15762 40126
rect 26910 40114 26962 40126
rect 1344 40010 38640 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 38640 40010
rect 1344 39924 38640 39958
rect 15598 39842 15650 39854
rect 22766 39842 22818 39854
rect 19506 39790 19518 39842
rect 19570 39839 19582 39842
rect 19954 39839 19966 39842
rect 19570 39793 19966 39839
rect 19570 39790 19582 39793
rect 19954 39790 19966 39793
rect 20018 39790 20030 39842
rect 15598 39778 15650 39790
rect 22766 39778 22818 39790
rect 23774 39842 23826 39854
rect 23774 39778 23826 39790
rect 24110 39842 24162 39854
rect 24110 39778 24162 39790
rect 29822 39842 29874 39854
rect 34302 39842 34354 39854
rect 33618 39790 33630 39842
rect 33682 39839 33694 39842
rect 34066 39839 34078 39842
rect 33682 39793 34078 39839
rect 33682 39790 33694 39793
rect 34066 39790 34078 39793
rect 34130 39790 34142 39842
rect 29822 39778 29874 39790
rect 34302 39778 34354 39790
rect 6750 39730 6802 39742
rect 6178 39678 6190 39730
rect 6242 39678 6254 39730
rect 6750 39666 6802 39678
rect 7198 39730 7250 39742
rect 7198 39666 7250 39678
rect 18510 39730 18562 39742
rect 18510 39666 18562 39678
rect 19966 39730 20018 39742
rect 19966 39666 20018 39678
rect 20302 39730 20354 39742
rect 20302 39666 20354 39678
rect 20862 39730 20914 39742
rect 29262 39730 29314 39742
rect 22194 39678 22206 39730
rect 22258 39678 22270 39730
rect 24434 39678 24446 39730
rect 24498 39678 24510 39730
rect 30370 39678 30382 39730
rect 30434 39678 30446 39730
rect 32498 39678 32510 39730
rect 32562 39678 32574 39730
rect 35746 39678 35758 39730
rect 35810 39678 35822 39730
rect 37874 39678 37886 39730
rect 37938 39678 37950 39730
rect 20862 39666 20914 39678
rect 29262 39666 29314 39678
rect 5854 39618 5906 39630
rect 3154 39566 3166 39618
rect 3218 39566 3230 39618
rect 4386 39566 4398 39618
rect 4450 39566 4462 39618
rect 5058 39566 5070 39618
rect 5122 39566 5134 39618
rect 5618 39566 5630 39618
rect 5682 39566 5694 39618
rect 5854 39554 5906 39566
rect 12910 39618 12962 39630
rect 18174 39618 18226 39630
rect 13794 39566 13806 39618
rect 13858 39566 13870 39618
rect 15138 39566 15150 39618
rect 15202 39566 15214 39618
rect 12910 39554 12962 39566
rect 18174 39554 18226 39566
rect 21870 39618 21922 39630
rect 21870 39554 21922 39566
rect 22654 39618 22706 39630
rect 22654 39554 22706 39566
rect 26462 39618 26514 39630
rect 33742 39618 33794 39630
rect 27010 39566 27022 39618
rect 27074 39566 27086 39618
rect 33170 39566 33182 39618
rect 33234 39566 33246 39618
rect 26462 39554 26514 39566
rect 33742 39554 33794 39566
rect 34526 39618 34578 39630
rect 34526 39554 34578 39566
rect 34974 39618 35026 39630
rect 34974 39554 35026 39566
rect 35310 39618 35362 39630
rect 35310 39554 35362 39566
rect 35870 39618 35922 39630
rect 35870 39554 35922 39566
rect 36094 39618 36146 39630
rect 36094 39554 36146 39566
rect 36206 39618 36258 39630
rect 37202 39566 37214 39618
rect 37266 39566 37278 39618
rect 36206 39554 36258 39566
rect 17726 39506 17778 39518
rect 15026 39454 15038 39506
rect 15090 39454 15102 39506
rect 17726 39442 17778 39454
rect 21646 39506 21698 39518
rect 21646 39442 21698 39454
rect 23662 39506 23714 39518
rect 23662 39442 23714 39454
rect 24334 39506 24386 39518
rect 27470 39506 27522 39518
rect 24882 39454 24894 39506
rect 24946 39454 24958 39506
rect 24334 39442 24386 39454
rect 27470 39442 27522 39454
rect 29934 39506 29986 39518
rect 35186 39454 35198 39506
rect 35250 39454 35262 39506
rect 29934 39442 29986 39454
rect 2942 39394 2994 39406
rect 2942 39330 2994 39342
rect 4622 39394 4674 39406
rect 4622 39330 4674 39342
rect 4734 39394 4786 39406
rect 4734 39330 4786 39342
rect 4846 39394 4898 39406
rect 4846 39330 4898 39342
rect 6078 39394 6130 39406
rect 6078 39330 6130 39342
rect 6190 39394 6242 39406
rect 6190 39330 6242 39342
rect 12462 39394 12514 39406
rect 12462 39330 12514 39342
rect 14030 39394 14082 39406
rect 16382 39394 16434 39406
rect 14914 39342 14926 39394
rect 14978 39342 14990 39394
rect 14030 39330 14082 39342
rect 16382 39330 16434 39342
rect 18174 39394 18226 39406
rect 18174 39330 18226 39342
rect 22094 39394 22146 39406
rect 22094 39330 22146 39342
rect 22206 39394 22258 39406
rect 22206 39330 22258 39342
rect 22766 39394 22818 39406
rect 22766 39330 22818 39342
rect 23326 39394 23378 39406
rect 35758 39394 35810 39406
rect 28466 39342 28478 39394
rect 28530 39342 28542 39394
rect 23326 39330 23378 39342
rect 35758 39330 35810 39342
rect 1344 39226 38640 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 38640 39226
rect 1344 39140 38640 39174
rect 5182 39058 5234 39070
rect 5182 38994 5234 39006
rect 5518 39058 5570 39070
rect 5518 38994 5570 39006
rect 10446 39058 10498 39070
rect 10446 38994 10498 39006
rect 13022 39058 13074 39070
rect 13022 38994 13074 39006
rect 18398 39058 18450 39070
rect 18398 38994 18450 39006
rect 22990 39058 23042 39070
rect 22990 38994 23042 39006
rect 24110 39058 24162 39070
rect 24110 38994 24162 39006
rect 24222 39058 24274 39070
rect 24222 38994 24274 39006
rect 31390 39058 31442 39070
rect 33618 39006 33630 39058
rect 33682 39006 33694 39058
rect 31390 38994 31442 39006
rect 6862 38946 6914 38958
rect 2482 38894 2494 38946
rect 2546 38894 2558 38946
rect 5954 38894 5966 38946
rect 6018 38894 6030 38946
rect 6290 38894 6302 38946
rect 6354 38894 6366 38946
rect 6862 38882 6914 38894
rect 17390 38946 17442 38958
rect 17390 38882 17442 38894
rect 17726 38946 17778 38958
rect 23326 38946 23378 38958
rect 21634 38894 21646 38946
rect 21698 38894 21710 38946
rect 17726 38882 17778 38894
rect 23326 38882 23378 38894
rect 24334 38946 24386 38958
rect 24334 38882 24386 38894
rect 25230 38946 25282 38958
rect 30606 38946 30658 38958
rect 26002 38894 26014 38946
rect 26066 38894 26078 38946
rect 25230 38882 25282 38894
rect 30606 38882 30658 38894
rect 32398 38946 32450 38958
rect 32398 38882 32450 38894
rect 5854 38834 5906 38846
rect 10110 38834 10162 38846
rect 19182 38834 19234 38846
rect 1810 38782 1822 38834
rect 1874 38782 1886 38834
rect 6402 38782 6414 38834
rect 6466 38782 6478 38834
rect 16258 38782 16270 38834
rect 16322 38782 16334 38834
rect 23998 38834 24050 38846
rect 26238 38834 26290 38846
rect 31838 38834 31890 38846
rect 5854 38770 5906 38782
rect 10110 38770 10162 38782
rect 19182 38770 19234 38782
rect 22306 38770 22318 38822
rect 22370 38770 22382 38822
rect 24546 38782 24558 38834
rect 24610 38782 24622 38834
rect 25778 38782 25790 38834
rect 25842 38782 25854 38834
rect 26450 38782 26462 38834
rect 26514 38782 26526 38834
rect 27234 38782 27246 38834
rect 27298 38782 27310 38834
rect 32162 38782 32174 38834
rect 32226 38782 32238 38834
rect 38098 38782 38110 38834
rect 38162 38782 38174 38834
rect 23998 38770 24050 38782
rect 26238 38770 26290 38782
rect 31838 38770 31890 38782
rect 16830 38722 16882 38734
rect 18958 38722 19010 38734
rect 32510 38722 32562 38734
rect 4610 38670 4622 38722
rect 4674 38670 4686 38722
rect 13346 38670 13358 38722
rect 13410 38670 13422 38722
rect 15474 38670 15486 38722
rect 15538 38670 15550 38722
rect 18610 38670 18622 38722
rect 18674 38670 18686 38722
rect 19506 38670 19518 38722
rect 19570 38670 19582 38722
rect 28018 38670 28030 38722
rect 28082 38670 28094 38722
rect 30146 38670 30158 38722
rect 30210 38670 30222 38722
rect 16830 38658 16882 38670
rect 18958 38658 19010 38670
rect 32510 38658 32562 38670
rect 33070 38722 33122 38734
rect 35298 38670 35310 38722
rect 35362 38670 35374 38722
rect 37426 38670 37438 38722
rect 37490 38670 37502 38722
rect 33070 38658 33122 38670
rect 33294 38610 33346 38622
rect 17938 38558 17950 38610
rect 18002 38607 18014 38610
rect 18386 38607 18398 38610
rect 18002 38561 18398 38607
rect 18002 38558 18014 38561
rect 18386 38558 18398 38561
rect 18450 38558 18462 38610
rect 33294 38546 33346 38558
rect 1344 38442 38640 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 38640 38442
rect 1344 38356 38640 38390
rect 26450 38222 26462 38274
rect 26514 38271 26526 38274
rect 26898 38271 26910 38274
rect 26514 38225 26910 38271
rect 26514 38222 26526 38225
rect 26898 38222 26910 38225
rect 26962 38222 26974 38274
rect 4846 38162 4898 38174
rect 4846 38098 4898 38110
rect 5742 38162 5794 38174
rect 14814 38162 14866 38174
rect 16382 38162 16434 38174
rect 26462 38162 26514 38174
rect 38222 38162 38274 38174
rect 7410 38110 7422 38162
rect 7474 38110 7486 38162
rect 15922 38110 15934 38162
rect 15986 38110 15998 38162
rect 18386 38110 18398 38162
rect 18450 38110 18462 38162
rect 20514 38110 20526 38162
rect 20578 38110 20590 38162
rect 22194 38110 22206 38162
rect 22258 38110 22270 38162
rect 23090 38110 23102 38162
rect 23154 38110 23166 38162
rect 25218 38110 25230 38162
rect 25282 38110 25294 38162
rect 30482 38110 30494 38162
rect 30546 38110 30558 38162
rect 35522 38110 35534 38162
rect 35586 38110 35598 38162
rect 5742 38098 5794 38110
rect 14814 38098 14866 38110
rect 16382 38098 16434 38110
rect 26462 38098 26514 38110
rect 38222 38098 38274 38110
rect 4622 38050 4674 38062
rect 11454 38050 11506 38062
rect 10210 37998 10222 38050
rect 10274 37998 10286 38050
rect 4622 37986 4674 37998
rect 11454 37986 11506 37998
rect 14590 38050 14642 38062
rect 14590 37986 14642 37998
rect 15822 38050 15874 38062
rect 37774 38050 37826 38062
rect 17042 37998 17054 38050
rect 17106 37998 17118 38050
rect 17714 37998 17726 38050
rect 17778 37998 17790 38050
rect 22306 37998 22318 38050
rect 22370 37998 22382 38050
rect 26002 37998 26014 38050
rect 26066 37998 26078 38050
rect 33394 37998 33406 38050
rect 33458 37998 33470 38050
rect 36418 37998 36430 38050
rect 36482 37998 36494 38050
rect 15822 37986 15874 37998
rect 37774 37986 37826 37998
rect 3278 37938 3330 37950
rect 10670 37938 10722 37950
rect 9538 37886 9550 37938
rect 9602 37886 9614 37938
rect 3278 37874 3330 37886
rect 10670 37874 10722 37886
rect 11006 37938 11058 37950
rect 11006 37874 11058 37886
rect 15374 37938 15426 37950
rect 15374 37874 15426 37886
rect 16606 37938 16658 37950
rect 21646 37938 21698 37950
rect 16818 37886 16830 37938
rect 16882 37886 16894 37938
rect 16606 37874 16658 37886
rect 21646 37874 21698 37886
rect 21870 37938 21922 37950
rect 36990 37938 37042 37950
rect 32610 37886 32622 37938
rect 32674 37886 32686 37938
rect 21870 37874 21922 37886
rect 36990 37874 37042 37886
rect 37326 37938 37378 37950
rect 37326 37874 37378 37886
rect 2942 37826 2994 37838
rect 13918 37826 13970 37838
rect 15598 37826 15650 37838
rect 4274 37774 4286 37826
rect 4338 37774 4350 37826
rect 14242 37774 14254 37826
rect 14306 37774 14318 37826
rect 2942 37762 2994 37774
rect 13918 37762 13970 37774
rect 15598 37762 15650 37774
rect 15934 37826 15986 37838
rect 15934 37762 15986 37774
rect 17390 37826 17442 37838
rect 17390 37762 17442 37774
rect 22094 37826 22146 37838
rect 22094 37762 22146 37774
rect 22766 37826 22818 37838
rect 22766 37762 22818 37774
rect 26910 37826 26962 37838
rect 26910 37762 26962 37774
rect 33854 37826 33906 37838
rect 33854 37762 33906 37774
rect 1344 37658 38640 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 38640 37658
rect 1344 37572 38640 37606
rect 5070 37490 5122 37502
rect 10558 37490 10610 37502
rect 10098 37438 10110 37490
rect 10162 37438 10174 37490
rect 5070 37426 5122 37438
rect 10558 37426 10610 37438
rect 15374 37490 15426 37502
rect 15374 37426 15426 37438
rect 15710 37490 15762 37502
rect 15710 37426 15762 37438
rect 16606 37490 16658 37502
rect 16606 37426 16658 37438
rect 18286 37490 18338 37502
rect 18286 37426 18338 37438
rect 19518 37490 19570 37502
rect 21870 37490 21922 37502
rect 20738 37438 20750 37490
rect 20802 37438 20814 37490
rect 19518 37426 19570 37438
rect 21870 37426 21922 37438
rect 23438 37490 23490 37502
rect 23438 37426 23490 37438
rect 23886 37490 23938 37502
rect 23886 37426 23938 37438
rect 24334 37490 24386 37502
rect 24334 37426 24386 37438
rect 25790 37490 25842 37502
rect 25790 37426 25842 37438
rect 28254 37490 28306 37502
rect 28254 37426 28306 37438
rect 28926 37490 28978 37502
rect 28926 37426 28978 37438
rect 13470 37378 13522 37390
rect 2482 37326 2494 37378
rect 2546 37326 2558 37378
rect 13470 37314 13522 37326
rect 13806 37378 13858 37390
rect 13806 37314 13858 37326
rect 16046 37378 16098 37390
rect 16046 37314 16098 37326
rect 22430 37378 22482 37390
rect 22430 37314 22482 37326
rect 27806 37378 27858 37390
rect 27806 37314 27858 37326
rect 28142 37378 28194 37390
rect 28142 37314 28194 37326
rect 5518 37266 5570 37278
rect 1810 37214 1822 37266
rect 1874 37214 1886 37266
rect 5518 37202 5570 37214
rect 5630 37266 5682 37278
rect 5630 37202 5682 37214
rect 5742 37266 5794 37278
rect 9774 37266 9826 37278
rect 5954 37214 5966 37266
rect 6018 37214 6030 37266
rect 5742 37202 5794 37214
rect 9774 37202 9826 37214
rect 12574 37266 12626 37278
rect 12574 37202 12626 37214
rect 22654 37266 22706 37278
rect 28466 37214 28478 37266
rect 28530 37214 28542 37266
rect 38210 37214 38222 37266
rect 38274 37214 38286 37266
rect 22654 37202 22706 37214
rect 6750 37154 6802 37166
rect 4610 37102 4622 37154
rect 4674 37102 4686 37154
rect 6750 37090 6802 37102
rect 9550 37154 9602 37166
rect 9550 37090 9602 37102
rect 11678 37154 11730 37166
rect 11678 37090 11730 37102
rect 13022 37154 13074 37166
rect 13022 37090 13074 37102
rect 17726 37154 17778 37166
rect 17726 37090 17778 37102
rect 19966 37154 20018 37166
rect 19966 37090 20018 37102
rect 20526 37154 20578 37166
rect 20526 37090 20578 37102
rect 21310 37154 21362 37166
rect 21310 37090 21362 37102
rect 25342 37154 25394 37166
rect 25342 37090 25394 37102
rect 31614 37154 31666 37166
rect 35298 37102 35310 37154
rect 35362 37102 35374 37154
rect 37426 37102 37438 37154
rect 37490 37102 37502 37154
rect 31614 37090 31666 37102
rect 6414 37042 6466 37054
rect 12350 37042 12402 37054
rect 12002 36990 12014 37042
rect 12066 36990 12078 37042
rect 6414 36978 6466 36990
rect 12350 36978 12402 36990
rect 21086 37042 21138 37054
rect 21086 36978 21138 36990
rect 22990 37042 23042 37054
rect 22990 36978 23042 36990
rect 1344 36874 38640 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 38640 36874
rect 1344 36788 38640 36822
rect 22642 36654 22654 36706
rect 22706 36703 22718 36706
rect 23314 36703 23326 36706
rect 22706 36657 23326 36703
rect 22706 36654 22718 36657
rect 23314 36654 23326 36657
rect 23378 36654 23390 36706
rect 37538 36654 37550 36706
rect 37602 36654 37614 36706
rect 5182 36594 5234 36606
rect 5182 36530 5234 36542
rect 5966 36594 6018 36606
rect 5966 36530 6018 36542
rect 6750 36594 6802 36606
rect 6750 36530 6802 36542
rect 8542 36594 8594 36606
rect 8542 36530 8594 36542
rect 15150 36594 15202 36606
rect 15150 36530 15202 36542
rect 16606 36594 16658 36606
rect 16606 36530 16658 36542
rect 17278 36594 17330 36606
rect 17278 36530 17330 36542
rect 18510 36594 18562 36606
rect 18510 36530 18562 36542
rect 22766 36594 22818 36606
rect 22766 36530 22818 36542
rect 23102 36594 23154 36606
rect 38222 36594 38274 36606
rect 28130 36542 28142 36594
rect 28194 36542 28206 36594
rect 23102 36530 23154 36542
rect 38222 36530 38274 36542
rect 5854 36482 5906 36494
rect 5854 36418 5906 36430
rect 6078 36482 6130 36494
rect 6078 36418 6130 36430
rect 8990 36482 9042 36494
rect 8990 36418 9042 36430
rect 9102 36482 9154 36494
rect 23998 36482 24050 36494
rect 29150 36482 29202 36494
rect 31054 36482 31106 36494
rect 36990 36482 37042 36494
rect 9426 36430 9438 36482
rect 9490 36430 9502 36482
rect 11666 36430 11678 36482
rect 11730 36430 11742 36482
rect 25218 36430 25230 36482
rect 25282 36430 25294 36482
rect 30146 36430 30158 36482
rect 30210 36430 30222 36482
rect 31826 36430 31838 36482
rect 31890 36430 31902 36482
rect 36194 36430 36206 36482
rect 36258 36430 36270 36482
rect 9102 36418 9154 36430
rect 23998 36418 24050 36430
rect 29150 36418 29202 36430
rect 31054 36418 31106 36430
rect 36990 36418 37042 36430
rect 37214 36482 37266 36494
rect 37214 36418 37266 36430
rect 5630 36370 5682 36382
rect 5630 36306 5682 36318
rect 9214 36370 9266 36382
rect 9214 36306 9266 36318
rect 24334 36370 24386 36382
rect 36430 36370 36482 36382
rect 26002 36318 26014 36370
rect 26066 36318 26078 36370
rect 24334 36306 24386 36318
rect 36430 36306 36482 36318
rect 6190 36258 6242 36270
rect 6190 36194 6242 36206
rect 7198 36258 7250 36270
rect 7198 36194 7250 36206
rect 9886 36258 9938 36270
rect 9886 36194 9938 36206
rect 11454 36258 11506 36270
rect 11454 36194 11506 36206
rect 21534 36258 21586 36270
rect 21534 36194 21586 36206
rect 22206 36258 22258 36270
rect 22206 36194 22258 36206
rect 23550 36258 23602 36270
rect 23550 36194 23602 36206
rect 28590 36258 28642 36270
rect 32846 36258 32898 36270
rect 30930 36206 30942 36258
rect 30994 36206 31006 36258
rect 28590 36194 28642 36206
rect 32846 36194 32898 36206
rect 35758 36258 35810 36270
rect 35758 36194 35810 36206
rect 1344 36090 38640 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 38640 36090
rect 1344 36004 38640 36038
rect 9774 35922 9826 35934
rect 9774 35858 9826 35870
rect 9886 35922 9938 35934
rect 9886 35858 9938 35870
rect 10670 35922 10722 35934
rect 10670 35858 10722 35870
rect 15710 35922 15762 35934
rect 15710 35858 15762 35870
rect 20526 35922 20578 35934
rect 20526 35858 20578 35870
rect 20862 35922 20914 35934
rect 20862 35858 20914 35870
rect 23326 35922 23378 35934
rect 31054 35922 31106 35934
rect 28690 35870 28702 35922
rect 28754 35870 28766 35922
rect 23326 35858 23378 35870
rect 31054 35858 31106 35870
rect 31166 35922 31218 35934
rect 31166 35858 31218 35870
rect 35086 35922 35138 35934
rect 36418 35870 36430 35922
rect 36482 35870 36494 35922
rect 35086 35858 35138 35870
rect 4174 35810 4226 35822
rect 4174 35746 4226 35758
rect 7310 35810 7362 35822
rect 7310 35746 7362 35758
rect 9550 35810 9602 35822
rect 19742 35810 19794 35822
rect 26686 35810 26738 35822
rect 30606 35810 30658 35822
rect 12786 35758 12798 35810
rect 12850 35758 12862 35810
rect 17490 35758 17502 35810
rect 17554 35758 17566 35810
rect 17826 35758 17838 35810
rect 17890 35758 17902 35810
rect 19954 35758 19966 35810
rect 20018 35758 20030 35810
rect 28914 35758 28926 35810
rect 28978 35758 28990 35810
rect 9550 35746 9602 35758
rect 19742 35746 19794 35758
rect 26686 35746 26738 35758
rect 30606 35746 30658 35758
rect 3950 35698 4002 35710
rect 3950 35634 4002 35646
rect 4510 35698 4562 35710
rect 4510 35634 4562 35646
rect 4734 35698 4786 35710
rect 4734 35634 4786 35646
rect 5518 35698 5570 35710
rect 5518 35634 5570 35646
rect 6974 35698 7026 35710
rect 6974 35634 7026 35646
rect 9998 35698 10050 35710
rect 9998 35634 10050 35646
rect 10110 35698 10162 35710
rect 10110 35634 10162 35646
rect 11118 35698 11170 35710
rect 15598 35698 15650 35710
rect 12002 35646 12014 35698
rect 12066 35646 12078 35698
rect 11118 35634 11170 35646
rect 15598 35634 15650 35646
rect 15934 35698 15986 35710
rect 19518 35698 19570 35710
rect 27022 35698 27074 35710
rect 30830 35698 30882 35710
rect 16146 35646 16158 35698
rect 16210 35646 16222 35698
rect 17938 35646 17950 35698
rect 18002 35646 18014 35698
rect 20066 35646 20078 35698
rect 20130 35646 20142 35698
rect 28242 35646 28254 35698
rect 28306 35646 28318 35698
rect 29138 35646 29150 35698
rect 29202 35646 29214 35698
rect 15934 35634 15986 35646
rect 19518 35634 19570 35646
rect 27022 35634 27074 35646
rect 30830 35634 30882 35646
rect 32398 35698 32450 35710
rect 32398 35634 32450 35646
rect 6638 35586 6690 35598
rect 15822 35586 15874 35598
rect 14914 35534 14926 35586
rect 14978 35534 14990 35586
rect 6638 35522 6690 35534
rect 15822 35522 15874 35534
rect 17390 35586 17442 35598
rect 17390 35522 17442 35534
rect 18734 35586 18786 35598
rect 18734 35522 18786 35534
rect 19294 35586 19346 35598
rect 19294 35522 19346 35534
rect 30942 35586 30994 35598
rect 30942 35522 30994 35534
rect 33182 35586 33234 35598
rect 33182 35522 33234 35534
rect 35534 35586 35586 35598
rect 35534 35522 35586 35534
rect 36094 35586 36146 35598
rect 36094 35522 36146 35534
rect 36766 35586 36818 35598
rect 36766 35522 36818 35534
rect 36990 35586 37042 35598
rect 36990 35522 37042 35534
rect 3614 35474 3666 35486
rect 18398 35474 18450 35486
rect 32174 35474 32226 35486
rect 5058 35422 5070 35474
rect 5122 35422 5134 35474
rect 10770 35422 10782 35474
rect 10834 35471 10846 35474
rect 11218 35471 11230 35474
rect 10834 35425 11230 35471
rect 10834 35422 10846 35425
rect 11218 35422 11230 35425
rect 11282 35422 11294 35474
rect 18610 35422 18622 35474
rect 18674 35471 18686 35474
rect 19282 35471 19294 35474
rect 18674 35425 19294 35471
rect 18674 35422 18686 35425
rect 19282 35422 19294 35425
rect 19346 35422 19358 35474
rect 31826 35422 31838 35474
rect 31890 35422 31902 35474
rect 35522 35422 35534 35474
rect 35586 35471 35598 35474
rect 36194 35471 36206 35474
rect 35586 35425 36206 35471
rect 35586 35422 35598 35425
rect 36194 35422 36206 35425
rect 36258 35422 36270 35474
rect 3614 35410 3666 35422
rect 18398 35410 18450 35422
rect 32174 35410 32226 35422
rect 1344 35306 38640 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 38640 35306
rect 1344 35220 38640 35254
rect 28478 35138 28530 35150
rect 28478 35074 28530 35086
rect 4398 35026 4450 35038
rect 15374 35026 15426 35038
rect 7522 34974 7534 35026
rect 7586 34974 7598 35026
rect 9650 34974 9662 35026
rect 9714 34974 9726 35026
rect 10770 34974 10782 35026
rect 10834 34974 10846 35026
rect 12898 34974 12910 35026
rect 12962 34974 12974 35026
rect 4398 34962 4450 34974
rect 15374 34962 15426 34974
rect 19630 35026 19682 35038
rect 22194 34974 22206 35026
rect 22258 34974 22270 35026
rect 34850 34974 34862 35026
rect 34914 34974 34926 35026
rect 35634 34974 35646 35026
rect 35698 34974 35710 35026
rect 19630 34962 19682 34974
rect 3278 34914 3330 34926
rect 3278 34850 3330 34862
rect 5854 34914 5906 34926
rect 5854 34850 5906 34862
rect 5966 34914 6018 34926
rect 5966 34850 6018 34862
rect 6302 34914 6354 34926
rect 15150 34914 15202 34926
rect 6738 34862 6750 34914
rect 6802 34862 6814 34914
rect 10098 34862 10110 34914
rect 10162 34862 10174 34914
rect 6302 34850 6354 34862
rect 15150 34850 15202 34862
rect 17838 34914 17890 34926
rect 17838 34850 17890 34862
rect 18622 34914 18674 34926
rect 25566 34914 25618 34926
rect 25106 34862 25118 34914
rect 25170 34862 25182 34914
rect 18622 34850 18674 34862
rect 25566 34850 25618 34862
rect 30270 34914 30322 34926
rect 35870 34914 35922 34926
rect 31378 34862 31390 34914
rect 31442 34862 31454 34914
rect 31938 34862 31950 34914
rect 32002 34862 32014 34914
rect 30270 34850 30322 34862
rect 35870 34850 35922 34862
rect 35982 34914 36034 34926
rect 35982 34850 36034 34862
rect 18062 34802 18114 34814
rect 18062 34738 18114 34750
rect 18174 34802 18226 34814
rect 28590 34802 28642 34814
rect 24322 34750 24334 34802
rect 24386 34750 24398 34802
rect 18174 34738 18226 34750
rect 28590 34738 28642 34750
rect 31614 34802 31666 34814
rect 35534 34802 35586 34814
rect 32722 34750 32734 34802
rect 32786 34750 32798 34802
rect 31614 34738 31666 34750
rect 35534 34738 35586 34750
rect 2942 34690 2994 34702
rect 2942 34626 2994 34638
rect 6078 34690 6130 34702
rect 6078 34626 6130 34638
rect 6190 34690 6242 34702
rect 6190 34626 6242 34638
rect 13582 34690 13634 34702
rect 15822 34690 15874 34702
rect 14802 34638 14814 34690
rect 14866 34638 14878 34690
rect 13582 34626 13634 34638
rect 15822 34626 15874 34638
rect 18846 34690 18898 34702
rect 18846 34626 18898 34638
rect 19182 34690 19234 34702
rect 19182 34626 19234 34638
rect 35646 34690 35698 34702
rect 35646 34626 35698 34638
rect 1344 34522 38640 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 38640 34522
rect 1344 34436 38640 34470
rect 6974 34354 7026 34366
rect 6974 34290 7026 34302
rect 7422 34354 7474 34366
rect 7422 34290 7474 34302
rect 17726 34354 17778 34366
rect 17726 34290 17778 34302
rect 19630 34354 19682 34366
rect 19630 34290 19682 34302
rect 22990 34354 23042 34366
rect 22990 34290 23042 34302
rect 24558 34354 24610 34366
rect 24558 34290 24610 34302
rect 27022 34354 27074 34366
rect 31950 34354 32002 34366
rect 29362 34302 29374 34354
rect 29426 34302 29438 34354
rect 27022 34290 27074 34302
rect 31950 34290 32002 34302
rect 33406 34354 33458 34366
rect 33406 34290 33458 34302
rect 33742 34354 33794 34366
rect 33742 34290 33794 34302
rect 34078 34354 34130 34366
rect 34078 34290 34130 34302
rect 34526 34354 34578 34366
rect 34526 34290 34578 34302
rect 4958 34242 5010 34254
rect 2482 34190 2494 34242
rect 2546 34190 2558 34242
rect 4958 34178 5010 34190
rect 15038 34242 15090 34254
rect 15038 34178 15090 34190
rect 15374 34242 15426 34254
rect 15374 34178 15426 34190
rect 18622 34242 18674 34254
rect 31278 34242 31330 34254
rect 27346 34190 27358 34242
rect 27410 34190 27422 34242
rect 31042 34190 31054 34242
rect 31106 34190 31118 34242
rect 18622 34178 18674 34190
rect 31278 34178 31330 34190
rect 35198 34242 35250 34254
rect 35410 34190 35422 34242
rect 35474 34190 35486 34242
rect 35198 34178 35250 34190
rect 6078 34130 6130 34142
rect 1810 34078 1822 34130
rect 1874 34078 1886 34130
rect 5170 34078 5182 34130
rect 5234 34078 5246 34130
rect 6078 34066 6130 34078
rect 6190 34130 6242 34142
rect 6190 34066 6242 34078
rect 6302 34130 6354 34142
rect 7758 34130 7810 34142
rect 6514 34078 6526 34130
rect 6578 34078 6590 34130
rect 6302 34066 6354 34078
rect 7758 34066 7810 34078
rect 13134 34130 13186 34142
rect 17614 34130 17666 34142
rect 17378 34078 17390 34130
rect 17442 34078 17454 34130
rect 13134 34066 13186 34078
rect 17614 34066 17666 34078
rect 17838 34130 17890 34142
rect 17838 34066 17890 34078
rect 17950 34130 18002 34142
rect 19518 34130 19570 34142
rect 18834 34078 18846 34130
rect 18898 34078 18910 34130
rect 19282 34078 19294 34130
rect 19346 34078 19358 34130
rect 17950 34066 18002 34078
rect 19518 34066 19570 34078
rect 19742 34130 19794 34142
rect 19742 34066 19794 34078
rect 19854 34130 19906 34142
rect 19854 34066 19906 34078
rect 23550 34130 23602 34142
rect 24222 34130 24274 34142
rect 33854 34130 33906 34142
rect 34750 34130 34802 34142
rect 23874 34078 23886 34130
rect 23938 34078 23950 34130
rect 28466 34078 28478 34130
rect 28530 34078 28542 34130
rect 29138 34078 29150 34130
rect 29202 34078 29214 34130
rect 29474 34078 29486 34130
rect 29538 34078 29550 34130
rect 31490 34078 31502 34130
rect 31554 34078 31566 34130
rect 34290 34078 34302 34130
rect 34354 34078 34366 34130
rect 23550 34066 23602 34078
rect 24222 34066 24274 34078
rect 33854 34066 33906 34078
rect 34750 34066 34802 34078
rect 9886 34018 9938 34030
rect 4610 33966 4622 34018
rect 4674 33966 4686 34018
rect 9886 33954 9938 33966
rect 12238 34018 12290 34030
rect 12238 33954 12290 33966
rect 20974 34018 21026 34030
rect 20974 33954 21026 33966
rect 23326 34018 23378 34030
rect 23326 33954 23378 33966
rect 30942 34018 30994 34030
rect 30942 33954 30994 33966
rect 33966 34018 34018 34030
rect 33966 33954 34018 33966
rect 35534 34018 35586 34030
rect 35534 33954 35586 33966
rect 12910 33906 12962 33918
rect 12562 33854 12574 33906
rect 12626 33854 12638 33906
rect 12910 33842 12962 33854
rect 1344 33738 38640 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 38640 33738
rect 1344 33652 38640 33686
rect 6526 33570 6578 33582
rect 27022 33570 27074 33582
rect 4722 33518 4734 33570
rect 4786 33567 4798 33570
rect 4946 33567 4958 33570
rect 4786 33521 4958 33567
rect 4786 33518 4798 33521
rect 4946 33518 4958 33521
rect 5010 33518 5022 33570
rect 26338 33518 26350 33570
rect 26402 33567 26414 33570
rect 26786 33567 26798 33570
rect 26402 33521 26798 33567
rect 26402 33518 26414 33521
rect 26786 33518 26798 33521
rect 26850 33518 26862 33570
rect 6526 33506 6578 33518
rect 27022 33506 27074 33518
rect 27694 33570 27746 33582
rect 27694 33506 27746 33518
rect 29262 33570 29314 33582
rect 29262 33506 29314 33518
rect 33070 33570 33122 33582
rect 33070 33506 33122 33518
rect 5966 33458 6018 33470
rect 5966 33394 6018 33406
rect 7422 33458 7474 33470
rect 21870 33458 21922 33470
rect 15250 33406 15262 33458
rect 15314 33406 15326 33458
rect 17378 33406 17390 33458
rect 17442 33406 17454 33458
rect 18610 33406 18622 33458
rect 18674 33406 18686 33458
rect 20738 33406 20750 33458
rect 20802 33406 20814 33458
rect 7422 33394 7474 33406
rect 21870 33394 21922 33406
rect 26350 33458 26402 33470
rect 26350 33394 26402 33406
rect 26798 33458 26850 33470
rect 26798 33394 26850 33406
rect 31278 33458 31330 33470
rect 31278 33394 31330 33406
rect 35310 33458 35362 33470
rect 35310 33394 35362 33406
rect 6190 33346 6242 33358
rect 6190 33282 6242 33294
rect 6974 33346 7026 33358
rect 21646 33346 21698 33358
rect 31502 33346 31554 33358
rect 12562 33294 12574 33346
rect 12626 33294 12638 33346
rect 14578 33294 14590 33346
rect 14642 33294 14654 33346
rect 17826 33294 17838 33346
rect 17890 33294 17902 33346
rect 27346 33294 27358 33346
rect 27410 33294 27422 33346
rect 28018 33294 28030 33346
rect 28082 33294 28094 33346
rect 6974 33282 7026 33294
rect 21646 33282 21698 33294
rect 31502 33282 31554 33294
rect 33294 33346 33346 33358
rect 33294 33282 33346 33294
rect 33742 33346 33794 33358
rect 33742 33282 33794 33294
rect 34078 33346 34130 33358
rect 34078 33282 34130 33294
rect 34974 33346 35026 33358
rect 34974 33282 35026 33294
rect 35534 33346 35586 33358
rect 35534 33282 35586 33294
rect 28478 33234 28530 33246
rect 28478 33170 28530 33182
rect 29150 33234 29202 33246
rect 29150 33170 29202 33182
rect 32174 33234 32226 33246
rect 32174 33170 32226 33182
rect 32510 33234 32562 33246
rect 36990 33234 37042 33246
rect 33954 33182 33966 33234
rect 34018 33182 34030 33234
rect 35858 33182 35870 33234
rect 35922 33182 35934 33234
rect 32510 33170 32562 33182
rect 36990 33170 37042 33182
rect 4846 33122 4898 33134
rect 4846 33058 4898 33070
rect 12798 33122 12850 33134
rect 24110 33122 24162 33134
rect 21298 33070 21310 33122
rect 21362 33070 21374 33122
rect 12798 33058 12850 33070
rect 24110 33058 24162 33070
rect 27134 33122 27186 33134
rect 27134 33058 27186 33070
rect 27806 33122 27858 33134
rect 27806 33058 27858 33070
rect 30942 33122 30994 33134
rect 37326 33122 37378 33134
rect 31826 33070 31838 33122
rect 31890 33070 31902 33122
rect 30942 33058 30994 33070
rect 37326 33058 37378 33070
rect 1344 32954 38640 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 38640 32954
rect 1344 32868 38640 32902
rect 16830 32786 16882 32798
rect 16830 32722 16882 32734
rect 17502 32786 17554 32798
rect 18386 32734 18398 32786
rect 18450 32734 18462 32786
rect 17502 32722 17554 32734
rect 8094 32674 8146 32686
rect 21422 32674 21474 32686
rect 33070 32674 33122 32686
rect 4610 32622 4622 32674
rect 4674 32622 4686 32674
rect 12562 32622 12574 32674
rect 12626 32622 12638 32674
rect 27570 32622 27582 32674
rect 27634 32622 27646 32674
rect 8094 32610 8146 32622
rect 21422 32610 21474 32622
rect 33070 32610 33122 32622
rect 33406 32674 33458 32686
rect 37426 32622 37438 32674
rect 37490 32622 37502 32674
rect 33406 32610 33458 32622
rect 7310 32562 7362 32574
rect 15150 32562 15202 32574
rect 3938 32510 3950 32562
rect 4002 32510 4014 32562
rect 11778 32510 11790 32562
rect 11842 32510 11854 32562
rect 7310 32498 7362 32510
rect 15150 32498 15202 32510
rect 17838 32562 17890 32574
rect 21186 32510 21198 32562
rect 21250 32510 21262 32562
rect 26898 32510 26910 32562
rect 26962 32510 26974 32562
rect 38210 32510 38222 32562
rect 38274 32510 38286 32562
rect 17838 32498 17890 32510
rect 7086 32450 7138 32462
rect 30158 32450 30210 32462
rect 6738 32398 6750 32450
rect 6802 32398 6814 32450
rect 14690 32398 14702 32450
rect 14754 32398 14766 32450
rect 29698 32398 29710 32450
rect 29762 32398 29774 32450
rect 35298 32398 35310 32450
rect 35362 32398 35374 32450
rect 7086 32386 7138 32398
rect 30158 32386 30210 32398
rect 18062 32338 18114 32350
rect 7634 32286 7646 32338
rect 7698 32286 7710 32338
rect 18062 32274 18114 32286
rect 1344 32170 38640 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 38640 32170
rect 1344 32084 38640 32118
rect 35870 32002 35922 32014
rect 35870 31938 35922 31950
rect 10558 31890 10610 31902
rect 10098 31838 10110 31890
rect 10162 31838 10174 31890
rect 10558 31826 10610 31838
rect 15598 31890 15650 31902
rect 15598 31826 15650 31838
rect 17614 31890 17666 31902
rect 29262 31890 29314 31902
rect 21298 31838 21310 31890
rect 21362 31838 21374 31890
rect 23426 31838 23438 31890
rect 23490 31838 23502 31890
rect 26450 31838 26462 31890
rect 26514 31838 26526 31890
rect 28578 31838 28590 31890
rect 28642 31838 28654 31890
rect 17614 31826 17666 31838
rect 29262 31826 29314 31838
rect 35422 31890 35474 31902
rect 35422 31826 35474 31838
rect 35646 31890 35698 31902
rect 35646 31826 35698 31838
rect 15822 31778 15874 31790
rect 24670 31778 24722 31790
rect 7298 31726 7310 31778
rect 7362 31726 7374 31778
rect 24210 31726 24222 31778
rect 24274 31726 24286 31778
rect 25666 31726 25678 31778
rect 25730 31726 25742 31778
rect 15822 31714 15874 31726
rect 24670 31714 24722 31726
rect 15262 31666 15314 31678
rect 36990 31666 37042 31678
rect 7970 31614 7982 31666
rect 8034 31614 8046 31666
rect 36194 31614 36206 31666
rect 36258 31614 36270 31666
rect 15262 31602 15314 31614
rect 36990 31602 37042 31614
rect 37326 31554 37378 31566
rect 16146 31502 16158 31554
rect 16210 31502 16222 31554
rect 37326 31490 37378 31502
rect 38222 31554 38274 31566
rect 38222 31490 38274 31502
rect 1344 31386 38640 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 38640 31386
rect 1344 31300 38640 31334
rect 5742 31218 5794 31230
rect 5742 31154 5794 31166
rect 7982 31218 8034 31230
rect 7982 31154 8034 31166
rect 8990 31218 9042 31230
rect 8990 31154 9042 31166
rect 24222 31218 24274 31230
rect 24222 31154 24274 31166
rect 31950 31218 32002 31230
rect 31950 31154 32002 31166
rect 7646 31106 7698 31118
rect 7646 31042 7698 31054
rect 16270 31106 16322 31118
rect 16270 31042 16322 31054
rect 16606 31106 16658 31118
rect 16606 31042 16658 31054
rect 19966 31106 20018 31118
rect 33842 31054 33854 31106
rect 33906 31054 33918 31106
rect 19966 31042 20018 31054
rect 9886 30994 9938 31006
rect 2482 30942 2494 30994
rect 2546 30942 2558 30994
rect 9886 30930 9938 30942
rect 10110 30994 10162 31006
rect 10110 30930 10162 30942
rect 19854 30994 19906 31006
rect 33170 30942 33182 30994
rect 33234 30942 33246 30994
rect 19854 30930 19906 30942
rect 19070 30882 19122 30894
rect 3154 30830 3166 30882
rect 3218 30830 3230 30882
rect 5282 30830 5294 30882
rect 5346 30830 5358 30882
rect 19070 30818 19122 30830
rect 19518 30882 19570 30894
rect 19518 30818 19570 30830
rect 22878 30882 22930 30894
rect 22878 30818 22930 30830
rect 23214 30882 23266 30894
rect 23214 30818 23266 30830
rect 30494 30882 30546 30894
rect 30494 30818 30546 30830
rect 31278 30882 31330 30894
rect 31278 30818 31330 30830
rect 32398 30882 32450 30894
rect 36430 30882 36482 30894
rect 35970 30830 35982 30882
rect 36034 30830 36046 30882
rect 32398 30818 32450 30830
rect 36430 30818 36482 30830
rect 19966 30770 20018 30782
rect 10434 30718 10446 30770
rect 10498 30718 10510 30770
rect 19966 30706 20018 30718
rect 23438 30770 23490 30782
rect 23438 30706 23490 30718
rect 23774 30770 23826 30782
rect 23774 30706 23826 30718
rect 1344 30602 38640 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 38640 30602
rect 1344 30516 38640 30550
rect 19406 30434 19458 30446
rect 19406 30370 19458 30382
rect 31838 30434 31890 30446
rect 31838 30370 31890 30382
rect 19182 30322 19234 30334
rect 16706 30270 16718 30322
rect 16770 30270 16782 30322
rect 18834 30270 18846 30322
rect 18898 30270 18910 30322
rect 19182 30258 19234 30270
rect 4734 30210 4786 30222
rect 4734 30146 4786 30158
rect 10670 30210 10722 30222
rect 22206 30210 22258 30222
rect 12674 30158 12686 30210
rect 12738 30158 12750 30210
rect 15922 30158 15934 30210
rect 15986 30158 15998 30210
rect 10670 30146 10722 30158
rect 22206 30146 22258 30158
rect 22430 30210 22482 30222
rect 22430 30146 22482 30158
rect 24110 30210 24162 30222
rect 24110 30146 24162 30158
rect 26910 30210 26962 30222
rect 26910 30146 26962 30158
rect 31614 30210 31666 30222
rect 32162 30158 32174 30210
rect 32226 30158 32238 30210
rect 32722 30158 32734 30210
rect 32786 30158 32798 30210
rect 31614 30146 31666 30158
rect 3502 30098 3554 30110
rect 3502 30034 3554 30046
rect 3838 30098 3890 30110
rect 3838 30034 3890 30046
rect 20078 30098 20130 30110
rect 20078 30034 20130 30046
rect 29822 30098 29874 30110
rect 29822 30034 29874 30046
rect 30494 30098 30546 30110
rect 30494 30034 30546 30046
rect 30830 30098 30882 30110
rect 30830 30034 30882 30046
rect 32510 30098 32562 30110
rect 32510 30034 32562 30046
rect 32958 30098 33010 30110
rect 32958 30034 33010 30046
rect 11006 29986 11058 29998
rect 11006 29922 11058 29934
rect 12910 29986 12962 29998
rect 20414 29986 20466 29998
rect 23214 29986 23266 29998
rect 19730 29934 19742 29986
rect 19794 29934 19806 29986
rect 22754 29934 22766 29986
rect 22818 29934 22830 29986
rect 12910 29922 12962 29934
rect 20414 29922 20466 29934
rect 23214 29922 23266 29934
rect 24446 29986 24498 29998
rect 24446 29922 24498 29934
rect 30158 29986 30210 29998
rect 30158 29922 30210 29934
rect 31054 29986 31106 29998
rect 31054 29922 31106 29934
rect 31278 29986 31330 29998
rect 31278 29922 31330 29934
rect 31390 29986 31442 29998
rect 31390 29922 31442 29934
rect 33070 29986 33122 29998
rect 33070 29922 33122 29934
rect 1344 29818 38640 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 38640 29818
rect 1344 29732 38640 29766
rect 9886 29650 9938 29662
rect 16606 29650 16658 29662
rect 4946 29598 4958 29650
rect 5010 29598 5022 29650
rect 15698 29598 15710 29650
rect 15762 29598 15774 29650
rect 9886 29586 9938 29598
rect 16606 29586 16658 29598
rect 17502 29650 17554 29662
rect 17502 29586 17554 29598
rect 23438 29650 23490 29662
rect 23438 29586 23490 29598
rect 25902 29650 25954 29662
rect 25902 29586 25954 29598
rect 27246 29650 27298 29662
rect 28130 29598 28142 29650
rect 28194 29598 28206 29650
rect 33618 29598 33630 29650
rect 33682 29598 33694 29650
rect 27246 29586 27298 29598
rect 10782 29538 10834 29550
rect 22430 29538 22482 29550
rect 13458 29486 13470 29538
rect 13522 29486 13534 29538
rect 15474 29486 15486 29538
rect 15538 29486 15550 29538
rect 20514 29486 20526 29538
rect 20578 29486 20590 29538
rect 10782 29474 10834 29486
rect 22430 29474 22482 29486
rect 22766 29538 22818 29550
rect 30370 29486 30382 29538
rect 30434 29486 30446 29538
rect 37426 29486 37438 29538
rect 37490 29486 37502 29538
rect 22766 29474 22818 29486
rect 5518 29426 5570 29438
rect 1698 29374 1710 29426
rect 1762 29374 1774 29426
rect 5518 29362 5570 29374
rect 10558 29426 10610 29438
rect 14702 29426 14754 29438
rect 21758 29426 21810 29438
rect 14130 29374 14142 29426
rect 14194 29374 14206 29426
rect 15810 29374 15822 29426
rect 15874 29374 15886 29426
rect 16258 29374 16270 29426
rect 16322 29374 16334 29426
rect 21186 29374 21198 29426
rect 21250 29374 21262 29426
rect 10558 29362 10610 29374
rect 14702 29362 14754 29374
rect 21758 29362 21810 29374
rect 24110 29426 24162 29438
rect 24110 29362 24162 29374
rect 24334 29426 24386 29438
rect 24334 29362 24386 29374
rect 26686 29426 26738 29438
rect 33070 29426 33122 29438
rect 27010 29374 27022 29426
rect 27074 29374 27086 29426
rect 29698 29374 29710 29426
rect 29762 29374 29774 29426
rect 38210 29374 38222 29426
rect 38274 29374 38286 29426
rect 26686 29362 26738 29374
rect 33070 29362 33122 29374
rect 7086 29314 7138 29326
rect 26238 29314 26290 29326
rect 2482 29262 2494 29314
rect 2546 29262 2558 29314
rect 4610 29262 4622 29314
rect 4674 29262 4686 29314
rect 11330 29262 11342 29314
rect 11394 29262 11406 29314
rect 18386 29262 18398 29314
rect 18450 29262 18462 29314
rect 7086 29250 7138 29262
rect 26238 29250 26290 29262
rect 27358 29314 27410 29326
rect 27358 29250 27410 29262
rect 27582 29314 27634 29326
rect 32498 29262 32510 29314
rect 32562 29262 32574 29314
rect 35298 29262 35310 29314
rect 35362 29262 35374 29314
rect 27582 29250 27634 29262
rect 5294 29202 5346 29214
rect 5294 29138 5346 29150
rect 10222 29202 10274 29214
rect 27806 29202 27858 29214
rect 23762 29150 23774 29202
rect 23826 29150 23838 29202
rect 10222 29138 10274 29150
rect 27806 29138 27858 29150
rect 33294 29202 33346 29214
rect 33294 29138 33346 29150
rect 1344 29034 38640 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 38640 29034
rect 1344 28948 38640 28982
rect 13470 28866 13522 28878
rect 13470 28802 13522 28814
rect 13806 28866 13858 28878
rect 13806 28802 13858 28814
rect 19182 28866 19234 28878
rect 19182 28802 19234 28814
rect 20302 28866 20354 28878
rect 20302 28802 20354 28814
rect 27470 28866 27522 28878
rect 30718 28866 30770 28878
rect 30370 28814 30382 28866
rect 30434 28814 30446 28866
rect 32386 28814 32398 28866
rect 32450 28814 32462 28866
rect 27470 28802 27522 28814
rect 30718 28802 30770 28814
rect 4398 28754 4450 28766
rect 4398 28690 4450 28702
rect 4846 28754 4898 28766
rect 4846 28690 4898 28702
rect 6526 28754 6578 28766
rect 6526 28690 6578 28702
rect 7310 28754 7362 28766
rect 7310 28690 7362 28702
rect 9214 28754 9266 28766
rect 14030 28754 14082 28766
rect 10770 28702 10782 28754
rect 10834 28702 10846 28754
rect 12898 28702 12910 28754
rect 12962 28702 12974 28754
rect 9214 28690 9266 28702
rect 14030 28690 14082 28702
rect 17054 28754 17106 28766
rect 27246 28754 27298 28766
rect 24770 28702 24782 28754
rect 24834 28702 24846 28754
rect 26898 28702 26910 28754
rect 26962 28702 26974 28754
rect 17054 28690 17106 28702
rect 27246 28690 27298 28702
rect 30046 28754 30098 28766
rect 30046 28690 30098 28702
rect 30942 28754 30994 28766
rect 30942 28690 30994 28702
rect 31838 28754 31890 28766
rect 31838 28690 31890 28702
rect 32846 28754 32898 28766
rect 32846 28690 32898 28702
rect 3390 28642 3442 28654
rect 4174 28642 4226 28654
rect 3826 28590 3838 28642
rect 3890 28590 3902 28642
rect 3390 28578 3442 28590
rect 4174 28578 4226 28590
rect 6302 28642 6354 28654
rect 6302 28578 6354 28590
rect 6750 28642 6802 28654
rect 29262 28642 29314 28654
rect 8194 28590 8206 28642
rect 8258 28590 8270 28642
rect 10098 28590 10110 28642
rect 10162 28590 10174 28642
rect 18610 28590 18622 28642
rect 18674 28590 18686 28642
rect 23986 28590 23998 28642
rect 24050 28590 24062 28642
rect 27794 28590 27806 28642
rect 27858 28590 27870 28642
rect 28354 28590 28366 28642
rect 28418 28590 28430 28642
rect 6750 28578 6802 28590
rect 29262 28578 29314 28590
rect 32062 28642 32114 28654
rect 32062 28578 32114 28590
rect 3054 28530 3106 28542
rect 3054 28466 3106 28478
rect 6414 28530 6466 28542
rect 6414 28466 6466 28478
rect 6638 28530 6690 28542
rect 6638 28466 6690 28478
rect 7982 28530 8034 28542
rect 7982 28466 8034 28478
rect 20190 28530 20242 28542
rect 20190 28466 20242 28478
rect 20302 28418 20354 28430
rect 20302 28354 20354 28366
rect 28142 28418 28194 28430
rect 28142 28354 28194 28366
rect 38222 28418 38274 28430
rect 38222 28354 38274 28366
rect 1344 28250 38640 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 38640 28250
rect 1344 28164 38640 28198
rect 13246 28082 13298 28094
rect 13246 28018 13298 28030
rect 13582 28082 13634 28094
rect 13582 28018 13634 28030
rect 17614 28082 17666 28094
rect 17614 28018 17666 28030
rect 17838 28082 17890 28094
rect 17838 28018 17890 28030
rect 17950 28082 18002 28094
rect 17950 28018 18002 28030
rect 18510 28082 18562 28094
rect 18510 28018 18562 28030
rect 20526 28082 20578 28094
rect 20526 28018 20578 28030
rect 25342 28082 25394 28094
rect 25342 28018 25394 28030
rect 26798 28082 26850 28094
rect 26798 28018 26850 28030
rect 30718 28082 30770 28094
rect 30718 28018 30770 28030
rect 32622 28082 32674 28094
rect 32622 28018 32674 28030
rect 36878 28082 36930 28094
rect 36878 28018 36930 28030
rect 16830 27970 16882 27982
rect 8194 27918 8206 27970
rect 8258 27918 8270 27970
rect 16830 27906 16882 27918
rect 17726 27970 17778 27982
rect 25566 27970 25618 27982
rect 32062 27970 32114 27982
rect 22306 27918 22318 27970
rect 22370 27918 22382 27970
rect 28130 27918 28142 27970
rect 28194 27918 28206 27970
rect 17726 27906 17778 27918
rect 25566 27906 25618 27918
rect 32062 27906 32114 27918
rect 32510 27970 32562 27982
rect 32510 27906 32562 27918
rect 9886 27858 9938 27870
rect 8978 27806 8990 27858
rect 9042 27806 9054 27858
rect 9886 27794 9938 27806
rect 10558 27858 10610 27870
rect 20078 27858 20130 27870
rect 25678 27858 25730 27870
rect 36990 27858 37042 27870
rect 16594 27806 16606 27858
rect 16658 27806 16670 27858
rect 17378 27806 17390 27858
rect 17442 27806 17454 27858
rect 21634 27806 21646 27858
rect 21698 27806 21710 27858
rect 26338 27806 26350 27858
rect 26402 27806 26414 27858
rect 26562 27806 26574 27858
rect 26626 27806 26638 27858
rect 27458 27806 27470 27858
rect 27522 27806 27534 27858
rect 32274 27806 32286 27858
rect 32338 27806 32350 27858
rect 10558 27794 10610 27806
rect 20078 27794 20130 27806
rect 25678 27794 25730 27806
rect 36990 27794 37042 27806
rect 4622 27746 4674 27758
rect 10110 27746 10162 27758
rect 31502 27746 31554 27758
rect 6066 27694 6078 27746
rect 6130 27694 6142 27746
rect 24434 27694 24446 27746
rect 24498 27694 24510 27746
rect 26674 27694 26686 27746
rect 26738 27694 26750 27746
rect 30258 27694 30270 27746
rect 30322 27694 30334 27746
rect 4622 27682 4674 27694
rect 10110 27682 10162 27694
rect 31502 27682 31554 27694
rect 9550 27634 9602 27646
rect 30482 27582 30494 27634
rect 30546 27631 30558 27634
rect 30818 27631 30830 27634
rect 30546 27585 30830 27631
rect 30546 27582 30558 27585
rect 30818 27582 30830 27585
rect 30882 27582 30894 27634
rect 9550 27570 9602 27582
rect 1344 27466 38640 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 38640 27466
rect 1344 27380 38640 27414
rect 31502 27298 31554 27310
rect 5506 27246 5518 27298
rect 5570 27295 5582 27298
rect 6066 27295 6078 27298
rect 5570 27249 6078 27295
rect 5570 27246 5582 27249
rect 6066 27246 6078 27249
rect 6130 27246 6142 27298
rect 29922 27246 29934 27298
rect 29986 27295 29998 27298
rect 30706 27295 30718 27298
rect 29986 27249 30718 27295
rect 29986 27246 29998 27249
rect 30706 27246 30718 27249
rect 30770 27246 30782 27298
rect 31502 27234 31554 27246
rect 5742 27186 5794 27198
rect 24670 27186 24722 27198
rect 4722 27134 4734 27186
rect 4786 27134 4798 27186
rect 6290 27134 6302 27186
rect 6354 27134 6366 27186
rect 13458 27134 13470 27186
rect 13522 27134 13534 27186
rect 17714 27134 17726 27186
rect 17778 27134 17790 27186
rect 19842 27134 19854 27186
rect 19906 27134 19918 27186
rect 5742 27122 5794 27134
rect 24670 27122 24722 27134
rect 26910 27186 26962 27198
rect 26910 27122 26962 27134
rect 29934 27186 29986 27198
rect 29934 27122 29986 27134
rect 31838 27186 31890 27198
rect 36206 27186 36258 27198
rect 32386 27134 32398 27186
rect 32450 27134 32462 27186
rect 31838 27122 31890 27134
rect 36206 27122 36258 27134
rect 9662 27074 9714 27086
rect 20302 27074 20354 27086
rect 30830 27074 30882 27086
rect 1810 27022 1822 27074
rect 1874 27022 1886 27074
rect 9090 27022 9102 27074
rect 9154 27022 9166 27074
rect 16258 27022 16270 27074
rect 16322 27022 16334 27074
rect 16930 27022 16942 27074
rect 16994 27022 17006 27074
rect 26450 27022 26462 27074
rect 26514 27022 26526 27074
rect 9662 27010 9714 27022
rect 20302 27010 20354 27022
rect 30830 27010 30882 27022
rect 32062 27074 32114 27086
rect 32062 27010 32114 27022
rect 24222 26962 24274 26974
rect 30382 26962 30434 26974
rect 2594 26910 2606 26962
rect 2658 26910 2670 26962
rect 8418 26910 8430 26962
rect 8482 26910 8494 26962
rect 15586 26910 15598 26962
rect 15650 26910 15662 26962
rect 25890 26910 25902 26962
rect 25954 26910 25966 26962
rect 26338 26910 26350 26962
rect 26402 26910 26414 26962
rect 24222 26898 24274 26910
rect 30382 26898 30434 26910
rect 31390 26962 31442 26974
rect 31390 26898 31442 26910
rect 32622 26962 32674 26974
rect 32622 26898 32674 26910
rect 34974 26962 35026 26974
rect 36990 26962 37042 26974
rect 35186 26910 35198 26962
rect 35250 26910 35262 26962
rect 34974 26898 35026 26910
rect 36990 26898 37042 26910
rect 38222 26962 38274 26974
rect 38222 26898 38274 26910
rect 31166 26850 31218 26862
rect 25442 26798 25454 26850
rect 25506 26798 25518 26850
rect 31166 26786 31218 26798
rect 32398 26850 32450 26862
rect 32398 26786 32450 26798
rect 37326 26850 37378 26862
rect 37326 26786 37378 26798
rect 1344 26682 38640 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 38640 26682
rect 1344 26596 38640 26630
rect 8318 26514 8370 26526
rect 8318 26450 8370 26462
rect 15038 26514 15090 26526
rect 15038 26450 15090 26462
rect 16830 26514 16882 26526
rect 23438 26514 23490 26526
rect 17378 26462 17390 26514
rect 17442 26462 17454 26514
rect 16830 26450 16882 26462
rect 23438 26450 23490 26462
rect 24334 26514 24386 26526
rect 24334 26450 24386 26462
rect 25902 26514 25954 26526
rect 25902 26450 25954 26462
rect 26014 26514 26066 26526
rect 26014 26450 26066 26462
rect 31726 26514 31778 26526
rect 31726 26450 31778 26462
rect 32062 26514 32114 26526
rect 32062 26450 32114 26462
rect 23774 26402 23826 26414
rect 22082 26350 22094 26402
rect 22146 26350 22158 26402
rect 22642 26350 22654 26402
rect 22706 26350 22718 26402
rect 37426 26350 37438 26402
rect 37490 26350 37502 26402
rect 23774 26338 23826 26350
rect 5406 26290 5458 26302
rect 17950 26290 18002 26302
rect 8082 26238 8094 26290
rect 8146 26238 8158 26290
rect 14802 26238 14814 26290
rect 14866 26238 14878 26290
rect 15810 26238 15822 26290
rect 15874 26238 15886 26290
rect 5406 26226 5458 26238
rect 17950 26226 18002 26238
rect 22878 26290 22930 26302
rect 22878 26226 22930 26238
rect 24782 26290 24834 26302
rect 25442 26238 25454 26290
rect 25506 26238 25518 26290
rect 25666 26238 25678 26290
rect 25730 26238 25742 26290
rect 38210 26238 38222 26290
rect 38274 26238 38286 26290
rect 24782 26226 24834 26238
rect 4510 26178 4562 26190
rect 4510 26114 4562 26126
rect 15486 26178 15538 26190
rect 15486 26114 15538 26126
rect 16382 26178 16434 26190
rect 16382 26114 16434 26126
rect 22990 26178 23042 26190
rect 22990 26114 23042 26126
rect 26350 26178 26402 26190
rect 35298 26126 35310 26178
rect 35362 26126 35374 26178
rect 26350 26114 26402 26126
rect 5182 26066 5234 26078
rect 4834 26014 4846 26066
rect 4898 26014 4910 26066
rect 5182 26002 5234 26014
rect 16158 26066 16210 26078
rect 16158 26002 16210 26014
rect 17726 26066 17778 26078
rect 17726 26002 17778 26014
rect 1344 25898 38640 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 38640 25898
rect 1344 25812 38640 25846
rect 25230 25730 25282 25742
rect 25230 25666 25282 25678
rect 36990 25730 37042 25742
rect 36990 25666 37042 25678
rect 6190 25618 6242 25630
rect 6190 25554 6242 25566
rect 6638 25618 6690 25630
rect 6638 25554 6690 25566
rect 17054 25618 17106 25630
rect 17054 25554 17106 25566
rect 25902 25618 25954 25630
rect 25902 25554 25954 25566
rect 26350 25618 26402 25630
rect 26350 25554 26402 25566
rect 37326 25618 37378 25630
rect 37326 25554 37378 25566
rect 5966 25506 6018 25518
rect 22082 25454 22094 25506
rect 22146 25454 22158 25506
rect 25106 25454 25118 25506
rect 25170 25454 25182 25506
rect 5966 25442 6018 25454
rect 3726 25394 3778 25406
rect 3726 25330 3778 25342
rect 4062 25394 4114 25406
rect 4062 25330 4114 25342
rect 12686 25394 12738 25406
rect 26126 25394 26178 25406
rect 23538 25342 23550 25394
rect 23602 25342 23614 25394
rect 24434 25342 24446 25394
rect 24498 25342 24510 25394
rect 12686 25330 12738 25342
rect 26126 25330 26178 25342
rect 27022 25394 27074 25406
rect 27022 25330 27074 25342
rect 35422 25394 35474 25406
rect 35422 25330 35474 25342
rect 36094 25394 36146 25406
rect 36094 25330 36146 25342
rect 37550 25394 37602 25406
rect 37550 25330 37602 25342
rect 37886 25394 37938 25406
rect 37886 25330 37938 25342
rect 38222 25394 38274 25406
rect 38222 25330 38274 25342
rect 27358 25282 27410 25294
rect 5618 25230 5630 25282
rect 5682 25230 5694 25282
rect 26674 25230 26686 25282
rect 26738 25230 26750 25282
rect 27358 25218 27410 25230
rect 27806 25282 27858 25294
rect 27806 25218 27858 25230
rect 30158 25282 30210 25294
rect 30158 25218 30210 25230
rect 31054 25282 31106 25294
rect 31054 25218 31106 25230
rect 31502 25282 31554 25294
rect 31502 25218 31554 25230
rect 35758 25282 35810 25294
rect 35758 25218 35810 25230
rect 1344 25114 38640 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 38640 25114
rect 1344 25028 38640 25062
rect 14030 24946 14082 24958
rect 14030 24882 14082 24894
rect 24670 24946 24722 24958
rect 24670 24882 24722 24894
rect 25678 24946 25730 24958
rect 25678 24882 25730 24894
rect 31166 24946 31218 24958
rect 31166 24882 31218 24894
rect 3278 24834 3330 24846
rect 3278 24770 3330 24782
rect 3614 24834 3666 24846
rect 3614 24770 3666 24782
rect 3950 24834 4002 24846
rect 3950 24770 4002 24782
rect 4286 24834 4338 24846
rect 30270 24834 30322 24846
rect 27794 24782 27806 24834
rect 27858 24782 27870 24834
rect 4286 24770 4338 24782
rect 30270 24770 30322 24782
rect 31838 24834 31890 24846
rect 31838 24770 31890 24782
rect 33406 24834 33458 24846
rect 35746 24782 35758 24834
rect 35810 24782 35822 24834
rect 33406 24770 33458 24782
rect 13022 24722 13074 24734
rect 32062 24722 32114 24734
rect 9650 24670 9662 24722
rect 9714 24670 9726 24722
rect 21410 24670 21422 24722
rect 21474 24670 21486 24722
rect 27010 24670 27022 24722
rect 27074 24670 27086 24722
rect 31378 24670 31390 24722
rect 31442 24670 31454 24722
rect 13022 24658 13074 24670
rect 32062 24658 32114 24670
rect 33070 24722 33122 24734
rect 34962 24670 34974 24722
rect 35026 24670 35038 24722
rect 33070 24658 33122 24670
rect 30830 24610 30882 24622
rect 10322 24558 10334 24610
rect 10386 24558 10398 24610
rect 12450 24558 12462 24610
rect 12514 24558 12526 24610
rect 22082 24558 22094 24610
rect 22146 24558 22158 24610
rect 24210 24558 24222 24610
rect 24274 24558 24286 24610
rect 29922 24558 29934 24610
rect 29986 24558 29998 24610
rect 30830 24546 30882 24558
rect 32398 24610 32450 24622
rect 32398 24546 32450 24558
rect 34638 24610 34690 24622
rect 37874 24558 37886 24610
rect 37938 24558 37950 24610
rect 34638 24546 34690 24558
rect 13246 24498 13298 24510
rect 30494 24498 30546 24510
rect 13570 24446 13582 24498
rect 13634 24446 13646 24498
rect 13246 24434 13298 24446
rect 30494 24434 30546 24446
rect 1344 24330 38640 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 38640 24330
rect 1344 24244 38640 24278
rect 12798 24162 12850 24174
rect 5618 24110 5630 24162
rect 5682 24110 5694 24162
rect 12798 24098 12850 24110
rect 19630 24162 19682 24174
rect 19630 24098 19682 24110
rect 26126 24050 26178 24062
rect 38334 24050 38386 24062
rect 16930 23998 16942 24050
rect 16994 23998 17006 24050
rect 32610 23998 32622 24050
rect 32674 23998 32686 24050
rect 32946 23998 32958 24050
rect 33010 23998 33022 24050
rect 35074 23998 35086 24050
rect 35138 23998 35150 24050
rect 26126 23986 26178 23998
rect 38334 23986 38386 23998
rect 5966 23938 6018 23950
rect 5966 23874 6018 23886
rect 6190 23938 6242 23950
rect 13582 23938 13634 23950
rect 18510 23938 18562 23950
rect 25902 23938 25954 23950
rect 9762 23886 9774 23938
rect 9826 23886 9838 23938
rect 16258 23886 16270 23938
rect 16322 23886 16334 23938
rect 21858 23886 21870 23938
rect 21922 23886 21934 23938
rect 25554 23886 25566 23938
rect 25618 23886 25630 23938
rect 29698 23886 29710 23938
rect 29762 23886 29774 23938
rect 35746 23886 35758 23938
rect 35810 23886 35822 23938
rect 6190 23874 6242 23886
rect 13582 23874 13634 23886
rect 18510 23874 18562 23886
rect 25902 23874 25954 23886
rect 9998 23826 10050 23838
rect 9998 23762 10050 23774
rect 12686 23826 12738 23838
rect 18286 23826 18338 23838
rect 16370 23774 16382 23826
rect 16434 23774 16446 23826
rect 12686 23762 12738 23774
rect 18286 23762 18338 23774
rect 19518 23826 19570 23838
rect 19518 23762 19570 23774
rect 20414 23826 20466 23838
rect 20414 23762 20466 23774
rect 20750 23826 20802 23838
rect 20750 23762 20802 23774
rect 25230 23826 25282 23838
rect 25230 23762 25282 23774
rect 27918 23826 27970 23838
rect 30482 23774 30494 23826
rect 30546 23774 30558 23826
rect 27918 23762 27970 23774
rect 5070 23714 5122 23726
rect 5070 23650 5122 23662
rect 9214 23714 9266 23726
rect 9214 23650 9266 23662
rect 12350 23714 12402 23726
rect 12350 23650 12402 23662
rect 12798 23714 12850 23726
rect 12798 23650 12850 23662
rect 13918 23714 13970 23726
rect 19630 23714 19682 23726
rect 18834 23662 18846 23714
rect 18898 23662 18910 23714
rect 13918 23650 13970 23662
rect 19630 23650 19682 23662
rect 22094 23714 22146 23726
rect 22094 23650 22146 23662
rect 27582 23714 27634 23726
rect 27582 23650 27634 23662
rect 1344 23546 38640 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 38640 23546
rect 1344 23460 38640 23494
rect 5518 23378 5570 23390
rect 5518 23314 5570 23326
rect 6750 23378 6802 23390
rect 6750 23314 6802 23326
rect 8654 23378 8706 23390
rect 10558 23378 10610 23390
rect 10098 23326 10110 23378
rect 10162 23326 10174 23378
rect 8654 23314 8706 23326
rect 10558 23314 10610 23326
rect 16718 23378 16770 23390
rect 16718 23314 16770 23326
rect 19070 23378 19122 23390
rect 19070 23314 19122 23326
rect 19966 23378 20018 23390
rect 33182 23378 33234 23390
rect 29250 23326 29262 23378
rect 29314 23326 29326 23378
rect 19966 23314 20018 23326
rect 33182 23314 33234 23326
rect 33630 23378 33682 23390
rect 33630 23314 33682 23326
rect 34750 23378 34802 23390
rect 34750 23314 34802 23326
rect 34862 23378 34914 23390
rect 36082 23326 36094 23378
rect 36146 23326 36158 23378
rect 34862 23314 34914 23326
rect 11566 23266 11618 23278
rect 24670 23266 24722 23278
rect 28590 23266 28642 23278
rect 2594 23214 2606 23266
rect 2658 23214 2670 23266
rect 14130 23214 14142 23266
rect 14194 23214 14206 23266
rect 22642 23214 22654 23266
rect 22706 23214 22718 23266
rect 27346 23214 27358 23266
rect 27410 23214 27422 23266
rect 11566 23202 11618 23214
rect 24670 23202 24722 23214
rect 28590 23202 28642 23214
rect 5294 23154 5346 23166
rect 1810 23102 1822 23154
rect 1874 23102 1886 23154
rect 5294 23090 5346 23102
rect 5406 23154 5458 23166
rect 5406 23090 5458 23102
rect 5630 23154 5682 23166
rect 6302 23154 6354 23166
rect 8542 23154 8594 23166
rect 5842 23102 5854 23154
rect 5906 23102 5918 23154
rect 8306 23102 8318 23154
rect 8370 23102 8382 23154
rect 5630 23090 5682 23102
rect 6302 23090 6354 23102
rect 8542 23090 8594 23102
rect 8766 23154 8818 23166
rect 8766 23090 8818 23102
rect 8878 23154 8930 23166
rect 8878 23090 8930 23102
rect 9774 23154 9826 23166
rect 17950 23154 18002 23166
rect 29822 23154 29874 23166
rect 34974 23154 35026 23166
rect 35534 23154 35586 23166
rect 11778 23102 11790 23154
rect 11842 23102 11854 23154
rect 13458 23102 13470 23154
rect 13522 23102 13534 23154
rect 23426 23102 23438 23154
rect 23490 23102 23502 23154
rect 24434 23102 24446 23154
rect 24498 23102 24510 23154
rect 28018 23102 28030 23154
rect 28082 23102 28094 23154
rect 34514 23102 34526 23154
rect 34578 23102 34590 23154
rect 35186 23102 35198 23154
rect 35250 23102 35262 23154
rect 9774 23090 9826 23102
rect 17950 23090 18002 23102
rect 29822 23090 29874 23102
rect 34974 23090 35026 23102
rect 35534 23090 35586 23102
rect 9550 23042 9602 23054
rect 4722 22990 4734 23042
rect 4786 22990 4798 23042
rect 9550 22978 9602 22990
rect 11006 23042 11058 23054
rect 11006 22978 11058 22990
rect 12350 23042 12402 23054
rect 17614 23042 17666 23054
rect 16258 22990 16270 23042
rect 16322 22990 16334 23042
rect 12350 22978 12402 22990
rect 17614 22978 17666 22990
rect 18174 23042 18226 23054
rect 23886 23042 23938 23054
rect 34078 23042 34130 23054
rect 20514 22990 20526 23042
rect 20578 22990 20590 23042
rect 25218 22990 25230 23042
rect 25282 22990 25294 23042
rect 18174 22978 18226 22990
rect 23886 22978 23938 22990
rect 34078 22978 34130 22990
rect 29598 22930 29650 22942
rect 35758 22930 35810 22942
rect 18498 22878 18510 22930
rect 18562 22878 18574 22930
rect 33730 22878 33742 22930
rect 33794 22927 33806 22930
rect 34290 22927 34302 22930
rect 33794 22881 34302 22927
rect 33794 22878 33806 22881
rect 34290 22878 34302 22881
rect 34354 22878 34366 22930
rect 29598 22866 29650 22878
rect 35758 22866 35810 22878
rect 1344 22762 38640 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 38640 22762
rect 1344 22676 38640 22710
rect 11778 22542 11790 22594
rect 11842 22542 11854 22594
rect 21858 22542 21870 22594
rect 21922 22542 21934 22594
rect 5070 22482 5122 22494
rect 6862 22482 6914 22494
rect 2482 22430 2494 22482
rect 2546 22430 2558 22482
rect 4610 22430 4622 22482
rect 4674 22430 4686 22482
rect 6290 22430 6302 22482
rect 6354 22430 6366 22482
rect 5070 22418 5122 22430
rect 6862 22418 6914 22430
rect 7310 22482 7362 22494
rect 12350 22482 12402 22494
rect 11442 22430 11454 22482
rect 11506 22430 11518 22482
rect 7310 22418 7362 22430
rect 12350 22418 12402 22430
rect 12798 22482 12850 22494
rect 12798 22418 12850 22430
rect 15598 22482 15650 22494
rect 21534 22482 21586 22494
rect 16370 22430 16382 22482
rect 16434 22430 16446 22482
rect 15598 22418 15650 22430
rect 21534 22418 21586 22430
rect 22206 22482 22258 22494
rect 27694 22482 27746 22494
rect 24994 22430 25006 22482
rect 25058 22430 25070 22482
rect 27122 22430 27134 22482
rect 27186 22430 27198 22482
rect 22206 22418 22258 22430
rect 27694 22418 27746 22430
rect 32734 22482 32786 22494
rect 32734 22418 32786 22430
rect 5966 22370 6018 22382
rect 12126 22370 12178 22382
rect 1810 22318 1822 22370
rect 1874 22318 1886 22370
rect 8642 22318 8654 22370
rect 8706 22318 8718 22370
rect 5966 22306 6018 22318
rect 12126 22306 12178 22318
rect 14926 22370 14978 22382
rect 19966 22370 20018 22382
rect 15250 22318 15262 22370
rect 15314 22318 15326 22370
rect 15922 22318 15934 22370
rect 15986 22318 15998 22370
rect 19170 22318 19182 22370
rect 19234 22318 19246 22370
rect 14926 22306 14978 22318
rect 19966 22306 20018 22318
rect 20414 22370 20466 22382
rect 20414 22306 20466 22318
rect 22430 22370 22482 22382
rect 24210 22318 24222 22370
rect 24274 22318 24286 22370
rect 22430 22306 22482 22318
rect 5742 22258 5794 22270
rect 19630 22258 19682 22270
rect 9314 22206 9326 22258
rect 9378 22206 9390 22258
rect 18498 22206 18510 22258
rect 18562 22206 18574 22258
rect 5742 22194 5794 22206
rect 19630 22194 19682 22206
rect 6190 22146 6242 22158
rect 6190 22082 6242 22094
rect 6302 22146 6354 22158
rect 6302 22082 6354 22094
rect 15486 22146 15538 22158
rect 15486 22082 15538 22094
rect 15710 22146 15762 22158
rect 15710 22082 15762 22094
rect 29262 22146 29314 22158
rect 29262 22082 29314 22094
rect 34190 22146 34242 22158
rect 34190 22082 34242 22094
rect 35198 22146 35250 22158
rect 35198 22082 35250 22094
rect 1344 21978 38640 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 38640 21978
rect 1344 21892 38640 21926
rect 9550 21810 9602 21822
rect 9550 21746 9602 21758
rect 15934 21810 15986 21822
rect 15934 21746 15986 21758
rect 16046 21810 16098 21822
rect 16046 21746 16098 21758
rect 16158 21810 16210 21822
rect 16158 21746 16210 21758
rect 16830 21810 16882 21822
rect 21410 21758 21422 21810
rect 21474 21758 21486 21810
rect 16830 21746 16882 21758
rect 21982 21698 22034 21710
rect 4722 21646 4734 21698
rect 4786 21646 4798 21698
rect 11554 21646 11566 21698
rect 11618 21646 11630 21698
rect 21982 21634 22034 21646
rect 5294 21586 5346 21598
rect 14142 21586 14194 21598
rect 34526 21586 34578 21598
rect 5954 21534 5966 21586
rect 6018 21534 6030 21586
rect 9762 21534 9774 21586
rect 9826 21534 9838 21586
rect 10882 21534 10894 21586
rect 10946 21534 10958 21586
rect 15698 21534 15710 21586
rect 15762 21534 15774 21586
rect 16370 21534 16382 21586
rect 16434 21534 16446 21586
rect 17378 21534 17390 21586
rect 17442 21534 17454 21586
rect 32498 21534 32510 21586
rect 32562 21534 32574 21586
rect 37762 21534 37774 21586
rect 37826 21534 37838 21586
rect 5294 21522 5346 21534
rect 14142 21522 14194 21534
rect 34526 21522 34578 21534
rect 4398 21474 4450 21486
rect 21086 21474 21138 21486
rect 33630 21474 33682 21486
rect 6738 21422 6750 21474
rect 6802 21422 6814 21474
rect 8866 21422 8878 21474
rect 8930 21422 8942 21474
rect 13682 21422 13694 21474
rect 13746 21422 13758 21474
rect 18162 21422 18174 21474
rect 18226 21422 18238 21474
rect 20290 21422 20302 21474
rect 20354 21422 20366 21474
rect 29586 21422 29598 21474
rect 29650 21422 29662 21474
rect 31714 21422 31726 21474
rect 31778 21422 31790 21474
rect 34850 21422 34862 21474
rect 34914 21422 34926 21474
rect 36978 21422 36990 21474
rect 37042 21422 37054 21474
rect 4398 21410 4450 21422
rect 21086 21410 21138 21422
rect 33630 21410 33682 21422
rect 5070 21362 5122 21374
rect 5070 21298 5122 21310
rect 21758 21362 21810 21374
rect 33406 21362 33458 21374
rect 33058 21310 33070 21362
rect 33122 21310 33134 21362
rect 21758 21298 21810 21310
rect 33406 21298 33458 21310
rect 1344 21194 38640 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 38640 21194
rect 1344 21108 38640 21142
rect 8978 20974 8990 21026
rect 9042 20974 9054 21026
rect 5742 20914 5794 20926
rect 5742 20850 5794 20862
rect 9550 20914 9602 20926
rect 9550 20850 9602 20862
rect 16382 20914 16434 20926
rect 16382 20850 16434 20862
rect 16830 20914 16882 20926
rect 18286 20914 18338 20926
rect 17714 20862 17726 20914
rect 17778 20862 17790 20914
rect 16830 20850 16882 20862
rect 18286 20850 18338 20862
rect 20526 20914 20578 20926
rect 20526 20850 20578 20862
rect 21534 20914 21586 20926
rect 21534 20850 21586 20862
rect 27022 20914 27074 20926
rect 27022 20850 27074 20862
rect 34974 20914 35026 20926
rect 34974 20850 35026 20862
rect 4174 20802 4226 20814
rect 4174 20738 4226 20750
rect 5070 20802 5122 20814
rect 5070 20738 5122 20750
rect 5966 20802 6018 20814
rect 5966 20738 6018 20750
rect 7422 20802 7474 20814
rect 7422 20738 7474 20750
rect 8430 20802 8482 20814
rect 8430 20738 8482 20750
rect 8654 20802 8706 20814
rect 27246 20802 27298 20814
rect 17378 20750 17390 20802
rect 17442 20750 17454 20802
rect 8654 20738 8706 20750
rect 27246 20738 27298 20750
rect 31838 20802 31890 20814
rect 35858 20750 35870 20802
rect 35922 20750 35934 20802
rect 31838 20738 31890 20750
rect 6638 20690 6690 20702
rect 6290 20638 6302 20690
rect 6354 20638 6366 20690
rect 6638 20626 6690 20638
rect 6974 20690 7026 20702
rect 6974 20626 7026 20638
rect 31502 20690 31554 20702
rect 31502 20626 31554 20638
rect 36094 20690 36146 20702
rect 36094 20626 36146 20638
rect 3838 20578 3890 20590
rect 3838 20514 3890 20526
rect 8094 20578 8146 20590
rect 8094 20514 8146 20526
rect 26686 20578 26738 20590
rect 32734 20578 32786 20590
rect 27570 20526 27582 20578
rect 27634 20526 27646 20578
rect 26686 20514 26738 20526
rect 32734 20514 32786 20526
rect 1344 20410 38640 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 38640 20410
rect 1344 20324 38640 20358
rect 18174 20242 18226 20254
rect 18174 20178 18226 20190
rect 20638 20130 20690 20142
rect 3266 20078 3278 20130
rect 3330 20078 3342 20130
rect 20638 20066 20690 20078
rect 20974 20130 21026 20142
rect 20974 20066 21026 20078
rect 24558 20130 24610 20142
rect 24558 20066 24610 20078
rect 27806 20130 27858 20142
rect 27806 20066 27858 20078
rect 28142 20130 28194 20142
rect 28142 20066 28194 20078
rect 34638 20130 34690 20142
rect 34638 20066 34690 20078
rect 12014 20018 12066 20030
rect 2594 19966 2606 20018
rect 2658 19966 2670 20018
rect 12014 19954 12066 19966
rect 17838 20018 17890 20030
rect 17838 19954 17890 19966
rect 23886 20018 23938 20030
rect 23886 19954 23938 19966
rect 24110 20018 24162 20030
rect 24110 19954 24162 19966
rect 34414 20018 34466 20030
rect 34414 19954 34466 19966
rect 34526 20018 34578 20030
rect 34526 19954 34578 19966
rect 34750 20018 34802 20030
rect 34962 19966 34974 20018
rect 35026 19966 35038 20018
rect 38098 19966 38110 20018
rect 38162 19966 38174 20018
rect 34750 19954 34802 19966
rect 5966 19906 6018 19918
rect 5394 19854 5406 19906
rect 5458 19854 5470 19906
rect 5966 19842 6018 19854
rect 11118 19906 11170 19918
rect 11118 19842 11170 19854
rect 23214 19906 23266 19918
rect 23214 19842 23266 19854
rect 33294 19906 33346 19918
rect 33294 19842 33346 19854
rect 33742 19906 33794 19918
rect 35298 19854 35310 19906
rect 35362 19854 35374 19906
rect 37426 19854 37438 19906
rect 37490 19854 37502 19906
rect 33742 19842 33794 19854
rect 11790 19794 11842 19806
rect 11442 19742 11454 19794
rect 11506 19742 11518 19794
rect 23538 19742 23550 19794
rect 23602 19742 23614 19794
rect 11790 19730 11842 19742
rect 1344 19626 38640 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 38640 19626
rect 1344 19540 38640 19574
rect 4174 19458 4226 19470
rect 36082 19406 36094 19458
rect 36146 19406 36158 19458
rect 4174 19394 4226 19406
rect 4398 19346 4450 19358
rect 17278 19346 17330 19358
rect 29262 19346 29314 19358
rect 14242 19294 14254 19346
rect 14306 19294 14318 19346
rect 16370 19294 16382 19346
rect 16434 19294 16446 19346
rect 23762 19294 23774 19346
rect 23826 19294 23838 19346
rect 4398 19282 4450 19294
rect 17278 19282 17330 19294
rect 29262 19282 29314 19294
rect 29710 19346 29762 19358
rect 32398 19346 32450 19358
rect 30706 19294 30718 19346
rect 30770 19294 30782 19346
rect 29710 19282 29762 19294
rect 32398 19282 32450 19294
rect 32846 19346 32898 19358
rect 35534 19346 35586 19358
rect 33954 19294 33966 19346
rect 34018 19294 34030 19346
rect 32846 19282 32898 19294
rect 35534 19282 35586 19294
rect 16830 19234 16882 19246
rect 30382 19234 30434 19246
rect 13458 19182 13470 19234
rect 13522 19182 13534 19234
rect 17154 19182 17166 19234
rect 17218 19182 17230 19234
rect 23202 19182 23214 19234
rect 23266 19182 23278 19234
rect 26674 19182 26686 19234
rect 26738 19182 26750 19234
rect 16830 19170 16882 19182
rect 4846 19010 4898 19022
rect 17169 19010 17215 19182
rect 30382 19170 30434 19182
rect 30494 19234 30546 19246
rect 30494 19170 30546 19182
rect 30830 19234 30882 19246
rect 30830 19170 30882 19182
rect 33630 19234 33682 19246
rect 34862 19234 34914 19246
rect 34066 19182 34078 19234
rect 34130 19182 34142 19234
rect 33630 19170 33682 19182
rect 34862 19170 34914 19182
rect 35758 19234 35810 19246
rect 35758 19170 35810 19182
rect 33406 19122 33458 19134
rect 25890 19070 25902 19122
rect 25954 19070 25966 19122
rect 33406 19058 33458 19070
rect 34638 19122 34690 19134
rect 34638 19058 34690 19070
rect 36990 19122 37042 19134
rect 36990 19058 37042 19070
rect 37326 19122 37378 19134
rect 37326 19058 37378 19070
rect 23438 19010 23490 19022
rect 3826 18958 3838 19010
rect 3890 18958 3902 19010
rect 17154 18958 17166 19010
rect 17218 18958 17230 19010
rect 4846 18946 4898 18958
rect 23438 18946 23490 18958
rect 27134 19010 27186 19022
rect 27134 18946 27186 18958
rect 30718 19010 30770 19022
rect 30718 18946 30770 18958
rect 31390 19010 31442 19022
rect 31390 18946 31442 18958
rect 33854 19010 33906 19022
rect 35186 18958 35198 19010
rect 35250 18958 35262 19010
rect 33854 18946 33906 18958
rect 1344 18842 38640 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 38640 18842
rect 1344 18756 38640 18790
rect 34302 18674 34354 18686
rect 17714 18622 17726 18674
rect 17778 18622 17790 18674
rect 34302 18610 34354 18622
rect 9550 18562 9602 18574
rect 9550 18498 9602 18510
rect 10334 18562 10386 18574
rect 10334 18498 10386 18510
rect 10670 18562 10722 18574
rect 10670 18498 10722 18510
rect 19854 18562 19906 18574
rect 19854 18498 19906 18510
rect 19966 18562 20018 18574
rect 31726 18562 31778 18574
rect 28354 18510 28366 18562
rect 28418 18510 28430 18562
rect 19966 18498 20018 18510
rect 31726 18498 31778 18510
rect 33742 18562 33794 18574
rect 33742 18498 33794 18510
rect 9886 18450 9938 18462
rect 2258 18398 2270 18450
rect 2322 18398 2334 18450
rect 9886 18386 9938 18398
rect 16830 18450 16882 18462
rect 16830 18386 16882 18398
rect 20414 18450 20466 18462
rect 31054 18450 31106 18462
rect 27682 18398 27694 18450
rect 27746 18398 27758 18450
rect 20414 18386 20466 18398
rect 31054 18386 31106 18398
rect 32062 18450 32114 18462
rect 33506 18398 33518 18450
rect 33570 18398 33582 18450
rect 38098 18398 38110 18450
rect 38162 18398 38174 18450
rect 32062 18386 32114 18398
rect 5518 18338 5570 18350
rect 2930 18286 2942 18338
rect 2994 18286 3006 18338
rect 5058 18286 5070 18338
rect 5122 18286 5134 18338
rect 5518 18274 5570 18286
rect 18286 18338 18338 18350
rect 18286 18274 18338 18286
rect 20974 18338 21026 18350
rect 30830 18338 30882 18350
rect 30482 18286 30494 18338
rect 30546 18286 30558 18338
rect 20974 18274 21026 18286
rect 30830 18274 30882 18286
rect 31390 18338 31442 18350
rect 31390 18274 31442 18286
rect 32510 18338 32562 18350
rect 32510 18274 32562 18286
rect 34974 18338 35026 18350
rect 35298 18286 35310 18338
rect 35362 18286 35374 18338
rect 37426 18286 37438 18338
rect 37490 18286 37502 18338
rect 34974 18274 35026 18286
rect 18062 18226 18114 18238
rect 5282 18174 5294 18226
rect 5346 18223 5358 18226
rect 5618 18223 5630 18226
rect 5346 18177 5630 18223
rect 5346 18174 5358 18177
rect 5618 18174 5630 18177
rect 5682 18174 5694 18226
rect 18062 18162 18114 18174
rect 19854 18226 19906 18238
rect 19854 18162 19906 18174
rect 1344 18058 38640 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 38640 18058
rect 1344 17972 38640 18006
rect 5854 17890 5906 17902
rect 33618 17838 33630 17890
rect 33682 17838 33694 17890
rect 5854 17826 5906 17838
rect 5070 17778 5122 17790
rect 5070 17714 5122 17726
rect 5630 17778 5682 17790
rect 30046 17778 30098 17790
rect 34190 17778 34242 17790
rect 7970 17726 7982 17778
rect 8034 17726 8046 17778
rect 10098 17726 10110 17778
rect 10162 17726 10174 17778
rect 17826 17726 17838 17778
rect 17890 17726 17902 17778
rect 19954 17726 19966 17778
rect 20018 17726 20030 17778
rect 23426 17726 23438 17778
rect 23490 17726 23502 17778
rect 25554 17726 25566 17778
rect 25618 17726 25630 17778
rect 31154 17726 31166 17778
rect 31218 17726 31230 17778
rect 33282 17726 33294 17778
rect 33346 17726 33358 17778
rect 5630 17714 5682 17726
rect 30046 17714 30098 17726
rect 34190 17714 34242 17726
rect 3614 17666 3666 17678
rect 33966 17666 34018 17678
rect 6178 17614 6190 17666
rect 6242 17614 6254 17666
rect 6738 17614 6750 17666
rect 6802 17614 6814 17666
rect 10770 17614 10782 17666
rect 10834 17614 10846 17666
rect 13682 17614 13694 17666
rect 13746 17614 13758 17666
rect 20738 17614 20750 17666
rect 20802 17614 20814 17666
rect 22642 17614 22654 17666
rect 22706 17614 22718 17666
rect 26114 17614 26126 17666
rect 26178 17614 26190 17666
rect 30482 17614 30494 17666
rect 30546 17614 30558 17666
rect 3614 17602 3666 17614
rect 33966 17602 34018 17614
rect 35086 17666 35138 17678
rect 35086 17602 35138 17614
rect 3278 17554 3330 17566
rect 3278 17490 3330 17502
rect 14478 17554 14530 17566
rect 14478 17490 14530 17502
rect 21310 17554 21362 17566
rect 21310 17490 21362 17502
rect 25902 17554 25954 17566
rect 25902 17490 25954 17502
rect 34638 17554 34690 17566
rect 34638 17490 34690 17502
rect 6526 17442 6578 17454
rect 6526 17378 6578 17390
rect 11342 17442 11394 17454
rect 11342 17378 11394 17390
rect 13470 17442 13522 17454
rect 13470 17378 13522 17390
rect 14142 17442 14194 17454
rect 14142 17378 14194 17390
rect 14926 17442 14978 17454
rect 14926 17378 14978 17390
rect 21646 17442 21698 17454
rect 21646 17378 21698 17390
rect 26686 17442 26738 17454
rect 26686 17378 26738 17390
rect 1344 17274 38640 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 38640 17274
rect 1344 17188 38640 17222
rect 8654 17106 8706 17118
rect 16270 17106 16322 17118
rect 15026 17054 15038 17106
rect 15090 17054 15102 17106
rect 8654 17042 8706 17054
rect 16270 17042 16322 17054
rect 17502 17106 17554 17118
rect 26910 17106 26962 17118
rect 25890 17054 25902 17106
rect 25954 17054 25966 17106
rect 17502 17042 17554 17054
rect 26910 17042 26962 17054
rect 29262 17106 29314 17118
rect 29262 17042 29314 17054
rect 32510 17106 32562 17118
rect 32510 17042 32562 17054
rect 36654 17106 36706 17118
rect 36654 17042 36706 17054
rect 17950 16994 18002 17006
rect 23102 16994 23154 17006
rect 6066 16942 6078 16994
rect 6130 16942 6142 16994
rect 12562 16942 12574 16994
rect 12626 16942 12638 16994
rect 21858 16942 21870 16994
rect 21922 16942 21934 16994
rect 33842 16942 33854 16994
rect 33906 16942 33918 16994
rect 17950 16930 18002 16942
rect 23102 16930 23154 16942
rect 15598 16882 15650 16894
rect 5394 16830 5406 16882
rect 5458 16830 5470 16882
rect 11778 16830 11790 16882
rect 11842 16830 11854 16882
rect 15598 16818 15650 16830
rect 16158 16882 16210 16894
rect 16158 16818 16210 16830
rect 16494 16882 16546 16894
rect 26238 16882 26290 16894
rect 36318 16882 36370 16894
rect 16706 16830 16718 16882
rect 16770 16830 16782 16882
rect 22642 16830 22654 16882
rect 22706 16830 22718 16882
rect 33170 16830 33182 16882
rect 33234 16830 33246 16882
rect 16494 16818 16546 16830
rect 26238 16818 26290 16830
rect 36318 16818 36370 16830
rect 16382 16770 16434 16782
rect 8194 16718 8206 16770
rect 8258 16718 8270 16770
rect 14690 16718 14702 16770
rect 14754 16718 14766 16770
rect 16382 16706 16434 16718
rect 19070 16770 19122 16782
rect 26462 16770 26514 16782
rect 19730 16718 19742 16770
rect 19794 16718 19806 16770
rect 19070 16706 19122 16718
rect 26462 16706 26514 16718
rect 28814 16770 28866 16782
rect 35970 16718 35982 16770
rect 36034 16718 36046 16770
rect 28814 16706 28866 16718
rect 15374 16658 15426 16670
rect 28802 16606 28814 16658
rect 28866 16655 28878 16658
rect 29362 16655 29374 16658
rect 28866 16609 29374 16655
rect 28866 16606 28878 16609
rect 29362 16606 29374 16609
rect 29426 16606 29438 16658
rect 15374 16594 15426 16606
rect 1344 16490 38640 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 38640 16490
rect 1344 16404 38640 16438
rect 22094 16322 22146 16334
rect 13458 16270 13470 16322
rect 13522 16270 13534 16322
rect 22094 16258 22146 16270
rect 29486 16322 29538 16334
rect 35522 16270 35534 16322
rect 35586 16270 35598 16322
rect 29486 16258 29538 16270
rect 12910 16210 12962 16222
rect 9314 16158 9326 16210
rect 9378 16158 9390 16210
rect 11442 16158 11454 16210
rect 11506 16158 11518 16210
rect 12910 16146 12962 16158
rect 13806 16210 13858 16222
rect 21870 16210 21922 16222
rect 15922 16158 15934 16210
rect 15986 16158 15998 16210
rect 13806 16146 13858 16158
rect 21870 16146 21922 16158
rect 22878 16210 22930 16222
rect 22878 16146 22930 16158
rect 23438 16210 23490 16222
rect 34974 16210 35026 16222
rect 25666 16158 25678 16210
rect 25730 16158 25742 16210
rect 23438 16146 23490 16158
rect 34974 16146 35026 16158
rect 12014 16098 12066 16110
rect 14030 16098 14082 16110
rect 8642 16046 8654 16098
rect 8706 16046 8718 16098
rect 12450 16046 12462 16098
rect 12514 16046 12526 16098
rect 12014 16034 12066 16046
rect 14030 16034 14082 16046
rect 14478 16098 14530 16110
rect 21422 16098 21474 16110
rect 29710 16098 29762 16110
rect 18722 16046 18734 16098
rect 18786 16046 18798 16098
rect 19282 16046 19294 16098
rect 19346 16046 19358 16098
rect 20738 16046 20750 16098
rect 20802 16046 20814 16098
rect 28578 16046 28590 16098
rect 28642 16046 28654 16098
rect 14478 16034 14530 16046
rect 21422 16034 21474 16046
rect 29710 16034 29762 16046
rect 35198 16098 35250 16110
rect 35198 16034 35250 16046
rect 11790 15986 11842 15998
rect 20526 15986 20578 15998
rect 18050 15934 18062 15986
rect 18114 15934 18126 15986
rect 19394 15934 19406 15986
rect 19458 15934 19470 15986
rect 27794 15934 27806 15986
rect 27858 15934 27870 15986
rect 11790 15922 11842 15934
rect 20526 15922 20578 15934
rect 12126 15874 12178 15886
rect 12126 15810 12178 15822
rect 12238 15874 12290 15886
rect 12238 15810 12290 15822
rect 14926 15874 14978 15886
rect 34638 15874 34690 15886
rect 20402 15822 20414 15874
rect 20466 15822 20478 15874
rect 22418 15822 22430 15874
rect 22482 15822 22494 15874
rect 29138 15822 29150 15874
rect 29202 15822 29214 15874
rect 14926 15810 14978 15822
rect 34638 15810 34690 15822
rect 1344 15706 38640 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 38640 15706
rect 1344 15620 38640 15654
rect 7534 15538 7586 15550
rect 7534 15474 7586 15486
rect 8990 15538 9042 15550
rect 8990 15474 9042 15486
rect 11678 15538 11730 15550
rect 11678 15474 11730 15486
rect 12686 15538 12738 15550
rect 12686 15474 12738 15486
rect 16494 15538 16546 15550
rect 16494 15474 16546 15486
rect 17278 15538 17330 15550
rect 17278 15474 17330 15486
rect 18958 15538 19010 15550
rect 23102 15538 23154 15550
rect 21298 15486 21310 15538
rect 21362 15486 21374 15538
rect 18958 15474 19010 15486
rect 23102 15474 23154 15486
rect 23886 15538 23938 15550
rect 23886 15474 23938 15486
rect 23998 15538 24050 15550
rect 23998 15474 24050 15486
rect 25342 15538 25394 15550
rect 25342 15474 25394 15486
rect 26238 15538 26290 15550
rect 26238 15474 26290 15486
rect 27358 15538 27410 15550
rect 27358 15474 27410 15486
rect 28702 15538 28754 15550
rect 28702 15474 28754 15486
rect 32286 15538 32338 15550
rect 32286 15474 32338 15486
rect 19294 15426 19346 15438
rect 13906 15374 13918 15426
rect 13970 15374 13982 15426
rect 17826 15374 17838 15426
rect 17890 15374 17902 15426
rect 18162 15374 18174 15426
rect 18226 15374 18238 15426
rect 19294 15362 19346 15374
rect 19630 15426 19682 15438
rect 19630 15362 19682 15374
rect 22654 15426 22706 15438
rect 22654 15362 22706 15374
rect 24222 15426 24274 15438
rect 24222 15362 24274 15374
rect 26462 15426 26514 15438
rect 26462 15362 26514 15374
rect 6862 15314 6914 15326
rect 6862 15250 6914 15262
rect 7086 15314 7138 15326
rect 7086 15250 7138 15262
rect 10222 15314 10274 15326
rect 10222 15250 10274 15262
rect 10446 15314 10498 15326
rect 17502 15314 17554 15326
rect 13122 15262 13134 15314
rect 13186 15262 13198 15314
rect 10446 15250 10498 15262
rect 17502 15250 17554 15262
rect 19742 15314 19794 15326
rect 19742 15250 19794 15262
rect 20302 15314 20354 15326
rect 20302 15250 20354 15262
rect 21646 15314 21698 15326
rect 24110 15314 24162 15326
rect 22418 15262 22430 15314
rect 22482 15262 22494 15314
rect 24434 15262 24446 15314
rect 24498 15262 24510 15314
rect 26002 15262 26014 15314
rect 26066 15262 26078 15314
rect 26674 15262 26686 15314
rect 26738 15262 26750 15314
rect 27122 15262 27134 15314
rect 27186 15262 27198 15314
rect 29026 15262 29038 15314
rect 29090 15262 29102 15314
rect 21646 15250 21698 15262
rect 24110 15250 24162 15262
rect 18286 15202 18338 15214
rect 16034 15150 16046 15202
rect 16098 15150 16110 15202
rect 18286 15138 18338 15150
rect 19406 15202 19458 15214
rect 19406 15138 19458 15150
rect 21870 15202 21922 15214
rect 21870 15138 21922 15150
rect 26350 15202 26402 15214
rect 29698 15150 29710 15202
rect 29762 15150 29774 15202
rect 31826 15150 31838 15202
rect 31890 15150 31902 15202
rect 26350 15138 26402 15150
rect 6514 15038 6526 15090
rect 6578 15038 6590 15090
rect 9874 15038 9886 15090
rect 9938 15038 9950 15090
rect 1344 14922 38640 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 38640 14922
rect 1344 14836 38640 14870
rect 25890 14702 25902 14754
rect 25954 14751 25966 14754
rect 26338 14751 26350 14754
rect 25954 14705 26350 14751
rect 25954 14702 25966 14705
rect 26338 14702 26350 14705
rect 26402 14702 26414 14754
rect 27346 14702 27358 14754
rect 27410 14702 27422 14754
rect 14702 14642 14754 14654
rect 14702 14578 14754 14590
rect 18958 14642 19010 14654
rect 25454 14642 25506 14654
rect 22530 14590 22542 14642
rect 22594 14590 22606 14642
rect 24658 14590 24670 14642
rect 24722 14590 24734 14642
rect 18958 14578 19010 14590
rect 25454 14578 25506 14590
rect 25902 14642 25954 14654
rect 25902 14578 25954 14590
rect 26462 14642 26514 14654
rect 26462 14578 26514 14590
rect 30606 14642 30658 14654
rect 30606 14578 30658 14590
rect 30942 14642 30994 14654
rect 30942 14578 30994 14590
rect 31166 14642 31218 14654
rect 34738 14590 34750 14642
rect 34802 14590 34814 14642
rect 31166 14578 31218 14590
rect 6302 14530 6354 14542
rect 6302 14466 6354 14478
rect 14478 14530 14530 14542
rect 26798 14530 26850 14542
rect 17490 14478 17502 14530
rect 17554 14478 17566 14530
rect 21858 14478 21870 14530
rect 21922 14478 21934 14530
rect 14478 14466 14530 14478
rect 26798 14466 26850 14478
rect 27022 14530 27074 14542
rect 27022 14466 27074 14478
rect 29262 14530 29314 14542
rect 31938 14478 31950 14530
rect 32002 14478 32014 14530
rect 29262 14466 29314 14478
rect 17726 14418 17778 14430
rect 17726 14354 17778 14366
rect 29598 14418 29650 14430
rect 32610 14366 32622 14418
rect 32674 14366 32686 14418
rect 29598 14354 29650 14366
rect 5966 14306 6018 14318
rect 15150 14306 15202 14318
rect 14130 14254 14142 14306
rect 14194 14254 14206 14306
rect 31490 14254 31502 14306
rect 31554 14254 31566 14306
rect 5966 14242 6018 14254
rect 15150 14242 15202 14254
rect 1344 14138 38640 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 38640 14138
rect 1344 14052 38640 14086
rect 33070 13970 33122 13982
rect 17602 13918 17614 13970
rect 17666 13918 17678 13970
rect 33070 13906 33122 13918
rect 9550 13858 9602 13870
rect 5394 13806 5406 13858
rect 5458 13806 5470 13858
rect 9550 13794 9602 13806
rect 9886 13858 9938 13870
rect 9886 13794 9938 13806
rect 7982 13746 8034 13758
rect 4722 13694 4734 13746
rect 4786 13694 4798 13746
rect 33282 13694 33294 13746
rect 33346 13694 33358 13746
rect 7982 13682 8034 13694
rect 17950 13634 18002 13646
rect 7522 13582 7534 13634
rect 7586 13582 7598 13634
rect 17950 13570 18002 13582
rect 18174 13634 18226 13646
rect 18174 13570 18226 13582
rect 18622 13634 18674 13646
rect 18622 13570 18674 13582
rect 25342 13634 25394 13646
rect 25342 13570 25394 13582
rect 31502 13634 31554 13646
rect 31502 13570 31554 13582
rect 1344 13354 38640 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 38640 13354
rect 1344 13268 38640 13302
rect 24558 13186 24610 13198
rect 24558 13122 24610 13134
rect 31166 13186 31218 13198
rect 31166 13122 31218 13134
rect 7198 13074 7250 13086
rect 17054 13074 17106 13086
rect 8306 13022 8318 13074
rect 8370 13022 8382 13074
rect 10434 13022 10446 13074
rect 10498 13022 10510 13074
rect 7198 13010 7250 13022
rect 17054 13010 17106 13022
rect 17502 13074 17554 13086
rect 17502 13010 17554 13022
rect 18286 13074 18338 13086
rect 18286 13010 18338 13022
rect 24782 13074 24834 13086
rect 24782 13010 24834 13022
rect 25230 13074 25282 13086
rect 25230 13010 25282 13022
rect 30270 13074 30322 13086
rect 30270 13010 30322 13022
rect 13806 12962 13858 12974
rect 7634 12910 7646 12962
rect 7698 12910 7710 12962
rect 30706 12910 30718 12962
rect 30770 12910 30782 12962
rect 13806 12898 13858 12910
rect 10894 12738 10946 12750
rect 10894 12674 10946 12686
rect 13470 12738 13522 12750
rect 13470 12674 13522 12686
rect 18958 12738 19010 12750
rect 24210 12686 24222 12738
rect 24274 12686 24286 12738
rect 18958 12674 19010 12686
rect 1344 12570 38640 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 38640 12570
rect 1344 12484 38640 12518
rect 8094 12402 8146 12414
rect 6626 12350 6638 12402
rect 6690 12350 6702 12402
rect 8094 12338 8146 12350
rect 12238 12402 12290 12414
rect 12238 12338 12290 12350
rect 13358 12402 13410 12414
rect 13358 12338 13410 12350
rect 13806 12402 13858 12414
rect 13806 12338 13858 12350
rect 15038 12402 15090 12414
rect 15038 12338 15090 12350
rect 15486 12402 15538 12414
rect 15486 12338 15538 12350
rect 16158 12402 16210 12414
rect 16158 12338 16210 12350
rect 17278 12402 17330 12414
rect 17278 12338 17330 12350
rect 18846 12402 18898 12414
rect 18846 12338 18898 12350
rect 6302 12290 6354 12302
rect 6302 12226 6354 12238
rect 12014 12290 12066 12302
rect 12014 12226 12066 12238
rect 19070 12290 19122 12302
rect 19070 12226 19122 12238
rect 24222 12290 24274 12302
rect 24222 12226 24274 12238
rect 6974 12178 7026 12190
rect 6066 12126 6078 12178
rect 6130 12126 6142 12178
rect 6974 12114 7026 12126
rect 8430 12178 8482 12190
rect 8430 12114 8482 12126
rect 9886 12178 9938 12190
rect 9886 12114 9938 12126
rect 12462 12178 12514 12190
rect 16270 12178 16322 12190
rect 12674 12126 12686 12178
rect 12738 12126 12750 12178
rect 15922 12126 15934 12178
rect 15986 12126 15998 12178
rect 12462 12114 12514 12126
rect 16270 12114 16322 12126
rect 16382 12178 16434 12190
rect 17502 12178 17554 12190
rect 16594 12126 16606 12178
rect 16658 12126 16670 12178
rect 16382 12114 16434 12126
rect 17502 12114 17554 12126
rect 17950 12178 18002 12190
rect 17950 12114 18002 12126
rect 18062 12178 18114 12190
rect 18610 12126 18622 12178
rect 18674 12126 18686 12178
rect 19282 12126 19294 12178
rect 19346 12126 19358 12178
rect 23762 12126 23774 12178
rect 23826 12126 23838 12178
rect 29698 12126 29710 12178
rect 29762 12126 29774 12178
rect 18062 12114 18114 12126
rect 7198 12066 7250 12078
rect 7198 12002 7250 12014
rect 7646 12066 7698 12078
rect 7646 12002 7698 12014
rect 8990 12066 9042 12078
rect 8990 12002 9042 12014
rect 10110 12066 10162 12078
rect 10110 12002 10162 12014
rect 12350 12066 12402 12078
rect 12350 12002 12402 12014
rect 18286 12066 18338 12078
rect 18286 12002 18338 12014
rect 18958 12066 19010 12078
rect 18958 12002 19010 12014
rect 19742 12066 19794 12078
rect 30158 12066 30210 12078
rect 20850 12014 20862 12066
rect 20914 12014 20926 12066
rect 22978 12014 22990 12066
rect 23042 12014 23054 12066
rect 26786 12014 26798 12066
rect 26850 12014 26862 12066
rect 28914 12014 28926 12066
rect 28978 12014 28990 12066
rect 19742 12002 19794 12014
rect 30158 12002 30210 12014
rect 9538 11902 9550 11954
rect 9602 11902 9614 11954
rect 29922 11902 29934 11954
rect 29986 11951 29998 11954
rect 30146 11951 30158 11954
rect 29986 11905 30158 11951
rect 29986 11902 29998 11905
rect 30146 11902 30158 11905
rect 30210 11902 30222 11954
rect 1344 11786 38640 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 38640 11786
rect 1344 11700 38640 11734
rect 14478 11618 14530 11630
rect 14478 11554 14530 11566
rect 12910 11506 12962 11518
rect 6962 11454 6974 11506
rect 7026 11454 7038 11506
rect 12002 11454 12014 11506
rect 12066 11454 12078 11506
rect 12910 11442 12962 11454
rect 14814 11506 14866 11518
rect 19182 11506 19234 11518
rect 18722 11454 18734 11506
rect 18786 11454 18798 11506
rect 14814 11442 14866 11454
rect 19182 11442 19234 11454
rect 20750 11506 20802 11518
rect 20750 11442 20802 11454
rect 25902 11506 25954 11518
rect 25902 11442 25954 11454
rect 26350 11506 26402 11518
rect 26350 11442 26402 11454
rect 27134 11506 27186 11518
rect 30258 11454 30270 11506
rect 30322 11454 30334 11506
rect 27134 11442 27186 11454
rect 20190 11394 20242 11406
rect 5618 11342 5630 11394
rect 5682 11342 5694 11394
rect 9090 11342 9102 11394
rect 9154 11342 9166 11394
rect 15362 11342 15374 11394
rect 15426 11342 15438 11394
rect 15810 11342 15822 11394
rect 15874 11342 15886 11394
rect 19618 11342 19630 11394
rect 19682 11342 19694 11394
rect 20190 11330 20242 11342
rect 21422 11394 21474 11406
rect 21422 11330 21474 11342
rect 21758 11394 21810 11406
rect 22306 11342 22318 11394
rect 22370 11342 22382 11394
rect 24322 11342 24334 11394
rect 24386 11342 24398 11394
rect 33058 11342 33070 11394
rect 33122 11342 33134 11394
rect 21758 11330 21810 11342
rect 14254 11282 14306 11294
rect 19966 11282 20018 11294
rect 9874 11230 9886 11282
rect 9938 11230 9950 11282
rect 16594 11230 16606 11282
rect 16658 11230 16670 11282
rect 19730 11230 19742 11282
rect 19794 11230 19806 11282
rect 14254 11218 14306 11230
rect 19966 11218 20018 11230
rect 21310 11282 21362 11294
rect 21310 11218 21362 11230
rect 21646 11282 21698 11294
rect 21646 11218 21698 11230
rect 22542 11282 22594 11294
rect 22542 11218 22594 11230
rect 27694 11282 27746 11294
rect 27694 11218 27746 11230
rect 28030 11282 28082 11294
rect 32386 11230 32398 11282
rect 32450 11230 32462 11282
rect 28030 11218 28082 11230
rect 12462 11170 12514 11182
rect 12462 11106 12514 11118
rect 15150 11170 15202 11182
rect 15150 11106 15202 11118
rect 24110 11170 24162 11182
rect 24110 11106 24162 11118
rect 29934 11170 29986 11182
rect 29934 11106 29986 11118
rect 1344 11002 38640 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 38640 11002
rect 1344 10916 38640 10950
rect 8990 10834 9042 10846
rect 8990 10770 9042 10782
rect 9886 10834 9938 10846
rect 9886 10770 9938 10782
rect 10670 10834 10722 10846
rect 10670 10770 10722 10782
rect 10782 10834 10834 10846
rect 10782 10770 10834 10782
rect 11342 10834 11394 10846
rect 11342 10770 11394 10782
rect 11790 10834 11842 10846
rect 11790 10770 11842 10782
rect 16158 10834 16210 10846
rect 16158 10770 16210 10782
rect 17838 10834 17890 10846
rect 17838 10770 17890 10782
rect 20638 10834 20690 10846
rect 20638 10770 20690 10782
rect 21534 10834 21586 10846
rect 22878 10834 22930 10846
rect 22418 10782 22430 10834
rect 22482 10782 22494 10834
rect 21534 10770 21586 10782
rect 22878 10770 22930 10782
rect 24222 10834 24274 10846
rect 24222 10770 24274 10782
rect 25342 10834 25394 10846
rect 25342 10770 25394 10782
rect 25454 10834 25506 10846
rect 25454 10770 25506 10782
rect 26798 10834 26850 10846
rect 31390 10834 31442 10846
rect 27458 10782 27470 10834
rect 27522 10782 27534 10834
rect 26798 10770 26850 10782
rect 31390 10770 31442 10782
rect 9550 10722 9602 10734
rect 19742 10722 19794 10734
rect 5282 10670 5294 10722
rect 5346 10670 5358 10722
rect 6402 10670 6414 10722
rect 6466 10670 6478 10722
rect 12898 10670 12910 10722
rect 12962 10670 12974 10722
rect 9550 10658 9602 10670
rect 19742 10658 19794 10670
rect 20526 10722 20578 10734
rect 20526 10658 20578 10670
rect 10446 10610 10498 10622
rect 18062 10610 18114 10622
rect 5730 10558 5742 10610
rect 5794 10558 5806 10610
rect 10210 10558 10222 10610
rect 10274 10558 10286 10610
rect 12114 10558 12126 10610
rect 12178 10558 12190 10610
rect 15810 10558 15822 10610
rect 15874 10558 15886 10610
rect 10446 10546 10498 10558
rect 18062 10546 18114 10558
rect 18510 10610 18562 10622
rect 18510 10546 18562 10558
rect 18622 10610 18674 10622
rect 18622 10546 18674 10558
rect 18846 10610 18898 10622
rect 18846 10546 18898 10558
rect 19294 10610 19346 10622
rect 19294 10546 19346 10558
rect 19630 10610 19682 10622
rect 19630 10546 19682 10558
rect 19966 10610 20018 10622
rect 19966 10546 20018 10558
rect 20190 10610 20242 10622
rect 20190 10546 20242 10558
rect 20750 10610 20802 10622
rect 20750 10546 20802 10558
rect 20974 10610 21026 10622
rect 20974 10546 21026 10558
rect 22094 10610 22146 10622
rect 22094 10546 22146 10558
rect 24670 10610 24722 10622
rect 24670 10546 24722 10558
rect 25678 10610 25730 10622
rect 25678 10546 25730 10558
rect 25790 10610 25842 10622
rect 26686 10610 26738 10622
rect 26450 10558 26462 10610
rect 26514 10558 26526 10610
rect 25790 10546 25842 10558
rect 26686 10546 26738 10558
rect 26910 10610 26962 10622
rect 27122 10558 27134 10610
rect 27186 10558 27198 10610
rect 31154 10558 31166 10610
rect 31218 10558 31230 10610
rect 26910 10546 26962 10558
rect 4286 10498 4338 10510
rect 17502 10498 17554 10510
rect 8530 10446 8542 10498
rect 8594 10446 8606 10498
rect 10658 10446 10670 10498
rect 10722 10446 10734 10498
rect 15026 10446 15038 10498
rect 15090 10446 15102 10498
rect 4286 10434 4338 10446
rect 17502 10434 17554 10446
rect 21870 10498 21922 10510
rect 28030 10498 28082 10510
rect 25330 10446 25342 10498
rect 25394 10446 25406 10498
rect 21870 10434 21922 10446
rect 28030 10434 28082 10446
rect 27806 10386 27858 10398
rect 11330 10334 11342 10386
rect 11394 10383 11406 10386
rect 11554 10383 11566 10386
rect 11394 10337 11566 10383
rect 11394 10334 11406 10337
rect 11554 10334 11566 10337
rect 11618 10334 11630 10386
rect 27806 10322 27858 10334
rect 1344 10218 38640 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 38640 10218
rect 1344 10132 38640 10166
rect 11330 9998 11342 10050
rect 11394 10047 11406 10050
rect 12002 10047 12014 10050
rect 11394 10001 12014 10047
rect 11394 9998 11406 10001
rect 12002 9998 12014 10001
rect 12066 9998 12078 10050
rect 27234 9998 27246 10050
rect 27298 10047 27310 10050
rect 28018 10047 28030 10050
rect 27298 10001 28030 10047
rect 27298 9998 27310 10001
rect 28018 9998 28030 10001
rect 28082 9998 28094 10050
rect 31154 9998 31166 10050
rect 31218 9998 31230 10050
rect 11566 9938 11618 9950
rect 4722 9886 4734 9938
rect 4786 9886 4798 9938
rect 10994 9886 11006 9938
rect 11058 9886 11070 9938
rect 11566 9874 11618 9886
rect 12014 9938 12066 9950
rect 16830 9938 16882 9950
rect 18286 9938 18338 9950
rect 14242 9886 14254 9938
rect 14306 9886 14318 9938
rect 16370 9886 16382 9938
rect 16434 9886 16446 9938
rect 17602 9886 17614 9938
rect 17666 9886 17678 9938
rect 12014 9874 12066 9886
rect 16830 9874 16882 9886
rect 18286 9874 18338 9886
rect 18958 9938 19010 9950
rect 18958 9874 19010 9886
rect 19406 9938 19458 9950
rect 19406 9874 19458 9886
rect 19854 9938 19906 9950
rect 19854 9874 19906 9886
rect 20078 9938 20130 9950
rect 27470 9938 27522 9950
rect 23874 9886 23886 9938
rect 23938 9886 23950 9938
rect 26002 9886 26014 9938
rect 26066 9886 26078 9938
rect 26450 9886 26462 9938
rect 26514 9886 26526 9938
rect 20078 9874 20130 9886
rect 27470 9874 27522 9886
rect 27918 9938 27970 9950
rect 31726 9938 31778 9950
rect 30034 9886 30046 9938
rect 30098 9886 30110 9938
rect 27918 9874 27970 9886
rect 31726 9874 31778 9886
rect 10670 9826 10722 9838
rect 17726 9826 17778 9838
rect 5618 9774 5630 9826
rect 5682 9774 5694 9826
rect 10434 9774 10446 9826
rect 10498 9774 10510 9826
rect 11106 9774 11118 9826
rect 11170 9774 11182 9826
rect 13458 9774 13470 9826
rect 13522 9774 13534 9826
rect 17154 9774 17166 9826
rect 17218 9774 17230 9826
rect 10670 9762 10722 9774
rect 17726 9762 17778 9774
rect 20302 9826 20354 9838
rect 26798 9826 26850 9838
rect 31502 9826 31554 9838
rect 23090 9774 23102 9826
rect 23154 9774 23166 9826
rect 26338 9774 26350 9826
rect 26402 9774 26414 9826
rect 29698 9774 29710 9826
rect 29762 9774 29774 9826
rect 20302 9762 20354 9774
rect 26798 9762 26850 9774
rect 31502 9762 31554 9774
rect 32174 9826 32226 9838
rect 32174 9762 32226 9774
rect 5070 9714 5122 9726
rect 27022 9714 27074 9726
rect 7410 9662 7422 9714
rect 7474 9662 7486 9714
rect 5070 9650 5122 9662
rect 27022 9650 27074 9662
rect 30830 9714 30882 9726
rect 30830 9650 30882 9662
rect 10894 9602 10946 9614
rect 10894 9538 10946 9550
rect 17390 9602 17442 9614
rect 17390 9538 17442 9550
rect 17614 9602 17666 9614
rect 26574 9602 26626 9614
rect 20626 9550 20638 9602
rect 20690 9550 20702 9602
rect 17614 9538 17666 9550
rect 26574 9538 26626 9550
rect 28366 9602 28418 9614
rect 28366 9538 28418 9550
rect 1344 9434 38640 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 38640 9434
rect 1344 9348 38640 9382
rect 8990 9266 9042 9278
rect 8990 9202 9042 9214
rect 15710 9266 15762 9278
rect 15710 9202 15762 9214
rect 18174 9266 18226 9278
rect 18174 9202 18226 9214
rect 20526 9154 20578 9166
rect 20526 9090 20578 9102
rect 9886 9042 9938 9054
rect 9886 8978 9938 8990
rect 10110 9042 10162 9054
rect 16830 9042 16882 9054
rect 32510 9042 32562 9054
rect 15474 8990 15486 9042
rect 15538 8990 15550 9042
rect 20290 8990 20302 9042
rect 20354 8990 20366 9042
rect 25442 8990 25454 9042
rect 25506 8990 25518 9042
rect 31938 8990 31950 9042
rect 32002 8990 32014 9042
rect 38210 8990 38222 9042
rect 38274 8990 38286 9042
rect 10110 8978 10162 8990
rect 16830 8978 16882 8990
rect 32510 8978 32562 8990
rect 5294 8930 5346 8942
rect 19742 8930 19794 8942
rect 28702 8930 28754 8942
rect 37214 8930 37266 8942
rect 16258 8878 16270 8930
rect 16322 8878 16334 8930
rect 26114 8878 26126 8930
rect 26178 8878 26190 8930
rect 28242 8878 28254 8930
rect 28306 8878 28318 8930
rect 29138 8878 29150 8930
rect 29202 8878 29214 8930
rect 31266 8878 31278 8930
rect 31330 8878 31342 8930
rect 5294 8866 5346 8878
rect 19742 8866 19794 8878
rect 28702 8866 28754 8878
rect 37214 8866 37266 8878
rect 16606 8818 16658 8830
rect 9538 8766 9550 8818
rect 9602 8766 9614 8818
rect 16606 8754 16658 8766
rect 1344 8650 38640 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 38640 8650
rect 1344 8564 38640 8598
rect 29934 8482 29986 8494
rect 29934 8418 29986 8430
rect 26126 8370 26178 8382
rect 26126 8306 26178 8318
rect 27582 8370 27634 8382
rect 27582 8306 27634 8318
rect 38334 8370 38386 8382
rect 38334 8306 38386 8318
rect 8878 8258 8930 8270
rect 26350 8258 26402 8270
rect 27358 8258 27410 8270
rect 31278 8258 31330 8270
rect 25554 8206 25566 8258
rect 25618 8206 25630 8258
rect 27010 8206 27022 8258
rect 27074 8206 27086 8258
rect 29586 8206 29598 8258
rect 29650 8206 29662 8258
rect 8878 8194 8930 8206
rect 26350 8194 26402 8206
rect 27358 8194 27410 8206
rect 31278 8194 31330 8206
rect 31502 8258 31554 8270
rect 31502 8194 31554 8206
rect 25790 8146 25842 8158
rect 25790 8082 25842 8094
rect 8542 8034 8594 8046
rect 8542 7970 8594 7982
rect 15934 8034 15986 8046
rect 15934 7970 15986 7982
rect 25118 8034 25170 8046
rect 28030 8034 28082 8046
rect 31950 8034 32002 8046
rect 26674 7982 26686 8034
rect 26738 7982 26750 8034
rect 30930 7982 30942 8034
rect 30994 7982 31006 8034
rect 25118 7970 25170 7982
rect 28030 7970 28082 7982
rect 31950 7970 32002 7982
rect 1344 7866 38640 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 38640 7866
rect 1344 7780 38640 7814
rect 10670 7698 10722 7710
rect 10670 7634 10722 7646
rect 14478 7698 14530 7710
rect 14478 7634 14530 7646
rect 30830 7698 30882 7710
rect 30830 7634 30882 7646
rect 31390 7698 31442 7710
rect 31390 7634 31442 7646
rect 10222 7586 10274 7598
rect 26910 7586 26962 7598
rect 21186 7534 21198 7586
rect 21250 7534 21262 7586
rect 28018 7534 28030 7586
rect 28082 7534 28094 7586
rect 10222 7522 10274 7534
rect 26910 7522 26962 7534
rect 5954 7422 5966 7474
rect 6018 7422 6030 7474
rect 9986 7422 9998 7474
rect 10050 7422 10062 7474
rect 11106 7422 11118 7474
rect 11170 7422 11182 7474
rect 21970 7422 21982 7474
rect 22034 7422 22046 7474
rect 26674 7422 26686 7474
rect 26738 7422 26750 7474
rect 27234 7422 27246 7474
rect 27298 7422 27310 7474
rect 30594 7422 30606 7474
rect 30658 7422 30670 7474
rect 7422 7362 7474 7374
rect 22430 7362 22482 7374
rect 6626 7310 6638 7362
rect 6690 7310 6702 7362
rect 11890 7310 11902 7362
rect 11954 7310 11966 7362
rect 14018 7310 14030 7362
rect 14082 7310 14094 7362
rect 19058 7310 19070 7362
rect 19122 7310 19134 7362
rect 30146 7310 30158 7362
rect 30210 7310 30222 7362
rect 7422 7298 7474 7310
rect 22430 7298 22482 7310
rect 1344 7082 38640 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 38640 7082
rect 1344 6996 38640 7030
rect 10782 6914 10834 6926
rect 10782 6850 10834 6862
rect 12126 6914 12178 6926
rect 12126 6850 12178 6862
rect 14366 6914 14418 6926
rect 14366 6850 14418 6862
rect 11006 6802 11058 6814
rect 10098 6750 10110 6802
rect 10162 6750 10174 6802
rect 11006 6738 11058 6750
rect 11454 6802 11506 6814
rect 11454 6738 11506 6750
rect 13694 6802 13746 6814
rect 13694 6738 13746 6750
rect 14590 6802 14642 6814
rect 17826 6750 17838 6802
rect 17890 6750 17902 6802
rect 14590 6738 14642 6750
rect 12350 6690 12402 6702
rect 18286 6690 18338 6702
rect 7298 6638 7310 6690
rect 7362 6638 7374 6690
rect 7970 6638 7982 6690
rect 8034 6638 8046 6690
rect 10434 6638 10446 6690
rect 10498 6638 10510 6690
rect 15026 6638 15038 6690
rect 15090 6638 15102 6690
rect 12350 6626 12402 6638
rect 18286 6626 18338 6638
rect 23550 6690 23602 6702
rect 23550 6626 23602 6638
rect 30382 6690 30434 6702
rect 30382 6626 30434 6638
rect 15698 6526 15710 6578
rect 15762 6526 15774 6578
rect 21870 6466 21922 6478
rect 11778 6414 11790 6466
rect 11842 6414 11854 6466
rect 14018 6414 14030 6466
rect 14082 6414 14094 6466
rect 21870 6402 21922 6414
rect 22318 6466 22370 6478
rect 22318 6402 22370 6414
rect 24894 6466 24946 6478
rect 24894 6402 24946 6414
rect 1344 6298 38640 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 38640 6298
rect 1344 6212 38640 6246
rect 16270 6130 16322 6142
rect 16270 6066 16322 6078
rect 17390 6018 17442 6030
rect 17390 5954 17442 5966
rect 24222 5906 24274 5918
rect 9650 5854 9662 5906
rect 9714 5854 9726 5906
rect 13010 5854 13022 5906
rect 13074 5854 13086 5906
rect 17602 5854 17614 5906
rect 17666 5854 17678 5906
rect 18946 5854 18958 5906
rect 19010 5854 19022 5906
rect 22194 5854 22206 5906
rect 22258 5854 22270 5906
rect 24222 5842 24274 5854
rect 24446 5906 24498 5918
rect 24446 5842 24498 5854
rect 25566 5906 25618 5918
rect 25566 5842 25618 5854
rect 25790 5906 25842 5918
rect 25790 5842 25842 5854
rect 23214 5794 23266 5806
rect 10322 5742 10334 5794
rect 10386 5742 10398 5794
rect 12450 5742 12462 5794
rect 12514 5742 12526 5794
rect 13682 5742 13694 5794
rect 13746 5742 13758 5794
rect 15810 5742 15822 5794
rect 15874 5742 15886 5794
rect 19618 5742 19630 5794
rect 19682 5742 19694 5794
rect 21746 5742 21758 5794
rect 21810 5742 21822 5794
rect 23214 5730 23266 5742
rect 23874 5630 23886 5682
rect 23938 5630 23950 5682
rect 25218 5630 25230 5682
rect 25282 5630 25294 5682
rect 1344 5514 38640 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 38640 5514
rect 1344 5428 38640 5462
rect 20414 5346 20466 5358
rect 20414 5282 20466 5294
rect 21534 5346 21586 5358
rect 21534 5282 21586 5294
rect 9326 5234 9378 5246
rect 9326 5170 9378 5182
rect 10110 5234 10162 5246
rect 10110 5170 10162 5182
rect 12798 5234 12850 5246
rect 12798 5170 12850 5182
rect 15934 5234 15986 5246
rect 19742 5234 19794 5246
rect 17042 5182 17054 5234
rect 17106 5182 17118 5234
rect 19170 5182 19182 5234
rect 19234 5182 19246 5234
rect 15934 5170 15986 5182
rect 19742 5170 19794 5182
rect 20638 5234 20690 5246
rect 20638 5170 20690 5182
rect 21310 5234 21362 5246
rect 21310 5170 21362 5182
rect 23102 5234 23154 5246
rect 27010 5182 27022 5234
rect 27074 5182 27086 5234
rect 23102 5170 23154 5182
rect 8654 5122 8706 5134
rect 15038 5122 15090 5134
rect 12114 5070 12126 5122
rect 12178 5070 12190 5122
rect 14466 5070 14478 5122
rect 14530 5070 14542 5122
rect 8654 5058 8706 5070
rect 15038 5058 15090 5070
rect 15710 5122 15762 5134
rect 16370 5070 16382 5122
rect 16434 5070 16446 5122
rect 21858 5070 21870 5122
rect 21922 5070 21934 5122
rect 22418 5070 22430 5122
rect 22482 5070 22494 5122
rect 23538 5070 23550 5122
rect 23602 5070 23614 5122
rect 24210 5070 24222 5122
rect 24274 5070 24286 5122
rect 15710 5058 15762 5070
rect 8318 5010 8370 5022
rect 8318 4946 8370 4958
rect 14254 5010 14306 5022
rect 27470 5010 27522 5022
rect 24882 4958 24894 5010
rect 24946 4958 24958 5010
rect 14254 4946 14306 4958
rect 27470 4946 27522 4958
rect 7982 4898 8034 4910
rect 7982 4834 8034 4846
rect 8766 4898 8818 4910
rect 8766 4834 8818 4846
rect 8990 4898 9042 4910
rect 8990 4834 9042 4846
rect 11902 4898 11954 4910
rect 11902 4834 11954 4846
rect 14030 4898 14082 4910
rect 22206 4898 22258 4910
rect 15362 4846 15374 4898
rect 15426 4846 15438 4898
rect 20066 4846 20078 4898
rect 20130 4846 20142 4898
rect 14030 4834 14082 4846
rect 22206 4834 22258 4846
rect 23774 4898 23826 4910
rect 23774 4834 23826 4846
rect 1344 4730 38640 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 38640 4730
rect 1344 4644 38640 4678
rect 8990 4562 9042 4574
rect 8990 4498 9042 4510
rect 9774 4562 9826 4574
rect 9774 4498 9826 4510
rect 11342 4562 11394 4574
rect 11342 4498 11394 4510
rect 15822 4562 15874 4574
rect 15822 4498 15874 4510
rect 16830 4562 16882 4574
rect 19070 4562 19122 4574
rect 17378 4510 17390 4562
rect 17442 4510 17454 4562
rect 16830 4498 16882 4510
rect 19070 4498 19122 4510
rect 19630 4562 19682 4574
rect 19630 4498 19682 4510
rect 23326 4562 23378 4574
rect 23326 4498 23378 4510
rect 24670 4562 24722 4574
rect 24670 4498 24722 4510
rect 10222 4450 10274 4462
rect 14030 4450 14082 4462
rect 7746 4398 7758 4450
rect 7810 4398 7822 4450
rect 10882 4398 10894 4450
rect 10946 4398 10958 4450
rect 22082 4398 22094 4450
rect 22146 4398 22158 4450
rect 25218 4398 25230 4450
rect 25282 4398 25294 4450
rect 25554 4398 25566 4450
rect 25618 4398 25630 4450
rect 10222 4386 10274 4398
rect 14030 4386 14082 4398
rect 10110 4338 10162 4350
rect 8530 4286 8542 4338
rect 8594 4286 8606 4338
rect 10110 4274 10162 4286
rect 10446 4338 10498 4350
rect 17726 4338 17778 4350
rect 10770 4286 10782 4338
rect 10834 4286 10846 4338
rect 14578 4286 14590 4338
rect 14642 4286 14654 4338
rect 16034 4286 16046 4338
rect 16098 4286 16110 4338
rect 10446 4274 10498 4286
rect 17726 4274 17778 4286
rect 17950 4338 18002 4350
rect 19394 4286 19406 4338
rect 19458 4286 19470 4338
rect 22866 4286 22878 4338
rect 22930 4286 22942 4338
rect 24434 4286 24446 4338
rect 24498 4286 24510 4338
rect 25890 4286 25902 4338
rect 25954 4286 25966 4338
rect 34402 4286 34414 4338
rect 34466 4286 34478 4338
rect 34738 4286 34750 4338
rect 34802 4286 34814 4338
rect 17950 4274 18002 4286
rect 15038 4226 15090 4238
rect 5618 4174 5630 4226
rect 5682 4174 5694 4226
rect 15038 4162 15090 4174
rect 15486 4226 15538 4238
rect 15486 4162 15538 4174
rect 18398 4226 18450 4238
rect 26462 4226 26514 4238
rect 19954 4174 19966 4226
rect 20018 4174 20030 4226
rect 34514 4174 34526 4226
rect 34578 4174 34590 4226
rect 18398 4162 18450 4174
rect 26462 4162 26514 4174
rect 33954 4062 33966 4114
rect 34018 4062 34030 4114
rect 1344 3946 38640 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 38640 3946
rect 1344 3860 38640 3894
rect 12574 3666 12626 3678
rect 26574 3666 26626 3678
rect 8082 3614 8094 3666
rect 8146 3614 8158 3666
rect 10434 3614 10446 3666
rect 10498 3614 10510 3666
rect 23874 3614 23886 3666
rect 23938 3614 23950 3666
rect 26002 3614 26014 3666
rect 26066 3614 26078 3666
rect 12574 3602 12626 3614
rect 26574 3602 26626 3614
rect 18174 3554 18226 3566
rect 33182 3554 33234 3566
rect 8306 3502 8318 3554
rect 8370 3502 8382 3554
rect 8530 3502 8542 3554
rect 8594 3502 8606 3554
rect 10098 3502 10110 3554
rect 10162 3502 10174 3554
rect 10322 3502 10334 3554
rect 10386 3502 10398 3554
rect 14802 3502 14814 3554
rect 14866 3502 14878 3554
rect 15474 3502 15486 3554
rect 15538 3502 15550 3554
rect 16034 3502 16046 3554
rect 16098 3502 16110 3554
rect 23202 3502 23214 3554
rect 23266 3502 23278 3554
rect 27458 3502 27470 3554
rect 27522 3502 27534 3554
rect 27906 3502 27918 3554
rect 27970 3502 27982 3554
rect 31042 3502 31054 3554
rect 31106 3502 31118 3554
rect 18174 3490 18226 3502
rect 33182 3490 33234 3502
rect 6190 3442 6242 3454
rect 6190 3378 6242 3390
rect 6302 3442 6354 3454
rect 11118 3442 11170 3454
rect 7410 3390 7422 3442
rect 7474 3390 7486 3442
rect 6302 3378 6354 3390
rect 11118 3378 11170 3390
rect 13694 3442 13746 3454
rect 13694 3378 13746 3390
rect 13918 3442 13970 3454
rect 13918 3378 13970 3390
rect 14254 3442 14306 3454
rect 14254 3378 14306 3390
rect 15038 3442 15090 3454
rect 15038 3378 15090 3390
rect 15710 3442 15762 3454
rect 15710 3378 15762 3390
rect 17166 3442 17218 3454
rect 17166 3378 17218 3390
rect 18622 3442 18674 3454
rect 33630 3442 33682 3454
rect 26898 3390 26910 3442
rect 26962 3390 26974 3442
rect 28466 3390 28478 3442
rect 28530 3390 28542 3442
rect 31154 3390 31166 3442
rect 31218 3390 31230 3442
rect 18622 3378 18674 3390
rect 33630 3378 33682 3390
rect 11454 3330 11506 3342
rect 11454 3266 11506 3278
rect 12126 3330 12178 3342
rect 20862 3330 20914 3342
rect 16146 3278 16158 3330
rect 16210 3278 16222 3330
rect 12126 3266 12178 3278
rect 20862 3266 20914 3278
rect 22654 3330 22706 3342
rect 27010 3278 27022 3330
rect 27074 3278 27086 3330
rect 33058 3278 33070 3330
rect 33122 3278 33134 3330
rect 22654 3266 22706 3278
rect 1344 3162 38640 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 38640 3162
rect 1344 3076 38640 3110
rect 17390 2994 17442 3006
rect 10546 2942 10558 2994
rect 10610 2942 10622 2994
rect 13682 2942 13694 2994
rect 13746 2942 13758 2994
rect 19842 2942 19854 2994
rect 19906 2942 19918 2994
rect 25890 2942 25902 2994
rect 25954 2942 25966 2994
rect 17390 2930 17442 2942
rect 15262 2882 15314 2894
rect 6402 2830 6414 2882
rect 6466 2830 6478 2882
rect 10098 2830 10110 2882
rect 10162 2830 10174 2882
rect 11554 2830 11566 2882
rect 11618 2830 11630 2882
rect 12786 2830 12798 2882
rect 12850 2830 12862 2882
rect 15262 2818 15314 2830
rect 20302 2882 20354 2894
rect 20302 2818 20354 2830
rect 22318 2882 22370 2894
rect 25330 2830 25342 2882
rect 25394 2830 25406 2882
rect 26786 2830 26798 2882
rect 26850 2830 26862 2882
rect 33954 2830 33966 2882
rect 34018 2830 34030 2882
rect 22318 2818 22370 2830
rect 11118 2770 11170 2782
rect 14814 2770 14866 2782
rect 18174 2770 18226 2782
rect 21870 2770 21922 2782
rect 26350 2770 26402 2782
rect 4610 2718 4622 2770
rect 4674 2718 4686 2770
rect 10546 2718 10558 2770
rect 10610 2718 10622 2770
rect 12674 2718 12686 2770
rect 12738 2718 12750 2770
rect 17602 2718 17614 2770
rect 17666 2718 17678 2770
rect 19730 2718 19742 2770
rect 19794 2718 19806 2770
rect 25218 2718 25230 2770
rect 25282 2718 25294 2770
rect 33058 2718 33070 2770
rect 33122 2718 33134 2770
rect 34738 2718 34750 2770
rect 34802 2718 34814 2770
rect 11118 2706 11170 2718
rect 14814 2706 14866 2718
rect 18174 2706 18226 2718
rect 21870 2706 21922 2718
rect 26350 2706 26402 2718
rect 7646 2658 7698 2670
rect 7646 2594 7698 2606
rect 8542 2658 8594 2670
rect 8542 2594 8594 2606
rect 9102 2658 9154 2670
rect 9102 2594 9154 2606
rect 9774 2658 9826 2670
rect 9774 2594 9826 2606
rect 12462 2658 12514 2670
rect 12462 2594 12514 2606
rect 19070 2658 19122 2670
rect 19070 2594 19122 2606
rect 19518 2658 19570 2670
rect 19518 2594 19570 2606
rect 24334 2658 24386 2670
rect 24334 2594 24386 2606
rect 24782 2658 24834 2670
rect 24782 2594 24834 2606
rect 27358 2658 27410 2670
rect 27358 2594 27410 2606
rect 27806 2658 27858 2670
rect 27806 2594 27858 2606
rect 28366 2658 28418 2670
rect 28366 2594 28418 2606
rect 28926 2658 28978 2670
rect 28926 2594 28978 2606
rect 29822 2658 29874 2670
rect 29822 2594 29874 2606
rect 30718 2658 30770 2670
rect 30718 2594 30770 2606
rect 31950 2658 32002 2670
rect 31950 2594 32002 2606
rect 32622 2658 32674 2670
rect 32622 2594 32674 2606
rect 36094 2658 36146 2670
rect 36094 2594 36146 2606
rect 36542 2658 36594 2670
rect 36542 2594 36594 2606
rect 33182 2546 33234 2558
rect 33182 2482 33234 2494
rect 1344 2378 38640 2412
rect 1344 2326 4478 2378
rect 4530 2326 4582 2378
rect 4634 2326 4686 2378
rect 4738 2326 35198 2378
rect 35250 2326 35302 2378
rect 35354 2326 35406 2378
rect 35458 2326 38640 2378
rect 1344 2292 38640 2326
rect 13246 2210 13298 2222
rect 13246 2146 13298 2158
rect 11230 1986 11282 1998
rect 16270 1986 16322 1998
rect 21086 1986 21138 1998
rect 8530 1934 8542 1986
rect 8594 1934 8606 1986
rect 10434 1934 10446 1986
rect 10498 1934 10510 1986
rect 11666 1934 11678 1986
rect 11730 1934 11742 1986
rect 12338 1934 12350 1986
rect 12402 1934 12414 1986
rect 13458 1934 13470 1986
rect 13522 1934 13534 1986
rect 17602 1934 17614 1986
rect 17666 1934 17678 1986
rect 11230 1922 11282 1934
rect 16270 1922 16322 1934
rect 21086 1922 21138 1934
rect 21982 1986 22034 1998
rect 21982 1922 22034 1934
rect 22878 1986 22930 1998
rect 22878 1922 22930 1934
rect 23662 1986 23714 1998
rect 32174 1986 32226 1998
rect 34862 1986 34914 1998
rect 26002 1934 26014 1986
rect 26066 1934 26078 1986
rect 27570 1934 27582 1986
rect 27634 1934 27646 1986
rect 29362 1934 29374 1986
rect 29426 1934 29438 1986
rect 33730 1934 33742 1986
rect 33794 1934 33806 1986
rect 23662 1922 23714 1934
rect 32174 1922 32226 1934
rect 34862 1922 34914 1934
rect 35310 1986 35362 1998
rect 36194 1934 36206 1986
rect 36258 1934 36270 1986
rect 36866 1934 36878 1986
rect 36930 1934 36942 1986
rect 35310 1922 35362 1934
rect 3838 1874 3890 1886
rect 3838 1810 3890 1822
rect 4062 1874 4114 1886
rect 4062 1810 4114 1822
rect 4398 1874 4450 1886
rect 4398 1810 4450 1822
rect 5854 1874 5906 1886
rect 5854 1810 5906 1822
rect 6190 1874 6242 1886
rect 7646 1874 7698 1886
rect 7074 1822 7086 1874
rect 7138 1822 7150 1874
rect 6190 1810 6242 1822
rect 7646 1810 7698 1822
rect 7982 1874 8034 1886
rect 7982 1810 8034 1822
rect 8766 1874 8818 1886
rect 8766 1810 8818 1822
rect 9438 1874 9490 1886
rect 9438 1810 9490 1822
rect 9774 1874 9826 1886
rect 9774 1810 9826 1822
rect 10222 1874 10274 1886
rect 10222 1810 10274 1822
rect 10894 1874 10946 1886
rect 10894 1810 10946 1822
rect 11902 1874 11954 1886
rect 11902 1810 11954 1822
rect 12574 1874 12626 1886
rect 17838 1874 17890 1886
rect 13682 1822 13694 1874
rect 13746 1822 13758 1874
rect 14914 1822 14926 1874
rect 14978 1822 14990 1874
rect 12574 1810 12626 1822
rect 17838 1810 17890 1822
rect 18398 1874 18450 1886
rect 18398 1810 18450 1822
rect 18734 1874 18786 1886
rect 18734 1810 18786 1822
rect 19182 1874 19234 1886
rect 19182 1810 19234 1822
rect 19518 1874 19570 1886
rect 19518 1810 19570 1822
rect 19854 1874 19906 1886
rect 19854 1810 19906 1822
rect 20190 1874 20242 1886
rect 20190 1810 20242 1822
rect 21422 1874 21474 1886
rect 21422 1810 21474 1822
rect 22318 1874 22370 1886
rect 22318 1810 22370 1822
rect 23214 1874 23266 1886
rect 23214 1810 23266 1822
rect 24558 1874 24610 1886
rect 24558 1810 24610 1822
rect 24894 1874 24946 1886
rect 24894 1810 24946 1822
rect 25230 1874 25282 1886
rect 25230 1810 25282 1822
rect 25566 1874 25618 1886
rect 25566 1810 25618 1822
rect 26238 1874 26290 1886
rect 26238 1810 26290 1822
rect 26574 1874 26626 1886
rect 26574 1810 26626 1822
rect 27358 1874 27410 1886
rect 27358 1810 27410 1822
rect 28366 1874 28418 1886
rect 28366 1810 28418 1822
rect 28702 1874 28754 1886
rect 28702 1810 28754 1822
rect 30046 1874 30098 1886
rect 30046 1810 30098 1822
rect 30382 1874 30434 1886
rect 30382 1810 30434 1822
rect 30942 1874 30994 1886
rect 30942 1810 30994 1822
rect 31278 1874 31330 1886
rect 31278 1810 31330 1822
rect 32510 1874 32562 1886
rect 32510 1810 32562 1822
rect 32846 1874 32898 1886
rect 32846 1810 32898 1822
rect 33182 1874 33234 1886
rect 33182 1810 33234 1822
rect 34526 1874 34578 1886
rect 34526 1810 34578 1822
rect 35982 1874 36034 1886
rect 35982 1810 36034 1822
rect 36654 1874 36706 1886
rect 36654 1810 36706 1822
rect 3390 1762 3442 1774
rect 3390 1698 3442 1710
rect 5070 1762 5122 1774
rect 5070 1698 5122 1710
rect 6750 1762 6802 1774
rect 6750 1698 6802 1710
rect 17278 1762 17330 1774
rect 17278 1698 17330 1710
rect 26910 1762 26962 1774
rect 26910 1698 26962 1710
rect 29150 1762 29202 1774
rect 29150 1698 29202 1710
rect 33966 1762 34018 1774
rect 33966 1698 34018 1710
rect 37438 1762 37490 1774
rect 37438 1698 37490 1710
rect 1344 1594 38640 1628
rect 1344 1542 19838 1594
rect 19890 1542 19942 1594
rect 19994 1542 20046 1594
rect 20098 1542 38640 1594
rect 1344 1508 38640 1542
<< via1 >>
rect 4478 97974 4530 98026
rect 4582 97974 4634 98026
rect 4686 97974 4738 98026
rect 35198 97974 35250 98026
rect 35302 97974 35354 98026
rect 35406 97974 35458 98026
rect 14478 97582 14530 97634
rect 15262 97582 15314 97634
rect 13022 97470 13074 97522
rect 1710 97358 1762 97410
rect 4062 97358 4114 97410
rect 6526 97358 6578 97410
rect 9326 97358 9378 97410
rect 11454 97358 11506 97410
rect 15710 97358 15762 97410
rect 16270 97358 16322 97410
rect 16942 97358 16994 97410
rect 18846 97358 18898 97410
rect 19838 97190 19890 97242
rect 19942 97190 19994 97242
rect 20046 97190 20098 97242
rect 7982 96798 8034 96850
rect 8878 96798 8930 96850
rect 13918 96798 13970 96850
rect 14702 96798 14754 96850
rect 31278 96798 31330 96850
rect 32286 96798 32338 96850
rect 34302 96798 34354 96850
rect 35198 96798 35250 96850
rect 9662 96686 9714 96738
rect 10110 96686 10162 96738
rect 12350 96686 12402 96738
rect 15150 96686 15202 96738
rect 6862 96574 6914 96626
rect 30158 96574 30210 96626
rect 33182 96574 33234 96626
rect 4478 96406 4530 96458
rect 4582 96406 4634 96458
rect 4686 96406 4738 96458
rect 35198 96406 35250 96458
rect 35302 96406 35354 96458
rect 35406 96406 35458 96458
rect 15598 96238 15650 96290
rect 19518 96238 19570 96290
rect 23438 96238 23490 96290
rect 16158 96126 16210 96178
rect 2942 96014 2994 96066
rect 3838 96014 3890 96066
rect 6750 96014 6802 96066
rect 7646 96014 7698 96066
rect 9326 96014 9378 96066
rect 10334 96014 10386 96066
rect 13582 96014 13634 96066
rect 14478 96014 14530 96066
rect 17502 96014 17554 96066
rect 18398 96014 18450 96066
rect 21422 96014 21474 96066
rect 22318 96014 22370 96066
rect 29262 96014 29314 96066
rect 30158 96014 30210 96066
rect 32958 96014 33010 96066
rect 33854 96014 33906 96066
rect 8654 95902 8706 95954
rect 24222 95902 24274 95954
rect 25006 95902 25058 95954
rect 25342 95902 25394 95954
rect 26462 95902 26514 95954
rect 26798 95902 26850 95954
rect 5182 95790 5234 95842
rect 5742 95790 5794 95842
rect 11678 95790 11730 95842
rect 12014 95790 12066 95842
rect 20078 95790 20130 95842
rect 20750 95790 20802 95842
rect 23886 95790 23938 95842
rect 25678 95790 25730 95842
rect 26014 95790 26066 95842
rect 27358 95790 27410 95842
rect 31502 95790 31554 95842
rect 35198 95790 35250 95842
rect 19838 95622 19890 95674
rect 19942 95622 19994 95674
rect 20046 95622 20098 95674
rect 6190 95454 6242 95506
rect 9662 95454 9714 95506
rect 12350 95454 12402 95506
rect 15150 95454 15202 95506
rect 16830 95342 16882 95394
rect 3950 95230 4002 95282
rect 4846 95230 4898 95282
rect 6750 95230 6802 95282
rect 7646 95230 7698 95282
rect 13918 95230 13970 95282
rect 14702 95230 14754 95282
rect 16494 95230 16546 95282
rect 17502 95230 17554 95282
rect 18398 95230 18450 95282
rect 21198 95230 21250 95282
rect 22206 95230 22258 95282
rect 24670 95230 24722 95282
rect 25342 95230 25394 95282
rect 26014 95230 26066 95282
rect 28254 95230 28306 95282
rect 29150 95230 29202 95282
rect 33070 95230 33122 95282
rect 34078 95230 34130 95282
rect 35646 95230 35698 95282
rect 36430 95230 36482 95282
rect 9102 95118 9154 95170
rect 19854 95118 19906 95170
rect 23550 95118 23602 95170
rect 30494 95118 30546 95170
rect 19518 95006 19570 95058
rect 27358 95006 27410 95058
rect 35198 95006 35250 95058
rect 37774 95006 37826 95058
rect 4478 94838 4530 94890
rect 4582 94838 4634 94890
rect 4686 94838 4738 94890
rect 35198 94838 35250 94890
rect 35302 94838 35354 94890
rect 35406 94838 35458 94890
rect 4958 94670 5010 94722
rect 20638 94670 20690 94722
rect 25342 94670 25394 94722
rect 34974 94670 35026 94722
rect 5742 94558 5794 94610
rect 6302 94558 6354 94610
rect 15598 94558 15650 94610
rect 15934 94558 15986 94610
rect 22206 94558 22258 94610
rect 26238 94558 26290 94610
rect 2942 94446 2994 94498
rect 3838 94446 3890 94498
rect 16158 94446 16210 94498
rect 16718 94446 16770 94498
rect 18510 94446 18562 94498
rect 19294 94446 19346 94498
rect 21534 94446 21586 94498
rect 22318 94446 22370 94498
rect 22654 94446 22706 94498
rect 25006 94446 25058 94498
rect 25342 94446 25394 94498
rect 25678 94446 25730 94498
rect 27806 94446 27858 94498
rect 28590 94446 28642 94498
rect 29262 94446 29314 94498
rect 30158 94446 30210 94498
rect 32846 94446 32898 94498
rect 33854 94446 33906 94498
rect 1710 94334 1762 94386
rect 16830 94334 16882 94386
rect 21982 94334 22034 94386
rect 22766 94334 22818 94386
rect 24334 94334 24386 94386
rect 25790 94334 25842 94386
rect 17278 94222 17330 94274
rect 17726 94222 17778 94274
rect 21310 94222 21362 94274
rect 23214 94222 23266 94274
rect 24110 94222 24162 94274
rect 24670 94222 24722 94274
rect 31502 94222 31554 94274
rect 19838 94054 19890 94106
rect 19942 94054 19994 94106
rect 20046 94054 20098 94106
rect 4622 93886 4674 93938
rect 9102 93886 9154 93938
rect 16270 93886 16322 93938
rect 20638 93886 20690 93938
rect 23326 93886 23378 93938
rect 13246 93774 13298 93826
rect 3390 93662 3442 93714
rect 4174 93662 4226 93714
rect 6750 93662 6802 93714
rect 7646 93662 7698 93714
rect 12014 93662 12066 93714
rect 13358 93662 13410 93714
rect 16606 93662 16658 93714
rect 16830 93662 16882 93714
rect 17502 93662 17554 93714
rect 18398 93662 18450 93714
rect 20302 93662 20354 93714
rect 20974 93662 21026 93714
rect 21982 93662 22034 93714
rect 23886 93662 23938 93714
rect 25230 93662 25282 93714
rect 26014 93662 26066 93714
rect 28814 93662 28866 93714
rect 29598 93662 29650 93714
rect 33182 93662 33234 93714
rect 33854 93662 33906 93714
rect 9662 93550 9714 93602
rect 12686 93550 12738 93602
rect 20078 93550 20130 93602
rect 23998 93550 24050 93602
rect 24558 93550 24610 93602
rect 2046 93438 2098 93490
rect 12350 93438 12402 93490
rect 19518 93438 19570 93490
rect 27358 93438 27410 93490
rect 30830 93438 30882 93490
rect 35198 93438 35250 93490
rect 4478 93270 4530 93322
rect 4582 93270 4634 93322
rect 4686 93270 4738 93322
rect 35198 93270 35250 93322
rect 35302 93270 35354 93322
rect 35406 93270 35458 93322
rect 4958 93102 5010 93154
rect 10782 93102 10834 93154
rect 19294 93102 19346 93154
rect 23438 93102 23490 93154
rect 24110 93102 24162 93154
rect 24446 93102 24498 93154
rect 25678 93102 25730 93154
rect 5742 92990 5794 93042
rect 9326 92990 9378 93042
rect 17278 92990 17330 93042
rect 18622 92990 18674 93042
rect 20750 92990 20802 93042
rect 31502 92990 31554 93042
rect 2942 92878 2994 92930
rect 3838 92878 3890 92930
rect 6974 92878 7026 92930
rect 7758 92878 7810 92930
rect 12126 92878 12178 92930
rect 12910 92878 12962 92930
rect 17054 92878 17106 92930
rect 17950 92878 18002 92930
rect 21310 92878 21362 92930
rect 22318 92878 22370 92930
rect 24670 92878 24722 92930
rect 29262 92878 29314 92930
rect 30158 92878 30210 92930
rect 31838 92878 31890 92930
rect 32734 92878 32786 92930
rect 9662 92766 9714 92818
rect 10334 92766 10386 92818
rect 13470 92766 13522 92818
rect 13806 92766 13858 92818
rect 14142 92766 14194 92818
rect 14590 92766 14642 92818
rect 19406 92766 19458 92818
rect 25566 92766 25618 92818
rect 26686 92766 26738 92818
rect 27470 92766 27522 92818
rect 25118 92654 25170 92706
rect 26126 92654 26178 92706
rect 34078 92654 34130 92706
rect 19838 92486 19890 92538
rect 19942 92486 19994 92538
rect 20046 92486 20098 92538
rect 5630 92318 5682 92370
rect 8766 92318 8818 92370
rect 10782 92318 10834 92370
rect 23214 92318 23266 92370
rect 4846 92206 4898 92258
rect 9998 92206 10050 92258
rect 10222 92206 10274 92258
rect 13470 92206 13522 92258
rect 14702 92206 14754 92258
rect 15150 92206 15202 92258
rect 20750 92206 20802 92258
rect 26126 92206 26178 92258
rect 37886 92206 37938 92258
rect 2942 92094 2994 92146
rect 3838 92094 3890 92146
rect 6526 92094 6578 92146
rect 7310 92094 7362 92146
rect 10894 92094 10946 92146
rect 12350 92094 12402 92146
rect 12686 92094 12738 92146
rect 14366 92094 14418 92146
rect 20974 92094 21026 92146
rect 21646 92094 21698 92146
rect 25342 92094 25394 92146
rect 27358 92094 27410 92146
rect 33182 92094 33234 92146
rect 33854 92094 33906 92146
rect 38222 92094 38274 92146
rect 22318 91982 22370 92034
rect 23326 91982 23378 92034
rect 24222 91982 24274 92034
rect 24670 91982 24722 92034
rect 26126 91982 26178 92034
rect 27806 91982 27858 92034
rect 37662 91982 37714 92034
rect 10334 91870 10386 91922
rect 14590 91870 14642 91922
rect 35198 91870 35250 91922
rect 4478 91702 4530 91754
rect 4582 91702 4634 91754
rect 4686 91702 4738 91754
rect 35198 91702 35250 91754
rect 35302 91702 35354 91754
rect 35406 91702 35458 91754
rect 4958 91534 5010 91586
rect 12238 91534 12290 91586
rect 12574 91534 12626 91586
rect 14030 91534 14082 91586
rect 14590 91534 14642 91586
rect 32510 91534 32562 91586
rect 8878 91422 8930 91474
rect 14254 91422 14306 91474
rect 14702 91422 14754 91474
rect 2942 91310 2994 91362
rect 3838 91310 3890 91362
rect 11566 91310 11618 91362
rect 12014 91310 12066 91362
rect 13582 91310 13634 91362
rect 13806 91310 13858 91362
rect 27694 91310 27746 91362
rect 33854 91310 33906 91362
rect 34526 91310 34578 91362
rect 13470 91198 13522 91250
rect 23774 91198 23826 91250
rect 5742 91086 5794 91138
rect 11678 91086 11730 91138
rect 19838 90918 19890 90970
rect 19942 90918 19994 90970
rect 20046 90918 20098 90970
rect 12574 90750 12626 90802
rect 24110 90638 24162 90690
rect 26014 90638 26066 90690
rect 29710 90638 29762 90690
rect 30158 90638 30210 90690
rect 3166 90526 3218 90578
rect 3838 90526 3890 90578
rect 12350 90526 12402 90578
rect 22990 90526 23042 90578
rect 25678 90526 25730 90578
rect 30270 90526 30322 90578
rect 5742 90414 5794 90466
rect 21758 90414 21810 90466
rect 22206 90414 22258 90466
rect 22654 90414 22706 90466
rect 23550 90414 23602 90466
rect 24782 90414 24834 90466
rect 25454 90414 25506 90466
rect 26574 90414 26626 90466
rect 27022 90414 27074 90466
rect 27470 90414 27522 90466
rect 27918 90414 27970 90466
rect 28254 90414 28306 90466
rect 5182 90302 5234 90354
rect 12686 90302 12738 90354
rect 26238 90302 26290 90354
rect 26574 90302 26626 90354
rect 30158 90302 30210 90354
rect 4478 90134 4530 90186
rect 4582 90134 4634 90186
rect 4686 90134 4738 90186
rect 35198 90134 35250 90186
rect 35302 90134 35354 90186
rect 35406 90134 35458 90186
rect 30270 89966 30322 90018
rect 10782 89854 10834 89906
rect 21646 89854 21698 89906
rect 27358 89854 27410 89906
rect 30494 89854 30546 89906
rect 3390 89742 3442 89794
rect 4286 89742 4338 89794
rect 7310 89742 7362 89794
rect 7982 89742 8034 89794
rect 8430 89742 8482 89794
rect 9326 89742 9378 89794
rect 19966 89742 20018 89794
rect 22766 89742 22818 89794
rect 27022 89742 27074 89794
rect 30382 89742 30434 89794
rect 22094 89630 22146 89682
rect 23886 89630 23938 89682
rect 26574 89630 26626 89682
rect 2046 89518 2098 89570
rect 4846 89518 4898 89570
rect 5742 89518 5794 89570
rect 15934 89518 15986 89570
rect 16494 89518 16546 89570
rect 17278 89518 17330 89570
rect 19518 89518 19570 89570
rect 22542 89518 22594 89570
rect 22654 89518 22706 89570
rect 22990 89518 23042 89570
rect 23326 89518 23378 89570
rect 23438 89518 23490 89570
rect 23662 89518 23714 89570
rect 24222 89518 24274 89570
rect 24558 89518 24610 89570
rect 25118 89518 25170 89570
rect 25790 89518 25842 89570
rect 26014 89518 26066 89570
rect 26126 89518 26178 89570
rect 26238 89518 26290 89570
rect 28030 89518 28082 89570
rect 28478 89518 28530 89570
rect 29262 89518 29314 89570
rect 19838 89350 19890 89402
rect 19942 89350 19994 89402
rect 20046 89350 20098 89402
rect 24670 89182 24722 89234
rect 16718 89070 16770 89122
rect 6862 88958 6914 89010
rect 7534 88958 7586 89010
rect 12910 88958 12962 89010
rect 13358 88958 13410 89010
rect 16830 88958 16882 89010
rect 17502 88958 17554 89010
rect 20750 88958 20802 89010
rect 21982 88958 22034 89010
rect 23550 88958 23602 89010
rect 23998 88958 24050 89010
rect 24446 88958 24498 89010
rect 25230 88958 25282 89010
rect 37886 88958 37938 89010
rect 9102 88846 9154 88898
rect 14030 88846 14082 88898
rect 16158 88846 16210 88898
rect 18286 88846 18338 88898
rect 20414 88846 20466 88898
rect 21198 88846 21250 88898
rect 22766 88846 22818 88898
rect 24558 88846 24610 88898
rect 30158 88846 30210 88898
rect 31054 88846 31106 88898
rect 36542 88846 36594 88898
rect 16718 88734 16770 88786
rect 4478 88566 4530 88618
rect 4582 88566 4634 88618
rect 4686 88566 4738 88618
rect 35198 88566 35250 88618
rect 35302 88566 35354 88618
rect 35406 88566 35458 88618
rect 2158 88398 2210 88450
rect 21758 88398 21810 88450
rect 22094 88398 22146 88450
rect 25006 88398 25058 88450
rect 12798 88286 12850 88338
rect 15486 88286 15538 88338
rect 16942 88286 16994 88338
rect 24894 88286 24946 88338
rect 29934 88286 29986 88338
rect 32062 88286 32114 88338
rect 3278 88174 3330 88226
rect 4286 88174 4338 88226
rect 7086 88174 7138 88226
rect 7870 88174 7922 88226
rect 9662 88174 9714 88226
rect 10558 88174 10610 88226
rect 12574 88174 12626 88226
rect 14030 88174 14082 88226
rect 15262 88174 15314 88226
rect 16158 88174 16210 88226
rect 19518 88174 19570 88226
rect 19854 88174 19906 88226
rect 20638 88174 20690 88226
rect 21534 88174 21586 88226
rect 22430 88174 22482 88226
rect 24782 88174 24834 88226
rect 28590 88174 28642 88226
rect 29262 88174 29314 88226
rect 14366 88062 14418 88114
rect 14702 88062 14754 88114
rect 27806 88062 27858 88114
rect 35646 88062 35698 88114
rect 4734 87950 4786 88002
rect 9438 87950 9490 88002
rect 12014 87950 12066 88002
rect 12238 87950 12290 88002
rect 13806 87950 13858 88002
rect 14254 87950 14306 88002
rect 19182 87950 19234 88002
rect 19742 87950 19794 88002
rect 20302 87950 20354 88002
rect 20750 87950 20802 88002
rect 25566 87950 25618 88002
rect 32510 87950 32562 88002
rect 35086 87950 35138 88002
rect 35310 87950 35362 88002
rect 35534 87950 35586 88002
rect 19838 87782 19890 87834
rect 19942 87782 19994 87834
rect 20046 87782 20098 87834
rect 9102 87614 9154 87666
rect 11902 87614 11954 87666
rect 14366 87614 14418 87666
rect 15262 87614 15314 87666
rect 15710 87614 15762 87666
rect 17502 87614 17554 87666
rect 20078 87614 20130 87666
rect 22766 87614 22818 87666
rect 22990 87614 23042 87666
rect 23214 87614 23266 87666
rect 23550 87614 23602 87666
rect 23774 87614 23826 87666
rect 13582 87502 13634 87554
rect 16718 87502 16770 87554
rect 18174 87502 18226 87554
rect 18734 87502 18786 87554
rect 19070 87502 19122 87554
rect 21086 87502 21138 87554
rect 24334 87502 24386 87554
rect 24558 87502 24610 87554
rect 27246 87502 27298 87554
rect 31166 87502 31218 87554
rect 35646 87502 35698 87554
rect 3278 87390 3330 87442
rect 4286 87390 4338 87442
rect 6862 87390 6914 87442
rect 7758 87390 7810 87442
rect 9662 87390 9714 87442
rect 10558 87390 10610 87442
rect 12350 87390 12402 87442
rect 13022 87390 13074 87442
rect 13918 87390 13970 87442
rect 15598 87390 15650 87442
rect 16270 87390 16322 87442
rect 17838 87390 17890 87442
rect 19630 87390 19682 87442
rect 20638 87390 20690 87442
rect 20974 87390 21026 87442
rect 21198 87390 21250 87442
rect 22206 87390 22258 87442
rect 24222 87390 24274 87442
rect 24670 87390 24722 87442
rect 25678 87390 25730 87442
rect 30830 87390 30882 87442
rect 31054 87390 31106 87442
rect 32062 87390 32114 87442
rect 32958 87390 33010 87442
rect 33406 87390 33458 87442
rect 33630 87390 33682 87442
rect 34526 87390 34578 87442
rect 34862 87390 34914 87442
rect 4734 87278 4786 87330
rect 5182 87278 5234 87330
rect 23102 87278 23154 87330
rect 23662 87278 23714 87330
rect 32510 87278 32562 87330
rect 33518 87278 33570 87330
rect 37774 87278 37826 87330
rect 2158 87166 2210 87218
rect 12574 87166 12626 87218
rect 15710 87166 15762 87218
rect 31614 87166 31666 87218
rect 4478 86998 4530 87050
rect 4582 86998 4634 87050
rect 4686 86998 4738 87050
rect 35198 86998 35250 87050
rect 35302 86998 35354 87050
rect 35406 86998 35458 87050
rect 2158 86830 2210 86882
rect 24670 86830 24722 86882
rect 26014 86830 26066 86882
rect 16046 86718 16098 86770
rect 16830 86718 16882 86770
rect 18286 86718 18338 86770
rect 19182 86718 19234 86770
rect 19854 86718 19906 86770
rect 22094 86718 22146 86770
rect 22318 86718 22370 86770
rect 26126 86718 26178 86770
rect 29150 86718 29202 86770
rect 29598 86718 29650 86770
rect 32846 86718 32898 86770
rect 34974 86718 35026 86770
rect 36206 86718 36258 86770
rect 3278 86606 3330 86658
rect 4286 86606 4338 86658
rect 8430 86606 8482 86658
rect 9326 86606 9378 86658
rect 10110 86606 10162 86658
rect 10670 86606 10722 86658
rect 11678 86606 11730 86658
rect 16942 86606 16994 86658
rect 17502 86606 17554 86658
rect 20302 86606 20354 86658
rect 20750 86606 20802 86658
rect 21982 86606 22034 86658
rect 22766 86606 22818 86658
rect 23214 86606 23266 86658
rect 23550 86606 23602 86658
rect 24334 86606 24386 86658
rect 25118 86606 25170 86658
rect 25902 86606 25954 86658
rect 27134 86606 27186 86658
rect 28030 86606 28082 86658
rect 28478 86606 28530 86658
rect 32510 86606 32562 86658
rect 35646 86606 35698 86658
rect 10894 86494 10946 86546
rect 12574 86494 12626 86546
rect 20414 86494 20466 86546
rect 23774 86494 23826 86546
rect 24110 86494 24162 86546
rect 26910 86494 26962 86546
rect 31726 86494 31778 86546
rect 4734 86382 4786 86434
rect 6974 86382 7026 86434
rect 20638 86382 20690 86434
rect 23662 86382 23714 86434
rect 27022 86382 27074 86434
rect 27358 86382 27410 86434
rect 27806 86382 27858 86434
rect 27918 86382 27970 86434
rect 29262 86382 29314 86434
rect 19838 86214 19890 86266
rect 19942 86214 19994 86266
rect 20046 86214 20098 86266
rect 7310 86046 7362 86098
rect 11678 86046 11730 86098
rect 12126 86046 12178 86098
rect 31502 86046 31554 86098
rect 36318 86046 36370 86098
rect 11566 85934 11618 85986
rect 25342 85934 25394 85986
rect 27470 85934 27522 85986
rect 31614 85934 31666 85986
rect 3278 85822 3330 85874
rect 4286 85822 4338 85874
rect 4622 85822 4674 85874
rect 5406 85822 5458 85874
rect 6974 85822 7026 85874
rect 14142 85822 14194 85874
rect 23550 85822 23602 85874
rect 25230 85822 25282 85874
rect 30270 85822 30322 85874
rect 31166 85822 31218 85874
rect 31838 85822 31890 85874
rect 33630 85822 33682 85874
rect 34974 85822 35026 85874
rect 36206 85822 36258 85874
rect 13806 85710 13858 85762
rect 14254 85710 14306 85762
rect 19630 85710 19682 85762
rect 32510 85710 32562 85762
rect 33070 85710 33122 85762
rect 35086 85710 35138 85762
rect 35758 85710 35810 85762
rect 36878 85710 36930 85762
rect 37326 85710 37378 85762
rect 2158 85598 2210 85650
rect 14478 85598 14530 85650
rect 33294 85598 33346 85650
rect 36318 85598 36370 85650
rect 4478 85430 4530 85482
rect 4582 85430 4634 85482
rect 4686 85430 4738 85482
rect 35198 85430 35250 85482
rect 35302 85430 35354 85482
rect 35406 85430 35458 85482
rect 2158 85262 2210 85314
rect 14814 85262 14866 85314
rect 15150 85262 15202 85314
rect 19070 85262 19122 85314
rect 19630 85262 19682 85314
rect 20414 85262 20466 85314
rect 21758 85262 21810 85314
rect 32510 85262 32562 85314
rect 32846 85262 32898 85314
rect 29486 85150 29538 85202
rect 29934 85150 29986 85202
rect 30830 85150 30882 85202
rect 31726 85150 31778 85202
rect 37102 85150 37154 85202
rect 3278 85038 3330 85090
rect 4286 85038 4338 85090
rect 14030 85038 14082 85090
rect 14254 85038 14306 85090
rect 14590 85038 14642 85090
rect 15598 85038 15650 85090
rect 19182 85038 19234 85090
rect 20526 85038 20578 85090
rect 20750 85038 20802 85090
rect 21422 85038 21474 85090
rect 21870 85038 21922 85090
rect 22094 85038 22146 85090
rect 22318 85038 22370 85090
rect 22654 85038 22706 85090
rect 29374 85038 29426 85090
rect 31278 85038 31330 85090
rect 31614 85038 31666 85090
rect 31838 85038 31890 85090
rect 34414 85038 34466 85090
rect 35646 85038 35698 85090
rect 35870 85038 35922 85090
rect 25566 84926 25618 84978
rect 32062 84926 32114 84978
rect 34974 84926 35026 84978
rect 35310 84926 35362 84978
rect 35982 84926 36034 84978
rect 4734 84814 4786 84866
rect 12910 84814 12962 84866
rect 13806 84814 13858 84866
rect 14142 84814 14194 84866
rect 18734 84814 18786 84866
rect 19742 84814 19794 84866
rect 20078 84814 20130 84866
rect 28366 84814 28418 84866
rect 30382 84814 30434 84866
rect 32734 84814 32786 84866
rect 33966 84814 34018 84866
rect 34526 84814 34578 84866
rect 34750 84814 34802 84866
rect 35086 84814 35138 84866
rect 35422 84814 35474 84866
rect 36206 84814 36258 84866
rect 37662 84814 37714 84866
rect 19838 84646 19890 84698
rect 19942 84646 19994 84698
rect 20046 84646 20098 84698
rect 17614 84478 17666 84530
rect 18846 84478 18898 84530
rect 19070 84478 19122 84530
rect 21086 84478 21138 84530
rect 21310 84478 21362 84530
rect 23886 84478 23938 84530
rect 25678 84478 25730 84530
rect 25902 84478 25954 84530
rect 28590 84478 28642 84530
rect 29150 84478 29202 84530
rect 30158 84478 30210 84530
rect 30606 84478 30658 84530
rect 31054 84478 31106 84530
rect 34190 84478 34242 84530
rect 34974 84478 35026 84530
rect 14702 84366 14754 84418
rect 19966 84366 20018 84418
rect 20414 84366 20466 84418
rect 23326 84366 23378 84418
rect 24222 84366 24274 84418
rect 28030 84366 28082 84418
rect 29710 84366 29762 84418
rect 3278 84254 3330 84306
rect 4286 84254 4338 84306
rect 15486 84254 15538 84306
rect 18510 84254 18562 84306
rect 19406 84254 19458 84306
rect 20190 84254 20242 84306
rect 20638 84254 20690 84306
rect 22318 84254 22370 84306
rect 22990 84254 23042 84306
rect 23438 84254 23490 84306
rect 24446 84254 24498 84306
rect 25230 84254 25282 84306
rect 26910 84254 26962 84306
rect 27806 84254 27858 84306
rect 35310 84254 35362 84306
rect 4734 84142 4786 84194
rect 8766 84142 8818 84194
rect 12574 84142 12626 84194
rect 15934 84142 15986 84194
rect 18062 84142 18114 84194
rect 21198 84142 21250 84194
rect 22094 84142 22146 84194
rect 22878 84142 22930 84194
rect 25454 84142 25506 84194
rect 25790 84142 25842 84194
rect 27134 84142 27186 84194
rect 27470 84142 27522 84194
rect 33854 84142 33906 84194
rect 36094 84142 36146 84194
rect 38222 84142 38274 84194
rect 2158 84030 2210 84082
rect 18734 84030 18786 84082
rect 19854 84030 19906 84082
rect 28254 84030 28306 84082
rect 4478 83862 4530 83914
rect 4582 83862 4634 83914
rect 4686 83862 4738 83914
rect 35198 83862 35250 83914
rect 35302 83862 35354 83914
rect 35406 83862 35458 83914
rect 2158 83694 2210 83746
rect 9102 83694 9154 83746
rect 9774 83694 9826 83746
rect 14814 83694 14866 83746
rect 29262 83694 29314 83746
rect 37102 83694 37154 83746
rect 9774 83582 9826 83634
rect 16158 83582 16210 83634
rect 17726 83582 17778 83634
rect 19294 83582 19346 83634
rect 20414 83582 20466 83634
rect 30494 83582 30546 83634
rect 34750 83582 34802 83634
rect 37662 83582 37714 83634
rect 38110 83582 38162 83634
rect 3278 83470 3330 83522
rect 4286 83470 4338 83522
rect 8094 83470 8146 83522
rect 15374 83470 15426 83522
rect 17838 83470 17890 83522
rect 18398 83470 18450 83522
rect 18510 83470 18562 83522
rect 19182 83470 19234 83522
rect 19966 83470 20018 83522
rect 21870 83470 21922 83522
rect 24782 83470 24834 83522
rect 29038 83470 29090 83522
rect 34862 83470 34914 83522
rect 35646 83470 35698 83522
rect 35982 83470 36034 83522
rect 4734 83358 4786 83410
rect 8430 83358 8482 83410
rect 14142 83358 14194 83410
rect 14254 83358 14306 83410
rect 14366 83358 14418 83410
rect 15598 83358 15650 83410
rect 22878 83358 22930 83410
rect 26014 83358 26066 83410
rect 29598 83358 29650 83410
rect 31390 83358 31442 83410
rect 36206 83358 36258 83410
rect 36990 83358 37042 83410
rect 37102 83358 37154 83410
rect 8318 83246 8370 83298
rect 9326 83246 9378 83298
rect 13022 83246 13074 83298
rect 13694 83246 13746 83298
rect 15150 83246 15202 83298
rect 15262 83246 15314 83298
rect 16606 83246 16658 83298
rect 17166 83246 17218 83298
rect 18286 83246 18338 83298
rect 19518 83246 19570 83298
rect 22318 83246 22370 83298
rect 29374 83246 29426 83298
rect 30046 83246 30098 83298
rect 30942 83246 30994 83298
rect 34078 83246 34130 83298
rect 34414 83246 34466 83298
rect 34638 83246 34690 83298
rect 37550 83246 37602 83298
rect 19838 83078 19890 83130
rect 19942 83078 19994 83130
rect 20046 83078 20098 83130
rect 17614 82910 17666 82962
rect 28254 82910 28306 82962
rect 29038 82910 29090 82962
rect 30606 82910 30658 82962
rect 8206 82798 8258 82850
rect 10222 82798 10274 82850
rect 12686 82798 12738 82850
rect 18622 82798 18674 82850
rect 26462 82798 26514 82850
rect 28366 82798 28418 82850
rect 35758 82798 35810 82850
rect 8990 82686 9042 82738
rect 9550 82686 9602 82738
rect 9774 82686 9826 82738
rect 9998 82686 10050 82738
rect 12014 82686 12066 82738
rect 19630 82686 19682 82738
rect 25230 82686 25282 82738
rect 25902 82686 25954 82738
rect 27246 82686 27298 82738
rect 27918 82686 27970 82738
rect 28590 82686 28642 82738
rect 28814 82686 28866 82738
rect 29150 82686 29202 82738
rect 29374 82686 29426 82738
rect 34974 82686 35026 82738
rect 6078 82574 6130 82626
rect 9662 82574 9714 82626
rect 10670 82574 10722 82626
rect 11118 82574 11170 82626
rect 14814 82574 14866 82626
rect 15486 82574 15538 82626
rect 18174 82574 18226 82626
rect 23550 82574 23602 82626
rect 26238 82574 26290 82626
rect 27134 82574 27186 82626
rect 29822 82574 29874 82626
rect 30158 82574 30210 82626
rect 31166 82574 31218 82626
rect 31614 82574 31666 82626
rect 33182 82574 33234 82626
rect 34638 82574 34690 82626
rect 37886 82574 37938 82626
rect 18510 82462 18562 82514
rect 18846 82462 18898 82514
rect 27022 82462 27074 82514
rect 31390 82462 31442 82514
rect 31838 82462 31890 82514
rect 32286 82462 32338 82514
rect 4478 82294 4530 82346
rect 4582 82294 4634 82346
rect 4686 82294 4738 82346
rect 35198 82294 35250 82346
rect 35302 82294 35354 82346
rect 35406 82294 35458 82346
rect 14478 82126 14530 82178
rect 14926 82126 14978 82178
rect 15374 82126 15426 82178
rect 27358 82126 27410 82178
rect 11566 82014 11618 82066
rect 15262 82014 15314 82066
rect 18174 82014 18226 82066
rect 20302 82014 20354 82066
rect 23438 82014 23490 82066
rect 27022 82014 27074 82066
rect 5182 81902 5234 81954
rect 6302 81902 6354 81954
rect 6638 81902 6690 81954
rect 10446 81902 10498 81954
rect 13694 81902 13746 81954
rect 17390 81902 17442 81954
rect 25566 81902 25618 81954
rect 27470 81902 27522 81954
rect 27918 81902 27970 81954
rect 28366 81902 28418 81954
rect 28590 81902 28642 81954
rect 29934 81902 29986 81954
rect 30606 81902 30658 81954
rect 31166 81902 31218 81954
rect 32958 81902 33010 81954
rect 35198 81902 35250 81954
rect 36206 81902 36258 81954
rect 4846 81790 4898 81842
rect 6078 81790 6130 81842
rect 9662 81790 9714 81842
rect 10782 81790 10834 81842
rect 10894 81790 10946 81842
rect 11006 81790 11058 81842
rect 14142 81790 14194 81842
rect 14366 81790 14418 81842
rect 26910 81790 26962 81842
rect 27134 81790 27186 81842
rect 30718 81790 30770 81842
rect 32174 81790 32226 81842
rect 4622 81678 4674 81730
rect 4958 81678 5010 81730
rect 5854 81678 5906 81730
rect 6414 81678 6466 81730
rect 7422 81678 7474 81730
rect 13022 81678 13074 81730
rect 14030 81678 14082 81730
rect 14814 81678 14866 81730
rect 17054 81678 17106 81730
rect 28142 81678 28194 81730
rect 29598 81678 29650 81730
rect 31278 81678 31330 81730
rect 34190 81678 34242 81730
rect 35310 81678 35362 81730
rect 19838 81510 19890 81562
rect 19942 81510 19994 81562
rect 20046 81510 20098 81562
rect 7086 81342 7138 81394
rect 9886 81342 9938 81394
rect 14478 81342 14530 81394
rect 16942 81342 16994 81394
rect 26574 81342 26626 81394
rect 27806 81342 27858 81394
rect 31614 81342 31666 81394
rect 5854 81230 5906 81282
rect 10222 81230 10274 81282
rect 18174 81230 18226 81282
rect 20974 81230 21026 81282
rect 21982 81230 22034 81282
rect 25454 81230 25506 81282
rect 27694 81230 27746 81282
rect 28702 81230 28754 81282
rect 31054 81230 31106 81282
rect 6526 81118 6578 81170
rect 9662 81118 9714 81170
rect 9774 81118 9826 81170
rect 9998 81118 10050 81170
rect 13246 81118 13298 81170
rect 13470 81118 13522 81170
rect 17390 81118 17442 81170
rect 20862 81118 20914 81170
rect 21198 81118 21250 81170
rect 21422 81118 21474 81170
rect 22094 81118 22146 81170
rect 22430 81118 22482 81170
rect 22654 81118 22706 81170
rect 23102 81118 23154 81170
rect 24334 81118 24386 81170
rect 24558 81118 24610 81170
rect 25230 81118 25282 81170
rect 25678 81118 25730 81170
rect 25902 81118 25954 81170
rect 26462 81118 26514 81170
rect 27134 81118 27186 81170
rect 27470 81118 27522 81170
rect 27918 81118 27970 81170
rect 28254 81118 28306 81170
rect 28478 81118 28530 81170
rect 28814 81118 28866 81170
rect 29038 81118 29090 81170
rect 30718 81118 30770 81170
rect 3726 81006 3778 81058
rect 8990 81006 9042 81058
rect 10670 81006 10722 81058
rect 12574 81006 12626 81058
rect 14030 81006 14082 81058
rect 16382 81006 16434 81058
rect 20302 81006 20354 81058
rect 20638 81006 20690 81058
rect 25454 81006 25506 81058
rect 26686 81006 26738 81058
rect 21982 80894 22034 80946
rect 23998 80894 24050 80946
rect 26910 80894 26962 80946
rect 29262 81006 29314 81058
rect 29598 80894 29650 80946
rect 29934 80894 29986 80946
rect 30270 80894 30322 80946
rect 4478 80726 4530 80778
rect 4582 80726 4634 80778
rect 4686 80726 4738 80778
rect 35198 80726 35250 80778
rect 35302 80726 35354 80778
rect 35406 80726 35458 80778
rect 17390 80558 17442 80610
rect 19294 80558 19346 80610
rect 20302 80558 20354 80610
rect 29710 80558 29762 80610
rect 17054 80446 17106 80498
rect 27694 80446 27746 80498
rect 29262 80446 29314 80498
rect 16494 80334 16546 80386
rect 19406 80334 19458 80386
rect 20078 80334 20130 80386
rect 20526 80334 20578 80386
rect 20638 80334 20690 80386
rect 21534 80334 21586 80386
rect 22094 80334 22146 80386
rect 28478 80334 28530 80386
rect 30046 80334 30098 80386
rect 30718 80334 30770 80386
rect 11902 80222 11954 80274
rect 17614 80222 17666 80274
rect 18062 80222 18114 80274
rect 25454 80222 25506 80274
rect 27918 80222 27970 80274
rect 28142 80222 28194 80274
rect 30830 80222 30882 80274
rect 11566 80110 11618 80162
rect 16718 80110 16770 80162
rect 20638 80110 20690 80162
rect 21534 80110 21586 80162
rect 28254 80110 28306 80162
rect 19838 79942 19890 79994
rect 19942 79942 19994 79994
rect 20046 79942 20098 79994
rect 15374 79774 15426 79826
rect 17614 79774 17666 79826
rect 6078 79662 6130 79714
rect 11342 79662 11394 79714
rect 17950 79662 18002 79714
rect 23326 79662 23378 79714
rect 31502 79662 31554 79714
rect 31950 79662 32002 79714
rect 5966 79550 6018 79602
rect 6302 79550 6354 79602
rect 10558 79550 10610 79602
rect 14142 79550 14194 79602
rect 18286 79550 18338 79602
rect 18622 79550 18674 79602
rect 19070 79550 19122 79602
rect 22318 79550 22370 79602
rect 22654 79550 22706 79602
rect 23438 79550 23490 79602
rect 23662 79550 23714 79602
rect 23886 79550 23938 79602
rect 25902 79550 25954 79602
rect 5630 79438 5682 79490
rect 6862 79438 6914 79490
rect 7198 79438 7250 79490
rect 9662 79438 9714 79490
rect 13470 79438 13522 79490
rect 16382 79438 16434 79490
rect 16830 79438 16882 79490
rect 18398 79438 18450 79490
rect 22430 79438 22482 79490
rect 24446 79438 24498 79490
rect 27246 79438 27298 79490
rect 33294 79438 33346 79490
rect 21198 79326 21250 79378
rect 21870 79326 21922 79378
rect 24446 79326 24498 79378
rect 24782 79326 24834 79378
rect 30942 79326 30994 79378
rect 31278 79326 31330 79378
rect 4478 79158 4530 79210
rect 4582 79158 4634 79210
rect 4686 79158 4738 79210
rect 35198 79158 35250 79210
rect 35302 79158 35354 79210
rect 35406 79158 35458 79210
rect 11902 78990 11954 79042
rect 10110 78878 10162 78930
rect 12238 78878 12290 78930
rect 19070 78878 19122 78930
rect 25006 78878 25058 78930
rect 25342 78878 25394 78930
rect 25790 78878 25842 78930
rect 27358 78878 27410 78930
rect 28030 78878 28082 78930
rect 29150 78878 29202 78930
rect 29710 78878 29762 78930
rect 30494 78878 30546 78930
rect 31502 78878 31554 78930
rect 32398 78878 32450 78930
rect 33294 78878 33346 78930
rect 33742 78878 33794 78930
rect 6302 78766 6354 78818
rect 7534 78766 7586 78818
rect 10670 78766 10722 78818
rect 11566 78766 11618 78818
rect 12462 78766 12514 78818
rect 14590 78766 14642 78818
rect 14926 78766 14978 78818
rect 15038 78766 15090 78818
rect 16270 78766 16322 78818
rect 20078 78766 20130 78818
rect 20526 78766 20578 78818
rect 23998 78766 24050 78818
rect 24558 78766 24610 78818
rect 26126 78766 26178 78818
rect 27246 78766 27298 78818
rect 27694 78766 27746 78818
rect 28366 78766 28418 78818
rect 29486 78766 29538 78818
rect 30606 78766 30658 78818
rect 31054 78766 31106 78818
rect 31390 78766 31442 78818
rect 31838 78766 31890 78818
rect 5966 78654 6018 78706
rect 6526 78654 6578 78706
rect 8878 78654 8930 78706
rect 16942 78654 16994 78706
rect 20638 78654 20690 78706
rect 23438 78654 23490 78706
rect 24110 78654 24162 78706
rect 24782 78654 24834 78706
rect 25678 78654 25730 78706
rect 26014 78654 26066 78706
rect 27134 78654 27186 78706
rect 28590 78654 28642 78706
rect 31726 78654 31778 78706
rect 34974 78654 35026 78706
rect 6302 78542 6354 78594
rect 10110 78542 10162 78594
rect 10222 78542 10274 78594
rect 10446 78542 10498 78594
rect 11118 78542 11170 78594
rect 14366 78542 14418 78594
rect 14702 78542 14754 78594
rect 15822 78542 15874 78594
rect 19854 78542 19906 78594
rect 20750 78542 20802 78594
rect 21646 78542 21698 78594
rect 21870 78542 21922 78594
rect 21982 78542 22034 78594
rect 22094 78542 22146 78594
rect 22542 78542 22594 78594
rect 22766 78542 22818 78594
rect 22878 78542 22930 78594
rect 22990 78542 23042 78594
rect 24334 78542 24386 78594
rect 27470 78542 27522 78594
rect 30494 78542 30546 78594
rect 30830 78542 30882 78594
rect 32846 78542 32898 78594
rect 34638 78542 34690 78594
rect 34862 78542 34914 78594
rect 35646 78542 35698 78594
rect 35870 78542 35922 78594
rect 35982 78542 36034 78594
rect 36094 78542 36146 78594
rect 19838 78374 19890 78426
rect 19942 78374 19994 78426
rect 20046 78374 20098 78426
rect 6974 78206 7026 78258
rect 17726 78206 17778 78258
rect 18622 78206 18674 78258
rect 27582 78206 27634 78258
rect 29150 78206 29202 78258
rect 29262 78206 29314 78258
rect 29374 78206 29426 78258
rect 30158 78206 30210 78258
rect 31390 78206 31442 78258
rect 32174 78206 32226 78258
rect 33630 78206 33682 78258
rect 35198 78206 35250 78258
rect 35310 78206 35362 78258
rect 9886 78094 9938 78146
rect 14030 78094 14082 78146
rect 17614 78094 17666 78146
rect 20190 78094 20242 78146
rect 26126 78094 26178 78146
rect 34638 78094 34690 78146
rect 37102 78094 37154 78146
rect 6526 77982 6578 78034
rect 9550 77982 9602 78034
rect 13358 77982 13410 78034
rect 17390 77982 17442 78034
rect 17950 77982 18002 78034
rect 23550 77982 23602 78034
rect 25790 77982 25842 78034
rect 26350 77982 26402 78034
rect 26686 77982 26738 78034
rect 28478 77982 28530 78034
rect 29486 77982 29538 78034
rect 29710 77982 29762 78034
rect 30270 77982 30322 78034
rect 30494 77982 30546 78034
rect 30718 77982 30770 78034
rect 31166 77982 31218 78034
rect 31278 77982 31330 78034
rect 31502 77982 31554 78034
rect 31726 77982 31778 78034
rect 35086 77982 35138 78034
rect 35534 77982 35586 78034
rect 35870 77982 35922 78034
rect 36766 77982 36818 78034
rect 37214 77982 37266 78034
rect 3614 77870 3666 77922
rect 5742 77870 5794 77922
rect 8990 77870 9042 77922
rect 12910 77870 12962 77922
rect 16158 77870 16210 77922
rect 16830 77870 16882 77922
rect 24782 77870 24834 77922
rect 26574 77870 26626 77922
rect 27022 77870 27074 77922
rect 28030 77870 28082 77922
rect 30158 77870 30210 77922
rect 33182 77870 33234 77922
rect 34078 77870 34130 77922
rect 36318 77870 36370 77922
rect 9550 77758 9602 77810
rect 25230 77758 25282 77810
rect 25566 77758 25618 77810
rect 27246 77758 27298 77810
rect 34414 77758 34466 77810
rect 34750 77758 34802 77810
rect 36206 77758 36258 77810
rect 36542 77758 36594 77810
rect 4478 77590 4530 77642
rect 4582 77590 4634 77642
rect 4686 77590 4738 77642
rect 35198 77590 35250 77642
rect 35302 77590 35354 77642
rect 35406 77590 35458 77642
rect 35198 77422 35250 77474
rect 35982 77422 36034 77474
rect 37214 77422 37266 77474
rect 37886 77422 37938 77474
rect 7310 77310 7362 77362
rect 9438 77310 9490 77362
rect 12126 77310 12178 77362
rect 13806 77310 13858 77362
rect 15038 77310 15090 77362
rect 21534 77310 21586 77362
rect 28142 77310 28194 77362
rect 35422 77310 35474 77362
rect 35646 77310 35698 77362
rect 37998 77310 38050 77362
rect 10110 77198 10162 77250
rect 10670 77198 10722 77250
rect 12574 77198 12626 77250
rect 12910 77198 12962 77250
rect 14478 77198 14530 77250
rect 20638 77198 20690 77250
rect 25454 77198 25506 77250
rect 26910 77198 26962 77250
rect 27246 77198 27298 77250
rect 27358 77198 27410 77250
rect 29262 77198 29314 77250
rect 31278 77198 31330 77250
rect 32062 77198 32114 77250
rect 32174 77198 32226 77250
rect 32510 77198 32562 77250
rect 33070 77198 33122 77250
rect 34750 77198 34802 77250
rect 35758 77198 35810 77250
rect 36430 77198 36482 77250
rect 37102 77198 37154 77250
rect 37438 77198 37490 77250
rect 12350 77086 12402 77138
rect 13694 77086 13746 77138
rect 14142 77086 14194 77138
rect 15150 77086 15202 77138
rect 16830 77086 16882 77138
rect 28366 77086 28418 77138
rect 31166 77086 31218 77138
rect 31502 77086 31554 77138
rect 31726 77086 31778 77138
rect 32398 77086 32450 77138
rect 33294 77086 33346 77138
rect 33630 77086 33682 77138
rect 34190 77086 34242 77138
rect 34526 77086 34578 77138
rect 36318 77086 36370 77138
rect 38110 77086 38162 77138
rect 12462 76974 12514 77026
rect 13918 76974 13970 77026
rect 14926 76974 14978 77026
rect 27134 76974 27186 77026
rect 27806 76974 27858 77026
rect 29710 76974 29762 77026
rect 30270 76974 30322 77026
rect 30606 76974 30658 77026
rect 33518 76974 33570 77026
rect 34302 76974 34354 77026
rect 37102 76974 37154 77026
rect 19838 76806 19890 76858
rect 19942 76806 19994 76858
rect 20046 76806 20098 76858
rect 15038 76638 15090 76690
rect 15486 76638 15538 76690
rect 15934 76638 15986 76690
rect 16606 76638 16658 76690
rect 16718 76638 16770 76690
rect 16830 76638 16882 76690
rect 24334 76638 24386 76690
rect 25342 76638 25394 76690
rect 26238 76638 26290 76690
rect 27806 76638 27858 76690
rect 31390 76638 31442 76690
rect 33406 76638 33458 76690
rect 36990 76638 37042 76690
rect 37662 76638 37714 76690
rect 8766 76526 8818 76578
rect 12238 76526 12290 76578
rect 17726 76526 17778 76578
rect 20638 76526 20690 76578
rect 26798 76526 26850 76578
rect 27022 76526 27074 76578
rect 27134 76526 27186 76578
rect 27246 76526 27298 76578
rect 28366 76526 28418 76578
rect 30494 76526 30546 76578
rect 31166 76526 31218 76578
rect 31502 76526 31554 76578
rect 32398 76526 32450 76578
rect 32622 76526 32674 76578
rect 35870 76526 35922 76578
rect 36430 76526 36482 76578
rect 36878 76526 36930 76578
rect 37886 76526 37938 76578
rect 9550 76414 9602 76466
rect 9774 76414 9826 76466
rect 9998 76414 10050 76466
rect 10222 76414 10274 76466
rect 11454 76414 11506 76466
rect 16158 76414 16210 76466
rect 17278 76414 17330 76466
rect 17838 76414 17890 76466
rect 18734 76414 18786 76466
rect 25230 76414 25282 76466
rect 25566 76414 25618 76466
rect 25790 76414 25842 76466
rect 27358 76414 27410 76466
rect 27582 76414 27634 76466
rect 27918 76414 27970 76466
rect 29598 76414 29650 76466
rect 30382 76414 30434 76466
rect 31726 76414 31778 76466
rect 32286 76414 32338 76466
rect 33294 76414 33346 76466
rect 33518 76414 33570 76466
rect 33966 76414 34018 76466
rect 35310 76414 35362 76466
rect 35646 76414 35698 76466
rect 37102 76414 37154 76466
rect 37438 76414 37490 76466
rect 37998 76414 38050 76466
rect 8318 76302 8370 76354
rect 8878 76302 8930 76354
rect 9886 76302 9938 76354
rect 10670 76302 10722 76354
rect 11118 76302 11170 76354
rect 14366 76302 14418 76354
rect 17502 76302 17554 76354
rect 29150 76302 29202 76354
rect 34750 76302 34802 76354
rect 8990 76190 9042 76242
rect 28254 76190 28306 76242
rect 29038 76190 29090 76242
rect 29934 76190 29986 76242
rect 34190 76190 34242 76242
rect 34526 76190 34578 76242
rect 4478 76022 4530 76074
rect 4582 76022 4634 76074
rect 4686 76022 4738 76074
rect 35198 76022 35250 76074
rect 35302 76022 35354 76074
rect 35406 76022 35458 76074
rect 19518 75854 19570 75906
rect 32510 75854 32562 75906
rect 33294 75854 33346 75906
rect 34078 75854 34130 75906
rect 6862 75742 6914 75794
rect 7646 75742 7698 75794
rect 9774 75742 9826 75794
rect 11006 75742 11058 75794
rect 20750 75742 20802 75794
rect 22654 75742 22706 75794
rect 26126 75742 26178 75794
rect 29262 75742 29314 75794
rect 30046 75742 30098 75794
rect 31054 75742 31106 75794
rect 32958 75742 33010 75794
rect 35534 75742 35586 75794
rect 37102 75742 37154 75794
rect 5966 75630 6018 75682
rect 6302 75630 6354 75682
rect 6526 75630 6578 75682
rect 10446 75630 10498 75682
rect 14590 75630 14642 75682
rect 15934 75630 15986 75682
rect 16270 75630 16322 75682
rect 21646 75630 21698 75682
rect 24782 75630 24834 75682
rect 30158 75630 30210 75682
rect 30606 75630 30658 75682
rect 31278 75630 31330 75682
rect 31838 75630 31890 75682
rect 31950 75630 32002 75682
rect 34414 75630 34466 75682
rect 34526 75630 34578 75682
rect 35198 75630 35250 75682
rect 35310 75630 35362 75682
rect 36094 75630 36146 75682
rect 36206 75630 36258 75682
rect 6078 75518 6130 75570
rect 30942 75518 30994 75570
rect 31502 75518 31554 75570
rect 32174 75518 32226 75570
rect 32398 75518 32450 75570
rect 33518 75518 33570 75570
rect 33966 75518 34018 75570
rect 34638 75518 34690 75570
rect 34974 75518 35026 75570
rect 35646 75518 35698 75570
rect 36990 75518 37042 75570
rect 37214 75518 37266 75570
rect 7310 75406 7362 75458
rect 15038 75406 15090 75458
rect 30046 75406 30098 75458
rect 30382 75406 30434 75458
rect 33742 75406 33794 75458
rect 35870 75406 35922 75458
rect 37438 75406 37490 75458
rect 19838 75238 19890 75290
rect 19942 75238 19994 75290
rect 20046 75238 20098 75290
rect 17726 75070 17778 75122
rect 24558 75070 24610 75122
rect 25230 75070 25282 75122
rect 27470 75070 27522 75122
rect 31726 75070 31778 75122
rect 32510 75070 32562 75122
rect 33070 75070 33122 75122
rect 33742 75070 33794 75122
rect 33966 75070 34018 75122
rect 35310 75070 35362 75122
rect 36318 75070 36370 75122
rect 36766 75070 36818 75122
rect 8766 74958 8818 75010
rect 23774 74958 23826 75010
rect 24446 74958 24498 75010
rect 26462 74958 26514 75010
rect 27134 74958 27186 75010
rect 29038 74958 29090 75010
rect 33406 74958 33458 75010
rect 34078 74958 34130 75010
rect 35422 74958 35474 75010
rect 36654 74958 36706 75010
rect 37214 74958 37266 75010
rect 7198 74846 7250 74898
rect 7758 74846 7810 74898
rect 7870 74846 7922 74898
rect 8318 74846 8370 74898
rect 11342 74846 11394 74898
rect 17950 74846 18002 74898
rect 18174 74846 18226 74898
rect 18510 74846 18562 74898
rect 19070 74846 19122 74898
rect 22430 74846 22482 74898
rect 22878 74846 22930 74898
rect 22990 74846 23042 74898
rect 23102 74846 23154 74898
rect 23326 74846 23378 74898
rect 23886 74846 23938 74898
rect 24782 74846 24834 74898
rect 25790 74846 25842 74898
rect 26798 74846 26850 74898
rect 27582 74846 27634 74898
rect 28478 74846 28530 74898
rect 29150 74846 29202 74898
rect 30158 74846 30210 74898
rect 30494 74846 30546 74898
rect 30606 74846 30658 74898
rect 34750 74846 34802 74898
rect 34974 74846 35026 74898
rect 36878 74846 36930 74898
rect 38222 74846 38274 74898
rect 4398 74734 4450 74786
rect 6526 74734 6578 74786
rect 8094 74734 8146 74786
rect 11006 74734 11058 74786
rect 13694 74734 13746 74786
rect 18062 74734 18114 74786
rect 19742 74734 19794 74786
rect 21870 74734 21922 74786
rect 23550 74734 23602 74786
rect 29262 74734 29314 74786
rect 35758 74734 35810 74786
rect 37662 74734 37714 74786
rect 25566 74622 25618 74674
rect 34414 74622 34466 74674
rect 35982 74622 36034 74674
rect 4478 74454 4530 74506
rect 4582 74454 4634 74506
rect 4686 74454 4738 74506
rect 35198 74454 35250 74506
rect 35302 74454 35354 74506
rect 35406 74454 35458 74506
rect 7198 74286 7250 74338
rect 7758 74286 7810 74338
rect 18846 74286 18898 74338
rect 19630 74286 19682 74338
rect 27806 74286 27858 74338
rect 29710 74286 29762 74338
rect 30158 74286 30210 74338
rect 35758 74286 35810 74338
rect 36206 74286 36258 74338
rect 2158 74174 2210 74226
rect 4286 74174 4338 74226
rect 7758 74174 7810 74226
rect 8430 74174 8482 74226
rect 19070 74174 19122 74226
rect 19966 74174 20018 74226
rect 21422 74174 21474 74226
rect 23662 74174 23714 74226
rect 29822 74174 29874 74226
rect 30270 74174 30322 74226
rect 30718 74174 30770 74226
rect 38334 74174 38386 74226
rect 5070 74062 5122 74114
rect 5742 74062 5794 74114
rect 6078 74062 6130 74114
rect 6638 74062 6690 74114
rect 6974 74062 7026 74114
rect 7310 74062 7362 74114
rect 14366 74062 14418 74114
rect 19854 74062 19906 74114
rect 20078 74062 20130 74114
rect 20526 74062 20578 74114
rect 26126 74062 26178 74114
rect 28142 74062 28194 74114
rect 28366 74062 28418 74114
rect 33742 74062 33794 74114
rect 33966 74062 34018 74114
rect 34974 74062 35026 74114
rect 35310 74062 35362 74114
rect 35646 74062 35698 74114
rect 36318 74062 36370 74114
rect 5854 73950 5906 74002
rect 6750 73950 6802 74002
rect 15822 73950 15874 74002
rect 29262 73950 29314 74002
rect 29374 73950 29426 74002
rect 33518 73950 33570 74002
rect 35198 73950 35250 74002
rect 19518 73838 19570 73890
rect 29038 73838 29090 73890
rect 33854 73838 33906 73890
rect 35758 73838 35810 73890
rect 19838 73670 19890 73722
rect 19942 73670 19994 73722
rect 20046 73670 20098 73722
rect 5294 73502 5346 73554
rect 6190 73502 6242 73554
rect 17502 73502 17554 73554
rect 17838 73502 17890 73554
rect 17950 73502 18002 73554
rect 18846 73502 18898 73554
rect 26238 73502 26290 73554
rect 27246 73502 27298 73554
rect 28702 73502 28754 73554
rect 30494 73502 30546 73554
rect 31502 73502 31554 73554
rect 16046 73390 16098 73442
rect 23102 73390 23154 73442
rect 29822 73390 29874 73442
rect 31054 73390 31106 73442
rect 16830 73278 16882 73330
rect 17726 73278 17778 73330
rect 19406 73278 19458 73330
rect 26126 73278 26178 73330
rect 26910 73278 26962 73330
rect 28366 73278 28418 73330
rect 29038 73278 29090 73330
rect 29598 73278 29650 73330
rect 30158 73278 30210 73330
rect 13918 73166 13970 73218
rect 18398 73166 18450 73218
rect 26238 73166 26290 73218
rect 29262 73166 29314 73218
rect 29710 73166 29762 73218
rect 30606 73166 30658 73218
rect 4478 72886 4530 72938
rect 4582 72886 4634 72938
rect 4686 72886 4738 72938
rect 35198 72886 35250 72938
rect 35302 72886 35354 72938
rect 35406 72886 35458 72938
rect 28254 72718 28306 72770
rect 15150 72606 15202 72658
rect 22206 72606 22258 72658
rect 29822 72606 29874 72658
rect 31950 72606 32002 72658
rect 35086 72606 35138 72658
rect 11790 72494 11842 72546
rect 13694 72494 13746 72546
rect 19966 72494 20018 72546
rect 20414 72494 20466 72546
rect 27806 72494 27858 72546
rect 29374 72494 29426 72546
rect 31278 72494 31330 72546
rect 25006 72382 25058 72434
rect 28254 72382 28306 72434
rect 28366 72382 28418 72434
rect 29262 72382 29314 72434
rect 11566 72270 11618 72322
rect 13470 72270 13522 72322
rect 33630 72270 33682 72322
rect 34078 72270 34130 72322
rect 34638 72270 34690 72322
rect 35646 72270 35698 72322
rect 36094 72270 36146 72322
rect 19838 72102 19890 72154
rect 19942 72102 19994 72154
rect 20046 72102 20098 72154
rect 26126 71934 26178 71986
rect 26238 71934 26290 71986
rect 32398 71934 32450 71986
rect 36766 71934 36818 71986
rect 8542 71822 8594 71874
rect 22542 71822 22594 71874
rect 29934 71822 29986 71874
rect 33294 71822 33346 71874
rect 34414 71822 34466 71874
rect 34862 71822 34914 71874
rect 35982 71822 36034 71874
rect 8878 71710 8930 71762
rect 11118 71710 11170 71762
rect 14478 71710 14530 71762
rect 17502 71710 17554 71762
rect 18846 71710 18898 71762
rect 21870 71710 21922 71762
rect 25566 71710 25618 71762
rect 26014 71710 26066 71762
rect 27806 71710 27858 71762
rect 34190 71710 34242 71762
rect 34974 71710 35026 71762
rect 36094 71710 36146 71762
rect 36318 71710 36370 71762
rect 9998 71598 10050 71650
rect 11790 71598 11842 71650
rect 13918 71598 13970 71650
rect 21086 71598 21138 71650
rect 24670 71598 24722 71650
rect 25790 71598 25842 71650
rect 33966 71598 34018 71650
rect 37214 71598 37266 71650
rect 37662 71598 37714 71650
rect 33406 71486 33458 71538
rect 34862 71486 34914 71538
rect 35534 71486 35586 71538
rect 4478 71318 4530 71370
rect 4582 71318 4634 71370
rect 4686 71318 4738 71370
rect 35198 71318 35250 71370
rect 35302 71318 35354 71370
rect 35406 71318 35458 71370
rect 13470 71150 13522 71202
rect 13806 71150 13858 71202
rect 7534 71038 7586 71090
rect 9662 71038 9714 71090
rect 10782 71038 10834 71090
rect 12910 71038 12962 71090
rect 14478 71038 14530 71090
rect 17838 71038 17890 71090
rect 18286 71038 18338 71090
rect 22430 71038 22482 71090
rect 25006 71038 25058 71090
rect 30158 71038 30210 71090
rect 32510 71038 32562 71090
rect 37214 71038 37266 71090
rect 6750 70926 6802 70978
rect 9998 70926 10050 70978
rect 14030 70926 14082 70978
rect 15038 70926 15090 70978
rect 23886 70926 23938 70978
rect 25230 70926 25282 70978
rect 25566 70926 25618 70978
rect 26798 70926 26850 70978
rect 27358 70926 27410 70978
rect 29374 70926 29426 70978
rect 31726 70926 31778 70978
rect 32734 70926 32786 70978
rect 33742 70926 33794 70978
rect 35310 70926 35362 70978
rect 5630 70814 5682 70866
rect 15710 70814 15762 70866
rect 25790 70814 25842 70866
rect 27694 70814 27746 70866
rect 28030 70814 28082 70866
rect 31054 70814 31106 70866
rect 32622 70814 32674 70866
rect 35422 70814 35474 70866
rect 38222 70814 38274 70866
rect 5966 70702 6018 70754
rect 14590 70702 14642 70754
rect 18398 70702 18450 70754
rect 18846 70702 18898 70754
rect 24334 70702 24386 70754
rect 25454 70702 25506 70754
rect 26462 70702 26514 70754
rect 27918 70702 27970 70754
rect 36094 70702 36146 70754
rect 19838 70534 19890 70586
rect 19942 70534 19994 70586
rect 20046 70534 20098 70586
rect 11566 70366 11618 70418
rect 15262 70366 15314 70418
rect 15934 70366 15986 70418
rect 25342 70366 25394 70418
rect 26238 70366 26290 70418
rect 26462 70366 26514 70418
rect 27470 70366 27522 70418
rect 28142 70366 28194 70418
rect 33630 70366 33682 70418
rect 34078 70366 34130 70418
rect 6190 70254 6242 70306
rect 10670 70254 10722 70306
rect 12686 70254 12738 70306
rect 15710 70254 15762 70306
rect 18398 70254 18450 70306
rect 26686 70254 26738 70306
rect 28254 70254 28306 70306
rect 28926 70254 28978 70306
rect 30606 70254 30658 70306
rect 30830 70254 30882 70306
rect 34302 70254 34354 70306
rect 5518 70142 5570 70194
rect 11902 70142 11954 70194
rect 15598 70142 15650 70194
rect 18958 70142 19010 70194
rect 22318 70142 22370 70194
rect 26126 70142 26178 70194
rect 26798 70142 26850 70194
rect 27246 70142 27298 70194
rect 27582 70142 27634 70194
rect 27918 70142 27970 70194
rect 29150 70142 29202 70194
rect 30382 70142 30434 70194
rect 31166 70142 31218 70194
rect 31838 70142 31890 70194
rect 32174 70142 32226 70194
rect 33070 70142 33122 70194
rect 33294 70142 33346 70194
rect 33518 70142 33570 70194
rect 33742 70142 33794 70194
rect 34414 70142 34466 70194
rect 34862 70142 34914 70194
rect 36990 70142 37042 70194
rect 8318 70030 8370 70082
rect 8766 70030 8818 70082
rect 9886 70030 9938 70082
rect 10110 70030 10162 70082
rect 10334 70030 10386 70082
rect 11006 70030 11058 70082
rect 14814 70030 14866 70082
rect 16270 70030 16322 70082
rect 17838 70030 17890 70082
rect 18174 70030 18226 70082
rect 18510 70030 18562 70082
rect 19630 70030 19682 70082
rect 21758 70030 21810 70082
rect 25902 70030 25954 70082
rect 28478 70030 28530 70082
rect 29486 70030 29538 70082
rect 37326 70030 37378 70082
rect 11230 69918 11282 69970
rect 28702 69918 28754 69970
rect 29710 69918 29762 69970
rect 30046 69918 30098 69970
rect 32174 69918 32226 69970
rect 35758 69918 35810 69970
rect 4478 69750 4530 69802
rect 4582 69750 4634 69802
rect 4686 69750 4738 69802
rect 35198 69750 35250 69802
rect 35302 69750 35354 69802
rect 35406 69750 35458 69802
rect 5630 69582 5682 69634
rect 6750 69582 6802 69634
rect 7086 69582 7138 69634
rect 9102 69582 9154 69634
rect 26798 69582 26850 69634
rect 32174 69582 32226 69634
rect 5070 69470 5122 69522
rect 9550 69470 9602 69522
rect 10670 69470 10722 69522
rect 13582 69470 13634 69522
rect 14030 69470 14082 69522
rect 14478 69470 14530 69522
rect 17726 69470 17778 69522
rect 18174 69470 18226 69522
rect 28366 69470 28418 69522
rect 31390 69470 31442 69522
rect 32958 69470 33010 69522
rect 35646 69470 35698 69522
rect 38222 69470 38274 69522
rect 2158 69358 2210 69410
rect 5966 69358 6018 69410
rect 6190 69358 6242 69410
rect 8766 69358 8818 69410
rect 11230 69358 11282 69410
rect 14814 69358 14866 69410
rect 22094 69358 22146 69410
rect 26686 69358 26738 69410
rect 27358 69358 27410 69410
rect 27694 69358 27746 69410
rect 29150 69358 29202 69410
rect 29598 69358 29650 69410
rect 30270 69358 30322 69410
rect 31838 69358 31890 69410
rect 32846 69358 32898 69410
rect 34862 69358 34914 69410
rect 35870 69358 35922 69410
rect 36990 69358 37042 69410
rect 2942 69246 2994 69298
rect 8542 69246 8594 69298
rect 11566 69246 11618 69298
rect 15598 69246 15650 69298
rect 24446 69246 24498 69298
rect 27918 69246 27970 69298
rect 29486 69246 29538 69298
rect 33406 69246 33458 69298
rect 34526 69246 34578 69298
rect 37214 69246 37266 69298
rect 37326 69246 37378 69298
rect 6638 69134 6690 69186
rect 7086 69134 7138 69186
rect 9998 69134 10050 69186
rect 18062 69134 18114 69186
rect 29374 69134 29426 69186
rect 32062 69134 32114 69186
rect 37774 69134 37826 69186
rect 19838 68966 19890 69018
rect 19942 68966 19994 69018
rect 20046 68966 20098 69018
rect 3502 68798 3554 68850
rect 15822 68798 15874 68850
rect 16270 68798 16322 68850
rect 28254 68798 28306 68850
rect 28478 68798 28530 68850
rect 30942 68798 30994 68850
rect 33182 68798 33234 68850
rect 16382 68686 16434 68738
rect 20750 68686 20802 68738
rect 21198 68686 21250 68738
rect 33070 68686 33122 68738
rect 3838 68574 3890 68626
rect 4510 68574 4562 68626
rect 6078 68574 6130 68626
rect 17502 68574 17554 68626
rect 28590 68574 28642 68626
rect 31614 68574 31666 68626
rect 32622 68574 32674 68626
rect 33966 68574 34018 68626
rect 36094 68574 36146 68626
rect 36766 68574 36818 68626
rect 6862 68462 6914 68514
rect 8990 68462 9042 68514
rect 9550 68462 9602 68514
rect 10110 68462 10162 68514
rect 10558 68462 10610 68514
rect 15374 68462 15426 68514
rect 18174 68462 18226 68514
rect 20302 68462 20354 68514
rect 29038 68462 29090 68514
rect 29374 68462 29426 68514
rect 29486 68462 29538 68514
rect 5294 68350 5346 68402
rect 9886 68350 9938 68402
rect 16158 68350 16210 68402
rect 21086 68350 21138 68402
rect 30046 68462 30098 68514
rect 30382 68462 30434 68514
rect 31950 68462 32002 68514
rect 34974 68462 35026 68514
rect 37550 68462 37602 68514
rect 30382 68350 30434 68402
rect 31838 68350 31890 68402
rect 35198 68350 35250 68402
rect 4478 68182 4530 68234
rect 4582 68182 4634 68234
rect 4686 68182 4738 68234
rect 35198 68182 35250 68234
rect 35302 68182 35354 68234
rect 35406 68182 35458 68234
rect 8878 68014 8930 68066
rect 9214 68014 9266 68066
rect 17950 68014 18002 68066
rect 31950 68014 32002 68066
rect 33070 68014 33122 68066
rect 34414 68014 34466 68066
rect 34750 68014 34802 68066
rect 36878 68014 36930 68066
rect 9214 67902 9266 67954
rect 18622 67902 18674 67954
rect 19742 67902 19794 67954
rect 20190 67902 20242 67954
rect 24110 67902 24162 67954
rect 29598 67902 29650 67954
rect 31726 67902 31778 67954
rect 37326 67902 37378 67954
rect 20526 67790 20578 67842
rect 27022 67790 27074 67842
rect 27470 67790 27522 67842
rect 31278 67790 31330 67842
rect 33630 67790 33682 67842
rect 35534 67790 35586 67842
rect 36094 67790 36146 67842
rect 37550 67790 37602 67842
rect 37774 67790 37826 67842
rect 3166 67678 3218 67730
rect 7870 67678 7922 67730
rect 8206 67678 8258 67730
rect 16830 67678 16882 67730
rect 17614 67678 17666 67730
rect 17838 67678 17890 67730
rect 20638 67678 20690 67730
rect 23102 67678 23154 67730
rect 26238 67678 26290 67730
rect 30382 67678 30434 67730
rect 30718 67678 30770 67730
rect 31726 67678 31778 67730
rect 33182 67678 33234 67730
rect 33854 67678 33906 67730
rect 35310 67678 35362 67730
rect 2830 67566 2882 67618
rect 5742 67566 5794 67618
rect 17390 67566 17442 67618
rect 19406 67566 19458 67618
rect 19630 67566 19682 67618
rect 20862 67566 20914 67618
rect 21534 67566 21586 67618
rect 36094 67566 36146 67618
rect 19838 67398 19890 67450
rect 19942 67398 19994 67450
rect 20046 67398 20098 67450
rect 35086 67230 35138 67282
rect 2494 67118 2546 67170
rect 11118 67118 11170 67170
rect 20750 67118 20802 67170
rect 29262 67118 29314 67170
rect 30494 67118 30546 67170
rect 33406 67118 33458 67170
rect 34190 67118 34242 67170
rect 37438 67118 37490 67170
rect 1822 67006 1874 67058
rect 8766 67006 8818 67058
rect 15038 67006 15090 67058
rect 17614 67006 17666 67058
rect 17950 67006 18002 67058
rect 18734 67006 18786 67058
rect 19294 67006 19346 67058
rect 20078 67006 20130 67058
rect 29150 67006 29202 67058
rect 29486 67006 29538 67058
rect 33630 67006 33682 67058
rect 34302 67006 34354 67058
rect 35982 67006 36034 67058
rect 37886 67006 37938 67058
rect 4622 66894 4674 66946
rect 5070 66894 5122 66946
rect 8430 66894 8482 66946
rect 8990 66894 9042 66946
rect 15486 66894 15538 66946
rect 16046 66894 16098 66946
rect 16494 66894 16546 66946
rect 16942 66894 16994 66946
rect 18174 66894 18226 66946
rect 22878 66894 22930 66946
rect 23438 66894 23490 66946
rect 23886 66894 23938 66946
rect 24334 66894 24386 66946
rect 24782 66894 24834 66946
rect 30046 66894 30098 66946
rect 30942 66894 30994 66946
rect 31390 66894 31442 66946
rect 15262 66782 15314 66834
rect 16494 66782 16546 66834
rect 19070 66782 19122 66834
rect 23998 66782 24050 66834
rect 24334 66782 24386 66834
rect 24782 66782 24834 66834
rect 4478 66614 4530 66666
rect 4582 66614 4634 66666
rect 4686 66614 4738 66666
rect 35198 66614 35250 66666
rect 35302 66614 35354 66666
rect 35406 66614 35458 66666
rect 3390 66446 3442 66498
rect 17390 66446 17442 66498
rect 19182 66446 19234 66498
rect 29262 66446 29314 66498
rect 30046 66446 30098 66498
rect 30382 66446 30434 66498
rect 32958 66446 33010 66498
rect 5070 66334 5122 66386
rect 8654 66334 8706 66386
rect 9998 66334 10050 66386
rect 10894 66334 10946 66386
rect 14814 66334 14866 66386
rect 15598 66334 15650 66386
rect 16606 66334 16658 66386
rect 18734 66334 18786 66386
rect 21422 66334 21474 66386
rect 24894 66334 24946 66386
rect 26014 66334 26066 66386
rect 29710 66334 29762 66386
rect 31166 66334 31218 66386
rect 34638 66334 34690 66386
rect 3726 66222 3778 66274
rect 3950 66222 4002 66274
rect 4510 66222 4562 66274
rect 5854 66222 5906 66274
rect 9102 66222 9154 66274
rect 9326 66222 9378 66274
rect 10222 66222 10274 66274
rect 11118 66222 11170 66274
rect 16494 66222 16546 66274
rect 17726 66222 17778 66274
rect 17950 66222 18002 66274
rect 18174 66222 18226 66274
rect 18958 66222 19010 66274
rect 19406 66222 19458 66274
rect 20414 66222 20466 66274
rect 20638 66222 20690 66274
rect 22094 66222 22146 66274
rect 29486 66222 29538 66274
rect 30382 66222 30434 66274
rect 33294 66222 33346 66274
rect 34862 66222 34914 66274
rect 37326 66222 37378 66274
rect 6526 66110 6578 66162
rect 14254 66110 14306 66162
rect 22766 66110 22818 66162
rect 25230 66110 25282 66162
rect 25566 66110 25618 66162
rect 29822 66110 29874 66162
rect 30718 66110 30770 66162
rect 31838 66110 31890 66162
rect 33518 66110 33570 66162
rect 35422 66110 35474 66162
rect 37550 66110 37602 66162
rect 4286 65998 4338 66050
rect 9662 65998 9714 66050
rect 10558 65998 10610 66050
rect 11454 65998 11506 66050
rect 11902 65998 11954 66050
rect 14142 65998 14194 66050
rect 36318 65998 36370 66050
rect 36990 65998 37042 66050
rect 19838 65830 19890 65882
rect 19942 65830 19994 65882
rect 20046 65830 20098 65882
rect 9886 65662 9938 65714
rect 10782 65662 10834 65714
rect 22654 65662 22706 65714
rect 25790 65662 25842 65714
rect 33294 65662 33346 65714
rect 3614 65550 3666 65602
rect 7086 65550 7138 65602
rect 16270 65550 16322 65602
rect 17502 65550 17554 65602
rect 20526 65550 20578 65602
rect 30942 65550 30994 65602
rect 32398 65550 32450 65602
rect 33854 65550 33906 65602
rect 2942 65438 2994 65490
rect 7422 65438 7474 65490
rect 11790 65438 11842 65490
rect 15038 65438 15090 65490
rect 15598 65438 15650 65490
rect 19070 65438 19122 65490
rect 21198 65438 21250 65490
rect 22318 65438 22370 65490
rect 22990 65438 23042 65490
rect 23214 65438 23266 65490
rect 23438 65438 23490 65490
rect 23886 65438 23938 65490
rect 23998 65438 24050 65490
rect 25230 65438 25282 65490
rect 28814 65438 28866 65490
rect 30046 65438 30098 65490
rect 30606 65438 30658 65490
rect 32174 65438 32226 65490
rect 32510 65438 32562 65490
rect 33406 65438 33458 65490
rect 34190 65438 34242 65490
rect 35198 65438 35250 65490
rect 35870 65438 35922 65490
rect 37438 65438 37490 65490
rect 5742 65326 5794 65378
rect 6190 65326 6242 65378
rect 8878 65326 8930 65378
rect 12462 65326 12514 65378
rect 14590 65326 14642 65378
rect 16046 65326 16098 65378
rect 16718 65326 16770 65378
rect 19182 65326 19234 65378
rect 21870 65326 21922 65378
rect 24222 65326 24274 65378
rect 24670 65326 24722 65378
rect 26238 65326 26290 65378
rect 26686 65326 26738 65378
rect 28590 65326 28642 65378
rect 31614 65326 31666 65378
rect 33518 65326 33570 65378
rect 34526 65326 34578 65378
rect 35982 65326 36034 65378
rect 37774 65326 37826 65378
rect 21758 65214 21810 65266
rect 25454 65214 25506 65266
rect 4478 65046 4530 65098
rect 4582 65046 4634 65098
rect 4686 65046 4738 65098
rect 35198 65046 35250 65098
rect 35302 65046 35354 65098
rect 35406 65046 35458 65098
rect 3838 64878 3890 64930
rect 7870 64878 7922 64930
rect 13470 64878 13522 64930
rect 15038 64878 15090 64930
rect 22990 64878 23042 64930
rect 26350 64878 26402 64930
rect 28590 64878 28642 64930
rect 29598 64878 29650 64930
rect 34974 64878 35026 64930
rect 35534 64878 35586 64930
rect 4174 64766 4226 64818
rect 4398 64766 4450 64818
rect 12462 64766 12514 64818
rect 13022 64766 13074 64818
rect 13582 64766 13634 64818
rect 22094 64766 22146 64818
rect 25118 64766 25170 64818
rect 25454 64766 25506 64818
rect 28030 64766 28082 64818
rect 33630 64766 33682 64818
rect 36318 64766 36370 64818
rect 36990 64766 37042 64818
rect 8206 64654 8258 64706
rect 8430 64654 8482 64706
rect 13806 64654 13858 64706
rect 14366 64654 14418 64706
rect 15038 64654 15090 64706
rect 15486 64654 15538 64706
rect 16046 64654 16098 64706
rect 18622 64654 18674 64706
rect 20750 64654 20802 64706
rect 21310 64654 21362 64706
rect 23326 64654 23378 64706
rect 23550 64654 23602 64706
rect 24110 64654 24162 64706
rect 24334 64654 24386 64706
rect 24894 64654 24946 64706
rect 25678 64654 25730 64706
rect 28254 64654 28306 64706
rect 31166 64654 31218 64706
rect 32622 64654 32674 64706
rect 33406 64654 33458 64706
rect 34078 64654 34130 64706
rect 34638 64654 34690 64706
rect 35870 64654 35922 64706
rect 36094 64654 36146 64706
rect 37102 64654 37154 64706
rect 37886 64654 37938 64706
rect 4846 64542 4898 64594
rect 16158 64542 16210 64594
rect 16942 64542 16994 64594
rect 19518 64542 19570 64594
rect 21646 64542 21698 64594
rect 22542 64542 22594 64594
rect 24670 64542 24722 64594
rect 26462 64542 26514 64594
rect 27806 64542 27858 64594
rect 29262 64542 29314 64594
rect 33070 64542 33122 64594
rect 34414 64542 34466 64594
rect 34862 64542 34914 64594
rect 37326 64542 37378 64594
rect 38222 64542 38274 64594
rect 7534 64430 7586 64482
rect 14030 64430 14082 64482
rect 14254 64430 14306 64482
rect 18510 64430 18562 64482
rect 21534 64430 21586 64482
rect 26014 64430 26066 64482
rect 26910 64430 26962 64482
rect 29486 64430 29538 64482
rect 30046 64430 30098 64482
rect 32062 64430 32114 64482
rect 32174 64430 32226 64482
rect 32286 64430 32338 64482
rect 38110 64430 38162 64482
rect 19838 64262 19890 64314
rect 19942 64262 19994 64314
rect 20046 64262 20098 64314
rect 16830 64094 16882 64146
rect 23214 64094 23266 64146
rect 25342 64094 25394 64146
rect 26238 64094 26290 64146
rect 28702 64094 28754 64146
rect 32062 64094 32114 64146
rect 12126 63982 12178 64034
rect 14590 63982 14642 64034
rect 16382 63982 16434 64034
rect 17502 63982 17554 64034
rect 19966 63982 20018 64034
rect 21870 63982 21922 64034
rect 27134 63982 27186 64034
rect 29150 63982 29202 64034
rect 29262 63982 29314 64034
rect 30382 63982 30434 64034
rect 30942 63982 30994 64034
rect 31950 63982 32002 64034
rect 32286 63982 32338 64034
rect 32510 63982 32562 64034
rect 33518 63982 33570 64034
rect 34638 63982 34690 64034
rect 36094 63982 36146 64034
rect 37438 63982 37490 64034
rect 11454 63870 11506 63922
rect 15150 63870 15202 63922
rect 15710 63870 15762 63922
rect 16270 63870 16322 63922
rect 17390 63870 17442 63922
rect 21198 63870 21250 63922
rect 22990 63870 23042 63922
rect 23550 63870 23602 63922
rect 23774 63870 23826 63922
rect 24222 63870 24274 63922
rect 24334 63870 24386 63922
rect 24558 63870 24610 63922
rect 25790 63870 25842 63922
rect 27806 63870 27858 63922
rect 28590 63870 28642 63922
rect 28926 63870 28978 63922
rect 29486 63870 29538 63922
rect 29934 63870 29986 63922
rect 30830 63870 30882 63922
rect 33854 63870 33906 63922
rect 35086 63870 35138 63922
rect 36318 63870 36370 63922
rect 38222 63870 38274 63922
rect 14254 63758 14306 63810
rect 19630 63758 19682 63810
rect 26686 63758 26738 63810
rect 28254 63758 28306 63810
rect 31278 63758 31330 63810
rect 14702 63646 14754 63698
rect 4478 63478 4530 63530
rect 4582 63478 4634 63530
rect 4686 63478 4738 63530
rect 35198 63478 35250 63530
rect 35302 63478 35354 63530
rect 35406 63478 35458 63530
rect 14030 63310 14082 63362
rect 15150 63310 15202 63362
rect 30718 63310 30770 63362
rect 33406 63310 33458 63362
rect 37550 63310 37602 63362
rect 11902 63198 11954 63250
rect 13470 63198 13522 63250
rect 18622 63198 18674 63250
rect 20750 63198 20802 63250
rect 27358 63198 27410 63250
rect 35982 63198 36034 63250
rect 8990 63086 9042 63138
rect 13694 63086 13746 63138
rect 15038 63086 15090 63138
rect 15486 63086 15538 63138
rect 16046 63086 16098 63138
rect 17950 63086 18002 63138
rect 21422 63086 21474 63138
rect 23102 63086 23154 63138
rect 24558 63086 24610 63138
rect 27806 63086 27858 63138
rect 29934 63086 29986 63138
rect 30606 63086 30658 63138
rect 30830 63086 30882 63138
rect 32174 63086 32226 63138
rect 33518 63086 33570 63138
rect 33854 63086 33906 63138
rect 35534 63086 35586 63138
rect 36094 63086 36146 63138
rect 37550 63086 37602 63138
rect 37886 63086 37938 63138
rect 6414 62974 6466 63026
rect 9774 62974 9826 63026
rect 14478 62974 14530 63026
rect 16158 62974 16210 63026
rect 16606 62974 16658 63026
rect 17278 62974 17330 63026
rect 21870 62974 21922 63026
rect 25230 62974 25282 63026
rect 29262 62974 29314 63026
rect 29598 62974 29650 63026
rect 35198 62974 35250 63026
rect 36430 62974 36482 63026
rect 6750 62862 6802 62914
rect 12350 62862 12402 62914
rect 16494 62862 16546 62914
rect 16830 62862 16882 62914
rect 17054 62862 17106 62914
rect 21422 62862 21474 62914
rect 19838 62694 19890 62746
rect 19942 62694 19994 62746
rect 20046 62694 20098 62746
rect 9662 62526 9714 62578
rect 9998 62526 10050 62578
rect 14254 62526 14306 62578
rect 14702 62526 14754 62578
rect 16830 62526 16882 62578
rect 18174 62526 18226 62578
rect 18622 62526 18674 62578
rect 19070 62526 19122 62578
rect 23102 62526 23154 62578
rect 29822 62526 29874 62578
rect 30494 62526 30546 62578
rect 37998 62526 38050 62578
rect 6526 62414 6578 62466
rect 20078 62414 20130 62466
rect 21198 62414 21250 62466
rect 25902 62414 25954 62466
rect 31726 62414 31778 62466
rect 32286 62414 32338 62466
rect 32622 62414 32674 62466
rect 1710 62302 1762 62354
rect 5742 62302 5794 62354
rect 10334 62302 10386 62354
rect 15374 62302 15426 62354
rect 16494 62302 16546 62354
rect 19406 62302 19458 62354
rect 21086 62302 21138 62354
rect 22990 62302 23042 62354
rect 25678 62302 25730 62354
rect 29486 62302 29538 62354
rect 32510 62302 32562 62354
rect 33630 62302 33682 62354
rect 34750 62302 34802 62354
rect 35086 62302 35138 62354
rect 36430 62302 36482 62354
rect 36654 62302 36706 62354
rect 2494 62190 2546 62242
rect 4622 62190 4674 62242
rect 5070 62190 5122 62242
rect 8654 62190 8706 62242
rect 15822 62190 15874 62242
rect 17726 62190 17778 62242
rect 29038 62190 29090 62242
rect 29262 62190 29314 62242
rect 31054 62190 31106 62242
rect 38110 62190 38162 62242
rect 16270 62078 16322 62130
rect 19518 62078 19570 62130
rect 34414 62078 34466 62130
rect 4478 61910 4530 61962
rect 4582 61910 4634 61962
rect 4686 61910 4738 61962
rect 35198 61910 35250 61962
rect 35302 61910 35354 61962
rect 35406 61910 35458 61962
rect 6190 61742 6242 61794
rect 14030 61742 14082 61794
rect 16158 61742 16210 61794
rect 16718 61742 16770 61794
rect 27582 61742 27634 61794
rect 27806 61742 27858 61794
rect 29710 61742 29762 61794
rect 5966 61630 6018 61682
rect 6526 61630 6578 61682
rect 9998 61630 10050 61682
rect 16158 61630 16210 61682
rect 17726 61630 17778 61682
rect 20750 61630 20802 61682
rect 21422 61630 21474 61682
rect 24446 61630 24498 61682
rect 26574 61630 26626 61682
rect 27806 61630 27858 61682
rect 29374 61630 29426 61682
rect 35758 61630 35810 61682
rect 37774 61630 37826 61682
rect 15150 61518 15202 61570
rect 20190 61518 20242 61570
rect 21758 61518 21810 61570
rect 27358 61518 27410 61570
rect 29486 61518 29538 61570
rect 30494 61518 30546 61570
rect 31838 61518 31890 61570
rect 32286 61518 32338 61570
rect 33182 61518 33234 61570
rect 33630 61518 33682 61570
rect 34414 61518 34466 61570
rect 35422 61518 35474 61570
rect 36990 61518 37042 61570
rect 2830 61406 2882 61458
rect 3166 61406 3218 61458
rect 6750 61406 6802 61458
rect 13918 61406 13970 61458
rect 14590 61406 14642 61458
rect 14702 61406 14754 61458
rect 17054 61406 17106 61458
rect 20302 61406 20354 61458
rect 20526 61406 20578 61458
rect 23102 61406 23154 61458
rect 30942 61406 30994 61458
rect 31726 61406 31778 61458
rect 33294 61406 33346 61458
rect 36206 61406 36258 61458
rect 37214 61406 37266 61458
rect 37438 61406 37490 61458
rect 4174 61294 4226 61346
rect 7646 61294 7698 61346
rect 8094 61294 8146 61346
rect 9102 61294 9154 61346
rect 14366 61294 14418 61346
rect 16606 61294 16658 61346
rect 20078 61294 20130 61346
rect 23886 61294 23938 61346
rect 28590 61294 28642 61346
rect 31950 61294 32002 61346
rect 19838 61126 19890 61178
rect 19942 61126 19994 61178
rect 20046 61126 20098 61178
rect 3390 60958 3442 61010
rect 7982 60958 8034 61010
rect 10334 60958 10386 61010
rect 18958 60958 19010 61010
rect 23214 60958 23266 61010
rect 23662 60958 23714 61010
rect 25342 60958 25394 61010
rect 32286 60958 32338 61010
rect 32398 60958 32450 61010
rect 5742 60846 5794 60898
rect 6862 60846 6914 60898
rect 7422 60846 7474 60898
rect 9550 60846 9602 60898
rect 19406 60846 19458 60898
rect 19518 60846 19570 60898
rect 21422 60846 21474 60898
rect 28254 60846 28306 60898
rect 4286 60734 4338 60786
rect 6190 60734 6242 60786
rect 6974 60734 7026 60786
rect 9886 60734 9938 60786
rect 10670 60734 10722 60786
rect 19182 60734 19234 60786
rect 21198 60734 21250 60786
rect 3950 60622 4002 60674
rect 5294 60622 5346 60674
rect 6302 60622 6354 60674
rect 10894 60622 10946 60674
rect 11454 60622 11506 60674
rect 20302 60622 20354 60674
rect 20750 60622 20802 60674
rect 3726 60510 3778 60562
rect 4510 60510 4562 60562
rect 4846 60510 4898 60562
rect 11118 60510 11170 60562
rect 11454 60510 11506 60562
rect 20302 60510 20354 60562
rect 20526 60510 20578 60562
rect 28366 60846 28418 60898
rect 32510 60846 32562 60898
rect 33742 60846 33794 60898
rect 34862 60846 34914 60898
rect 22766 60734 22818 60786
rect 25566 60734 25618 60786
rect 27470 60734 27522 60786
rect 27918 60734 27970 60786
rect 29150 60734 29202 60786
rect 29598 60734 29650 60786
rect 30494 60734 30546 60786
rect 30830 60734 30882 60786
rect 33070 60734 33122 60786
rect 34190 60734 34242 60786
rect 35310 60734 35362 60786
rect 36430 60734 36482 60786
rect 37662 60734 37714 60786
rect 21646 60622 21698 60674
rect 31502 60622 31554 60674
rect 33518 60622 33570 60674
rect 35982 60622 36034 60674
rect 28366 60510 28418 60562
rect 28814 60510 28866 60562
rect 29150 60510 29202 60562
rect 4478 60342 4530 60394
rect 4582 60342 4634 60394
rect 4686 60342 4738 60394
rect 35198 60342 35250 60394
rect 35302 60342 35354 60394
rect 35406 60342 35458 60394
rect 19070 60174 19122 60226
rect 24670 60174 24722 60226
rect 25006 60174 25058 60226
rect 25342 60174 25394 60226
rect 29598 60174 29650 60226
rect 33070 60174 33122 60226
rect 37550 60174 37602 60226
rect 4622 60062 4674 60114
rect 6974 60062 7026 60114
rect 9102 60062 9154 60114
rect 12462 60062 12514 60114
rect 14254 60062 14306 60114
rect 16382 60062 16434 60114
rect 18734 60062 18786 60114
rect 21646 60062 21698 60114
rect 22430 60062 22482 60114
rect 24222 60062 24274 60114
rect 24670 60062 24722 60114
rect 32062 60062 32114 60114
rect 34638 60062 34690 60114
rect 37662 60062 37714 60114
rect 1822 59950 1874 60002
rect 5854 59950 5906 60002
rect 7758 59950 7810 60002
rect 8430 59950 8482 60002
rect 12014 59950 12066 60002
rect 13470 59950 13522 60002
rect 18958 59950 19010 60002
rect 19406 59950 19458 60002
rect 20414 59950 20466 60002
rect 20638 59950 20690 60002
rect 21982 59950 22034 60002
rect 23662 59950 23714 60002
rect 23886 59950 23938 60002
rect 25678 59950 25730 60002
rect 26350 59950 26402 60002
rect 29598 59950 29650 60002
rect 29934 59950 29986 60002
rect 31278 59950 31330 60002
rect 34862 59950 34914 60002
rect 37886 59950 37938 60002
rect 2494 59838 2546 59890
rect 8542 59838 8594 59890
rect 11230 59838 11282 59890
rect 21310 59838 21362 59890
rect 21534 59838 21586 59890
rect 24110 59838 24162 59890
rect 25902 59838 25954 59890
rect 27694 59838 27746 59890
rect 29262 59838 29314 59890
rect 31838 59838 31890 59890
rect 32846 59838 32898 59890
rect 35870 59838 35922 59890
rect 5070 59726 5122 59778
rect 5630 59726 5682 59778
rect 7534 59726 7586 59778
rect 7646 59726 7698 59778
rect 16830 59726 16882 59778
rect 18174 59726 18226 59778
rect 23214 59726 23266 59778
rect 28254 59726 28306 59778
rect 28702 59726 28754 59778
rect 33406 59726 33458 59778
rect 36318 59726 36370 59778
rect 19838 59558 19890 59610
rect 19942 59558 19994 59610
rect 20046 59558 20098 59610
rect 8990 59390 9042 59442
rect 10110 59390 10162 59442
rect 14254 59390 14306 59442
rect 18734 59390 18786 59442
rect 25454 59390 25506 59442
rect 29822 59390 29874 59442
rect 37662 59390 37714 59442
rect 37886 59390 37938 59442
rect 4622 59278 4674 59330
rect 9550 59278 9602 59330
rect 15486 59278 15538 59330
rect 17502 59278 17554 59330
rect 19518 59278 19570 59330
rect 21534 59278 21586 59330
rect 27918 59278 27970 59330
rect 30942 59278 30994 59330
rect 31614 59278 31666 59330
rect 32398 59278 32450 59330
rect 36318 59278 36370 59330
rect 37998 59278 38050 59330
rect 3838 59166 3890 59218
rect 9774 59166 9826 59218
rect 10894 59166 10946 59218
rect 14590 59166 14642 59218
rect 15710 59166 15762 59218
rect 17390 59166 17442 59218
rect 17614 59166 17666 59218
rect 18062 59166 18114 59218
rect 18958 59166 19010 59218
rect 22766 59166 22818 59218
rect 24446 59166 24498 59218
rect 24670 59166 24722 59218
rect 27582 59166 27634 59218
rect 29710 59166 29762 59218
rect 30494 59166 30546 59218
rect 31726 59166 31778 59218
rect 33294 59166 33346 59218
rect 35310 59166 35362 59218
rect 36206 59166 36258 59218
rect 36430 59166 36482 59218
rect 37102 59166 37154 59218
rect 6750 59054 6802 59106
rect 7198 59054 7250 59106
rect 7646 59054 7698 59106
rect 8542 59054 8594 59106
rect 11678 59054 11730 59106
rect 13806 59054 13858 59106
rect 15150 59054 15202 59106
rect 16382 59054 16434 59106
rect 16830 59054 16882 59106
rect 20974 59054 21026 59106
rect 23214 59054 23266 59106
rect 23774 59054 23826 59106
rect 27358 59054 27410 59106
rect 31278 59054 31330 59106
rect 33518 59054 33570 59106
rect 6974 58942 7026 58994
rect 7534 58942 7586 58994
rect 14814 58942 14866 58994
rect 24110 58942 24162 58994
rect 32510 58942 32562 58994
rect 34190 58942 34242 58994
rect 4478 58774 4530 58826
rect 4582 58774 4634 58826
rect 4686 58774 4738 58826
rect 35198 58774 35250 58826
rect 35302 58774 35354 58826
rect 35406 58774 35458 58826
rect 7310 58494 7362 58546
rect 4398 58382 4450 58434
rect 4846 58382 4898 58434
rect 5070 58382 5122 58434
rect 6862 58382 6914 58434
rect 7198 58382 7250 58434
rect 7310 58270 7362 58322
rect 7534 58270 7586 58322
rect 7982 58606 8034 58658
rect 27806 58606 27858 58658
rect 28142 58606 28194 58658
rect 28478 58606 28530 58658
rect 29486 58606 29538 58658
rect 9102 58494 9154 58546
rect 11230 58494 11282 58546
rect 13582 58494 13634 58546
rect 14702 58494 14754 58546
rect 16830 58494 16882 58546
rect 18622 58494 18674 58546
rect 20750 58494 20802 58546
rect 22094 58494 22146 58546
rect 24222 58494 24274 58546
rect 28478 58494 28530 58546
rect 30270 58494 30322 58546
rect 32734 58494 32786 58546
rect 34862 58494 34914 58546
rect 37438 58494 37490 58546
rect 8430 58382 8482 58434
rect 14030 58382 14082 58434
rect 17838 58382 17890 58434
rect 21422 58382 21474 58434
rect 24670 58382 24722 58434
rect 29374 58382 29426 58434
rect 30606 58382 30658 58434
rect 31726 58382 31778 58434
rect 31950 58382 32002 58434
rect 33182 58382 33234 58434
rect 33854 58382 33906 58434
rect 35534 58382 35586 58434
rect 36990 58382 37042 58434
rect 17278 58270 17330 58322
rect 27694 58270 27746 58322
rect 29934 58270 29986 58322
rect 30158 58270 30210 58322
rect 33406 58270 33458 58322
rect 33518 58270 33570 58322
rect 36206 58270 36258 58322
rect 37102 58270 37154 58322
rect 4622 58158 4674 58210
rect 4734 58158 4786 58210
rect 5742 58158 5794 58210
rect 6190 58158 6242 58210
rect 6974 58158 7026 58210
rect 7870 58158 7922 58210
rect 11678 58158 11730 58210
rect 28030 58158 28082 58210
rect 29486 58158 29538 58210
rect 19838 57990 19890 58042
rect 19942 57990 19994 58042
rect 20046 57990 20098 58042
rect 7534 57822 7586 57874
rect 10894 57822 10946 57874
rect 12126 57822 12178 57874
rect 16046 57822 16098 57874
rect 16830 57822 16882 57874
rect 17614 57822 17666 57874
rect 17838 57822 17890 57874
rect 18062 57822 18114 57874
rect 22318 57822 22370 57874
rect 31614 57822 31666 57874
rect 32286 57822 32338 57874
rect 37886 57822 37938 57874
rect 5070 57710 5122 57762
rect 7086 57710 7138 57762
rect 14142 57710 14194 57762
rect 16158 57710 16210 57762
rect 17390 57710 17442 57762
rect 19182 57710 19234 57762
rect 20190 57710 20242 57762
rect 24222 57710 24274 57762
rect 24558 57710 24610 57762
rect 27806 57710 27858 57762
rect 32510 57710 32562 57762
rect 34302 57710 34354 57762
rect 36542 57710 36594 57762
rect 38222 57710 38274 57762
rect 1822 57598 1874 57650
rect 10670 57598 10722 57650
rect 12462 57598 12514 57650
rect 18062 57598 18114 57650
rect 19966 57598 20018 57650
rect 21870 57598 21922 57650
rect 23214 57598 23266 57650
rect 27918 57598 27970 57650
rect 30606 57598 30658 57650
rect 31054 57598 31106 57650
rect 33854 57598 33906 57650
rect 34190 57598 34242 57650
rect 35534 57598 35586 57650
rect 35870 57598 35922 57650
rect 37214 57598 37266 57650
rect 2494 57486 2546 57538
rect 4622 57486 4674 57538
rect 6862 57486 6914 57538
rect 15038 57486 15090 57538
rect 20414 57486 20466 57538
rect 22766 57486 22818 57538
rect 27134 57486 27186 57538
rect 28814 57486 28866 57538
rect 32174 57486 32226 57538
rect 35758 57486 35810 57538
rect 37102 57486 37154 57538
rect 6526 57374 6578 57426
rect 4478 57206 4530 57258
rect 4582 57206 4634 57258
rect 4686 57206 4738 57258
rect 35198 57206 35250 57258
rect 35302 57206 35354 57258
rect 35406 57206 35458 57258
rect 16942 56926 16994 56978
rect 17950 56926 18002 56978
rect 22094 56926 22146 56978
rect 25342 56926 25394 56978
rect 27470 56926 27522 56978
rect 31950 56926 32002 56978
rect 33518 56926 33570 56978
rect 33854 56926 33906 56978
rect 35198 56926 35250 56978
rect 35646 56926 35698 56978
rect 38334 56926 38386 56978
rect 3054 56814 3106 56866
rect 6862 56814 6914 56866
rect 17166 56814 17218 56866
rect 18286 56814 18338 56866
rect 18510 56814 18562 56866
rect 19294 56814 19346 56866
rect 24894 56814 24946 56866
rect 28142 56814 28194 56866
rect 29150 56814 29202 56866
rect 30158 56814 30210 56866
rect 30718 56814 30770 56866
rect 31278 56814 31330 56866
rect 34974 56814 35026 56866
rect 2830 56702 2882 56754
rect 14590 56702 14642 56754
rect 14702 56702 14754 56754
rect 24222 56702 24274 56754
rect 30270 56702 30322 56754
rect 30942 56702 30994 56754
rect 6638 56590 6690 56642
rect 14142 56590 14194 56642
rect 14366 56590 14418 56642
rect 15598 56590 15650 56642
rect 16606 56590 16658 56642
rect 17502 56590 17554 56642
rect 18846 56590 18898 56642
rect 19838 56422 19890 56474
rect 19942 56422 19994 56474
rect 20046 56422 20098 56474
rect 2830 56254 2882 56306
rect 11230 56254 11282 56306
rect 23886 56254 23938 56306
rect 25342 56254 25394 56306
rect 30942 56254 30994 56306
rect 17502 56142 17554 56194
rect 17838 56142 17890 56194
rect 18510 56142 18562 56194
rect 3166 56030 3218 56082
rect 11566 56030 11618 56082
rect 12238 56030 12290 56082
rect 23662 56030 23714 56082
rect 26686 56030 26738 56082
rect 11790 55918 11842 55970
rect 27470 55918 27522 55970
rect 29598 55918 29650 55970
rect 30046 55918 30098 55970
rect 30494 55918 30546 55970
rect 4478 55638 4530 55690
rect 4582 55638 4634 55690
rect 4686 55638 4738 55690
rect 35198 55638 35250 55690
rect 35302 55638 35354 55690
rect 35406 55638 35458 55690
rect 27694 55470 27746 55522
rect 28030 55470 28082 55522
rect 30382 55470 30434 55522
rect 3614 55358 3666 55410
rect 6526 55358 6578 55410
rect 8654 55358 8706 55410
rect 9774 55358 9826 55410
rect 19742 55358 19794 55410
rect 20638 55358 20690 55410
rect 22094 55358 22146 55410
rect 22542 55358 22594 55410
rect 24222 55358 24274 55410
rect 32286 55358 32338 55410
rect 3950 55246 4002 55298
rect 4174 55246 4226 55298
rect 5742 55246 5794 55298
rect 23326 55246 23378 55298
rect 25678 55246 25730 55298
rect 27918 55246 27970 55298
rect 28142 55246 28194 55298
rect 28478 55246 28530 55298
rect 29150 55246 29202 55298
rect 29374 55246 29426 55298
rect 31166 55246 31218 55298
rect 35422 55246 35474 55298
rect 24558 55134 24610 55186
rect 34862 55134 34914 55186
rect 4622 55022 4674 55074
rect 9326 55022 9378 55074
rect 12238 55022 12290 55074
rect 12686 55022 12738 55074
rect 17950 55022 18002 55074
rect 18510 55022 18562 55074
rect 21422 55022 21474 55074
rect 25566 55022 25618 55074
rect 28366 55022 28418 55074
rect 35758 55022 35810 55074
rect 19838 54854 19890 54906
rect 19942 54854 19994 54906
rect 20046 54854 20098 54906
rect 3614 54686 3666 54738
rect 11678 54686 11730 54738
rect 21870 54686 21922 54738
rect 23886 54686 23938 54738
rect 30046 54686 30098 54738
rect 6862 54574 6914 54626
rect 9550 54574 9602 54626
rect 10446 54574 10498 54626
rect 13022 54574 13074 54626
rect 18174 54574 18226 54626
rect 21422 54574 21474 54626
rect 27918 54574 27970 54626
rect 33182 54574 33234 54626
rect 6190 54462 6242 54514
rect 9774 54462 9826 54514
rect 10894 54462 10946 54514
rect 11230 54462 11282 54514
rect 12350 54462 12402 54514
rect 16830 54462 16882 54514
rect 17390 54462 17442 54514
rect 21198 54462 21250 54514
rect 28814 54462 28866 54514
rect 33406 54462 33458 54514
rect 35310 54462 35362 54514
rect 3950 54350 4002 54402
rect 4174 54350 4226 54402
rect 4622 54350 4674 54402
rect 8990 54350 9042 54402
rect 10446 54350 10498 54402
rect 15150 54350 15202 54402
rect 15598 54350 15650 54402
rect 20302 54350 20354 54402
rect 20750 54350 20802 54402
rect 22430 54350 22482 54402
rect 22878 54350 22930 54402
rect 23438 54350 23490 54402
rect 24446 54350 24498 54402
rect 27022 54350 27074 54402
rect 30158 54350 30210 54402
rect 36094 54350 36146 54402
rect 38222 54350 38274 54402
rect 24222 54238 24274 54290
rect 27358 54238 27410 54290
rect 27694 54238 27746 54290
rect 4478 54070 4530 54122
rect 4582 54070 4634 54122
rect 4686 54070 4738 54122
rect 35198 54070 35250 54122
rect 35302 54070 35354 54122
rect 35406 54070 35458 54122
rect 8206 53902 8258 53954
rect 8542 53902 8594 53954
rect 21310 53902 21362 53954
rect 21646 53902 21698 53954
rect 4846 53790 4898 53842
rect 10782 53790 10834 53842
rect 12910 53790 12962 53842
rect 17054 53790 17106 53842
rect 22878 53790 22930 53842
rect 32062 53790 32114 53842
rect 33182 53790 33234 53842
rect 35310 53790 35362 53842
rect 8990 53678 9042 53730
rect 10110 53678 10162 53730
rect 15822 53678 15874 53730
rect 16718 53678 16770 53730
rect 20414 53678 20466 53730
rect 26798 53678 26850 53730
rect 29150 53678 29202 53730
rect 32398 53678 32450 53730
rect 3726 53566 3778 53618
rect 7982 53566 8034 53618
rect 13470 53566 13522 53618
rect 13806 53566 13858 53618
rect 17838 53566 17890 53618
rect 19294 53566 19346 53618
rect 21870 53566 21922 53618
rect 22430 53566 22482 53618
rect 29934 53566 29986 53618
rect 35982 53566 36034 53618
rect 36318 53566 36370 53618
rect 36990 53566 37042 53618
rect 3390 53454 3442 53506
rect 5854 53454 5906 53506
rect 14254 53454 14306 53506
rect 16382 53454 16434 53506
rect 20638 53454 20690 53506
rect 20862 53454 20914 53506
rect 22094 53454 22146 53506
rect 22318 53454 22370 53506
rect 23438 53454 23490 53506
rect 27022 53454 27074 53506
rect 37326 53454 37378 53506
rect 38222 53454 38274 53506
rect 19838 53286 19890 53338
rect 19942 53286 19994 53338
rect 20046 53286 20098 53338
rect 5406 53118 5458 53170
rect 6302 53118 6354 53170
rect 7310 53118 7362 53170
rect 8654 53118 8706 53170
rect 11454 53118 11506 53170
rect 12350 53118 12402 53170
rect 16270 53118 16322 53170
rect 18846 53118 18898 53170
rect 22430 53118 22482 53170
rect 33070 53118 33122 53170
rect 34974 53118 35026 53170
rect 2494 53006 2546 53058
rect 8206 53006 8258 53058
rect 15150 53006 15202 53058
rect 16606 53006 16658 53058
rect 17502 53006 17554 53058
rect 18510 53006 18562 53058
rect 19406 53006 19458 53058
rect 21534 53006 21586 53058
rect 22094 53006 22146 53058
rect 22654 53006 22706 53058
rect 27358 53006 27410 53058
rect 31166 53006 31218 53058
rect 37438 53006 37490 53058
rect 1822 52894 1874 52946
rect 4958 52894 5010 52946
rect 5182 52894 5234 52946
rect 5630 52894 5682 52946
rect 6638 52894 6690 52946
rect 7982 52894 8034 52946
rect 12014 52894 12066 52946
rect 15822 52894 15874 52946
rect 19182 52894 19234 52946
rect 20078 52894 20130 52946
rect 20638 52894 20690 52946
rect 21310 52894 21362 52946
rect 21982 52894 22034 52946
rect 28030 52894 28082 52946
rect 30830 52894 30882 52946
rect 32286 52894 32338 52946
rect 38222 52894 38274 52946
rect 4622 52782 4674 52834
rect 5294 52782 5346 52834
rect 6862 52782 6914 52834
rect 11790 52782 11842 52834
rect 13022 52782 13074 52834
rect 23438 52782 23490 52834
rect 23886 52782 23938 52834
rect 25230 52782 25282 52834
rect 28590 52782 28642 52834
rect 33630 52782 33682 52834
rect 34078 52782 34130 52834
rect 35310 52782 35362 52834
rect 7646 52670 7698 52722
rect 17390 52670 17442 52722
rect 17726 52670 17778 52722
rect 20414 52670 20466 52722
rect 33406 52670 33458 52722
rect 4478 52502 4530 52554
rect 4582 52502 4634 52554
rect 4686 52502 4738 52554
rect 35198 52502 35250 52554
rect 35302 52502 35354 52554
rect 35406 52502 35458 52554
rect 35870 52334 35922 52386
rect 36990 52334 37042 52386
rect 4846 52222 4898 52274
rect 12910 52222 12962 52274
rect 14702 52222 14754 52274
rect 16830 52222 16882 52274
rect 17278 52222 17330 52274
rect 19294 52222 19346 52274
rect 22094 52222 22146 52274
rect 24222 52222 24274 52274
rect 31278 52222 31330 52274
rect 33406 52222 33458 52274
rect 33854 52222 33906 52274
rect 2046 52110 2098 52162
rect 6078 52110 6130 52162
rect 15598 52110 15650 52162
rect 16270 52110 16322 52162
rect 17726 52110 17778 52162
rect 18398 52110 18450 52162
rect 20078 52110 20130 52162
rect 20190 52110 20242 52162
rect 20862 52110 20914 52162
rect 21310 52110 21362 52162
rect 24670 52110 24722 52162
rect 25118 52110 25170 52162
rect 29374 52110 29426 52162
rect 29710 52110 29762 52162
rect 30494 52110 30546 52162
rect 35310 52110 35362 52162
rect 35534 52110 35586 52162
rect 36318 52110 36370 52162
rect 37326 52110 37378 52162
rect 37550 52110 37602 52162
rect 38222 52110 38274 52162
rect 2718 51998 2770 52050
rect 16046 51998 16098 52050
rect 18062 51998 18114 52050
rect 20302 51998 20354 52050
rect 20526 51998 20578 52050
rect 14590 51886 14642 51938
rect 15374 51886 15426 51938
rect 15822 51886 15874 51938
rect 15934 51886 15986 51938
rect 29486 51886 29538 51938
rect 30046 51886 30098 51938
rect 19838 51718 19890 51770
rect 19942 51718 19994 51770
rect 20046 51718 20098 51770
rect 3838 51550 3890 51602
rect 5070 51550 5122 51602
rect 16830 51550 16882 51602
rect 17838 51550 17890 51602
rect 24558 51550 24610 51602
rect 25342 51550 25394 51602
rect 25790 51550 25842 51602
rect 30718 51550 30770 51602
rect 31166 51550 31218 51602
rect 36654 51550 36706 51602
rect 3166 51438 3218 51490
rect 3502 51438 3554 51490
rect 18062 51438 18114 51490
rect 19294 51438 19346 51490
rect 21534 51438 21586 51490
rect 23550 51438 23602 51490
rect 4174 51326 4226 51378
rect 16382 51326 16434 51378
rect 19182 51326 19234 51378
rect 19966 51326 20018 51378
rect 20414 51326 20466 51378
rect 20638 51326 20690 51378
rect 20862 51326 20914 51378
rect 22990 51326 23042 51378
rect 30382 51326 30434 51378
rect 10782 51214 10834 51266
rect 15934 51214 15986 51266
rect 30158 51214 30210 51266
rect 18286 51102 18338 51154
rect 18622 51102 18674 51154
rect 4478 50934 4530 50986
rect 4582 50934 4634 50986
rect 4686 50934 4738 50986
rect 35198 50934 35250 50986
rect 35302 50934 35354 50986
rect 35406 50934 35458 50986
rect 6302 50766 6354 50818
rect 6638 50766 6690 50818
rect 7310 50654 7362 50706
rect 9438 50654 9490 50706
rect 11342 50654 11394 50706
rect 14702 50654 14754 50706
rect 16606 50654 16658 50706
rect 23438 50654 23490 50706
rect 26798 50654 26850 50706
rect 27694 50654 27746 50706
rect 35198 50654 35250 50706
rect 9326 50542 9378 50594
rect 9662 50542 9714 50594
rect 10894 50542 10946 50594
rect 18622 50542 18674 50594
rect 20750 50542 20802 50594
rect 21758 50542 21810 50594
rect 23998 50542 24050 50594
rect 27246 50542 27298 50594
rect 6862 50430 6914 50482
rect 8878 50430 8930 50482
rect 15374 50430 15426 50482
rect 15598 50430 15650 50482
rect 15710 50430 15762 50482
rect 18062 50430 18114 50482
rect 19518 50430 19570 50482
rect 21422 50430 21474 50482
rect 24670 50430 24722 50482
rect 10110 50318 10162 50370
rect 10558 50318 10610 50370
rect 15934 50318 15986 50370
rect 17054 50318 17106 50370
rect 22430 50318 22482 50370
rect 34862 50318 34914 50370
rect 19838 50150 19890 50202
rect 19942 50150 19994 50202
rect 20046 50150 20098 50202
rect 5070 49982 5122 50034
rect 11118 49982 11170 50034
rect 18062 49982 18114 50034
rect 19406 49982 19458 50034
rect 20526 49982 20578 50034
rect 35646 49982 35698 50034
rect 2494 49870 2546 49922
rect 10222 49870 10274 49922
rect 16270 49870 16322 49922
rect 18622 49870 18674 49922
rect 20302 49870 20354 49922
rect 20750 49870 20802 49922
rect 23326 49870 23378 49922
rect 25566 49870 25618 49922
rect 33630 49870 33682 49922
rect 1822 49758 1874 49810
rect 10446 49758 10498 49810
rect 11678 49758 11730 49810
rect 14814 49758 14866 49810
rect 15262 49758 15314 49810
rect 15934 49758 15986 49810
rect 16494 49758 16546 49810
rect 17502 49758 17554 49810
rect 20190 49758 20242 49810
rect 22318 49758 22370 49810
rect 24558 49758 24610 49810
rect 25230 49758 25282 49810
rect 26126 49758 26178 49810
rect 26910 49758 26962 49810
rect 33966 49758 34018 49810
rect 34974 49758 35026 49810
rect 4622 49646 4674 49698
rect 8206 49646 8258 49698
rect 12350 49646 12402 49698
rect 14478 49646 14530 49698
rect 19182 49646 19234 49698
rect 19854 49646 19906 49698
rect 22990 49646 23042 49698
rect 25902 49646 25954 49698
rect 27694 49646 27746 49698
rect 29822 49646 29874 49698
rect 30270 49646 30322 49698
rect 7982 49534 8034 49586
rect 8206 49534 8258 49586
rect 30718 49646 30770 49698
rect 34638 49646 34690 49698
rect 35198 49646 35250 49698
rect 19854 49534 19906 49586
rect 26462 49534 26514 49586
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 13470 49198 13522 49250
rect 21422 49198 21474 49250
rect 7982 49086 8034 49138
rect 8318 49086 8370 49138
rect 10446 49086 10498 49138
rect 11678 49086 11730 49138
rect 12462 49086 12514 49138
rect 13582 49086 13634 49138
rect 15262 49086 15314 49138
rect 16158 49086 16210 49138
rect 24894 49086 24946 49138
rect 27022 49086 27074 49138
rect 29710 49086 29762 49138
rect 30494 49086 30546 49138
rect 31166 49086 31218 49138
rect 31726 49086 31778 49138
rect 33854 49086 33906 49138
rect 7758 48974 7810 49026
rect 11230 48974 11282 49026
rect 13806 48974 13858 49026
rect 14478 48974 14530 49026
rect 16046 48974 16098 49026
rect 18622 48974 18674 49026
rect 20750 48974 20802 49026
rect 22654 48974 22706 49026
rect 22878 48974 22930 49026
rect 27694 48974 27746 49026
rect 30046 48974 30098 49026
rect 30270 48974 30322 49026
rect 34638 48974 34690 49026
rect 35310 48974 35362 49026
rect 35758 48974 35810 49026
rect 37102 48974 37154 49026
rect 7086 48862 7138 48914
rect 7422 48862 7474 48914
rect 14142 48862 14194 48914
rect 15598 48862 15650 48914
rect 17614 48862 17666 48914
rect 20190 48862 20242 48914
rect 22094 48862 22146 48914
rect 23102 48862 23154 48914
rect 30606 48862 30658 48914
rect 6750 48750 6802 48802
rect 13022 48750 13074 48802
rect 14254 48750 14306 48802
rect 14926 48750 14978 48802
rect 15822 48750 15874 48802
rect 16158 48750 16210 48802
rect 17054 48750 17106 48802
rect 28254 48750 28306 48802
rect 29262 48750 29314 48802
rect 30494 48750 30546 48802
rect 35198 48750 35250 48802
rect 35422 48750 35474 48802
rect 35534 48750 35586 48802
rect 36206 48750 36258 48802
rect 37326 48750 37378 48802
rect 38222 48750 38274 48802
rect 19838 48582 19890 48634
rect 19942 48582 19994 48634
rect 20046 48582 20098 48634
rect 9662 48414 9714 48466
rect 10222 48414 10274 48466
rect 10334 48414 10386 48466
rect 10446 48414 10498 48466
rect 11342 48414 11394 48466
rect 13918 48414 13970 48466
rect 19406 48414 19458 48466
rect 24222 48414 24274 48466
rect 24670 48414 24722 48466
rect 25342 48414 25394 48466
rect 27134 48414 27186 48466
rect 28030 48414 28082 48466
rect 33854 48414 33906 48466
rect 34190 48414 34242 48466
rect 34750 48414 34802 48466
rect 3726 48302 3778 48354
rect 6750 48302 6802 48354
rect 11902 48302 11954 48354
rect 14590 48302 14642 48354
rect 17950 48302 18002 48354
rect 21086 48302 21138 48354
rect 22990 48302 23042 48354
rect 26798 48302 26850 48354
rect 33630 48302 33682 48354
rect 37438 48302 37490 48354
rect 4062 48190 4114 48242
rect 4734 48190 4786 48242
rect 5966 48190 6018 48242
rect 9998 48190 10050 48242
rect 10670 48190 10722 48242
rect 15374 48190 15426 48242
rect 16158 48190 16210 48242
rect 16382 48190 16434 48242
rect 17390 48190 17442 48242
rect 21198 48190 21250 48242
rect 21870 48190 21922 48242
rect 22654 48190 22706 48242
rect 23886 48190 23938 48242
rect 25678 48190 25730 48242
rect 28478 48190 28530 48242
rect 34078 48190 34130 48242
rect 38110 48190 38162 48242
rect 5294 48078 5346 48130
rect 8878 48078 8930 48130
rect 12350 48078 12402 48130
rect 12798 48078 12850 48130
rect 14366 48078 14418 48130
rect 15822 48078 15874 48130
rect 16494 48078 16546 48130
rect 22206 48078 22258 48130
rect 23102 48078 23154 48130
rect 23662 48078 23714 48130
rect 26126 48078 26178 48130
rect 27582 48078 27634 48130
rect 29262 48078 29314 48130
rect 31390 48078 31442 48130
rect 32286 48078 32338 48130
rect 33182 48078 33234 48130
rect 33966 48078 34018 48130
rect 35310 48078 35362 48130
rect 5070 47966 5122 48018
rect 11678 47966 11730 48018
rect 14702 47966 14754 48018
rect 21646 47966 21698 48018
rect 31726 47966 31778 48018
rect 32062 47966 32114 48018
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 14254 47630 14306 47682
rect 14702 47630 14754 47682
rect 2942 47518 2994 47570
rect 5070 47518 5122 47570
rect 8990 47518 9042 47570
rect 12910 47518 12962 47570
rect 14366 47518 14418 47570
rect 14814 47518 14866 47570
rect 15486 47518 15538 47570
rect 24782 47518 24834 47570
rect 27470 47518 27522 47570
rect 34750 47518 34802 47570
rect 37550 47518 37602 47570
rect 2270 47406 2322 47458
rect 6078 47406 6130 47458
rect 9438 47406 9490 47458
rect 10110 47406 10162 47458
rect 15710 47406 15762 47458
rect 16494 47406 16546 47458
rect 18510 47406 18562 47458
rect 21870 47406 21922 47458
rect 29710 47406 29762 47458
rect 30830 47406 30882 47458
rect 31278 47406 31330 47458
rect 31838 47406 31890 47458
rect 35086 47406 35138 47458
rect 35534 47406 35586 47458
rect 35758 47406 35810 47458
rect 36206 47406 36258 47458
rect 37326 47406 37378 47458
rect 6862 47294 6914 47346
rect 10782 47294 10834 47346
rect 15038 47294 15090 47346
rect 15486 47294 15538 47346
rect 17054 47294 17106 47346
rect 19070 47294 19122 47346
rect 29486 47294 29538 47346
rect 31502 47294 31554 47346
rect 32622 47294 32674 47346
rect 36990 47294 37042 47346
rect 5742 47182 5794 47234
rect 13582 47182 13634 47234
rect 15262 47182 15314 47234
rect 16270 47182 16322 47234
rect 20078 47182 20130 47234
rect 20750 47182 20802 47234
rect 27022 47182 27074 47234
rect 27918 47182 27970 47234
rect 28366 47182 28418 47234
rect 35310 47182 35362 47234
rect 35422 47182 35474 47234
rect 36430 47182 36482 47234
rect 37998 47182 38050 47234
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 7422 46846 7474 46898
rect 10782 46846 10834 46898
rect 11006 46846 11058 46898
rect 11230 46846 11282 46898
rect 13806 46846 13858 46898
rect 14254 46846 14306 46898
rect 17838 46846 17890 46898
rect 24222 46846 24274 46898
rect 26238 46846 26290 46898
rect 27246 46846 27298 46898
rect 29598 46846 29650 46898
rect 33406 46846 33458 46898
rect 34638 46846 34690 46898
rect 35086 46846 35138 46898
rect 14142 46734 14194 46786
rect 19406 46734 19458 46786
rect 19966 46734 20018 46786
rect 23662 46734 23714 46786
rect 25230 46734 25282 46786
rect 37438 46734 37490 46786
rect 7758 46622 7810 46674
rect 11454 46622 11506 46674
rect 19518 46622 19570 46674
rect 21534 46622 21586 46674
rect 21982 46622 22034 46674
rect 24670 46622 24722 46674
rect 25454 46622 25506 46674
rect 25678 46622 25730 46674
rect 25790 46622 25842 46674
rect 27694 46622 27746 46674
rect 28590 46622 28642 46674
rect 38110 46622 38162 46674
rect 5294 46510 5346 46562
rect 9662 46510 9714 46562
rect 15038 46510 15090 46562
rect 15598 46510 15650 46562
rect 15934 46510 15986 46562
rect 16494 46510 16546 46562
rect 16830 46510 16882 46562
rect 22318 46510 22370 46562
rect 25566 46510 25618 46562
rect 26798 46510 26850 46562
rect 28142 46510 28194 46562
rect 29038 46510 29090 46562
rect 30158 46510 30210 46562
rect 30606 46510 30658 46562
rect 35310 46510 35362 46562
rect 14254 46398 14306 46450
rect 16046 46398 16098 46450
rect 16718 46398 16770 46450
rect 18286 46398 18338 46450
rect 26574 46398 26626 46450
rect 29934 46398 29986 46450
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 13470 46062 13522 46114
rect 37550 46062 37602 46114
rect 4622 45950 4674 46002
rect 14030 45950 14082 46002
rect 21758 45950 21810 46002
rect 30606 45950 30658 46002
rect 31054 45950 31106 46002
rect 36990 45950 37042 46002
rect 3950 45838 4002 45890
rect 4174 45838 4226 45890
rect 12910 45838 12962 45890
rect 13806 45838 13858 45890
rect 15934 45838 15986 45890
rect 16382 45838 16434 45890
rect 18398 45838 18450 45890
rect 20526 45838 20578 45890
rect 21534 45838 21586 45890
rect 24110 45838 24162 45890
rect 26238 45838 26290 45890
rect 28478 45838 28530 45890
rect 37214 45838 37266 45890
rect 16158 45726 16210 45778
rect 16830 45726 16882 45778
rect 19854 45726 19906 45778
rect 22766 45726 22818 45778
rect 23550 45726 23602 45778
rect 23662 45726 23714 45778
rect 23886 45726 23938 45778
rect 24222 45726 24274 45778
rect 26798 45726 26850 45778
rect 28366 45726 28418 45778
rect 3614 45614 3666 45666
rect 14814 45614 14866 45666
rect 15150 45614 15202 45666
rect 15598 45614 15650 45666
rect 16942 45614 16994 45666
rect 27806 45614 27858 45666
rect 28142 45614 28194 45666
rect 29262 45614 29314 45666
rect 29710 45614 29762 45666
rect 30158 45614 30210 45666
rect 34974 45614 35026 45666
rect 36430 45614 36482 45666
rect 38222 45614 38274 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 7982 45278 8034 45330
rect 11342 45278 11394 45330
rect 14366 45278 14418 45330
rect 17502 45278 17554 45330
rect 25342 45278 25394 45330
rect 17950 45166 18002 45218
rect 23214 45166 23266 45218
rect 25566 45166 25618 45218
rect 26014 45166 26066 45218
rect 28254 45166 28306 45218
rect 1822 45054 1874 45106
rect 14030 45054 14082 45106
rect 15374 45054 15426 45106
rect 17502 45054 17554 45106
rect 19182 45054 19234 45106
rect 20526 45054 20578 45106
rect 23438 45054 23490 45106
rect 23662 45054 23714 45106
rect 27134 45110 27186 45162
rect 23774 45054 23826 45106
rect 26350 45054 26402 45106
rect 26574 45054 26626 45106
rect 26910 45054 26962 45106
rect 27582 45054 27634 45106
rect 2494 44942 2546 44994
rect 4622 44942 4674 44994
rect 5070 44942 5122 44994
rect 7646 44942 7698 44994
rect 8542 44942 8594 44994
rect 11006 44942 11058 44994
rect 11678 44942 11730 44994
rect 11902 44942 11954 44994
rect 12462 44942 12514 44994
rect 14814 44942 14866 44994
rect 15262 44942 15314 44994
rect 16830 44942 16882 44994
rect 30382 44942 30434 44994
rect 30830 44942 30882 44994
rect 31278 44942 31330 44994
rect 31726 44942 31778 44994
rect 8318 44830 8370 44882
rect 21310 44830 21362 44882
rect 24222 44830 24274 44882
rect 27246 44830 27298 44882
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 14478 44382 14530 44434
rect 20302 44382 20354 44434
rect 20750 44382 20802 44434
rect 22542 44382 22594 44434
rect 28478 44382 28530 44434
rect 29710 44382 29762 44434
rect 31950 44382 32002 44434
rect 2270 44270 2322 44322
rect 3278 44270 3330 44322
rect 3614 44270 3666 44322
rect 3950 44270 4002 44322
rect 4174 44270 4226 44322
rect 15934 44270 15986 44322
rect 18062 44270 18114 44322
rect 21310 44270 21362 44322
rect 24670 44270 24722 44322
rect 26798 44270 26850 44322
rect 27134 44270 27186 44322
rect 27358 44270 27410 44322
rect 27582 44270 27634 44322
rect 30270 44270 30322 44322
rect 30494 44270 30546 44322
rect 32398 44270 32450 44322
rect 2942 44158 2994 44210
rect 6638 44158 6690 44210
rect 17054 44158 17106 44210
rect 18510 44158 18562 44210
rect 21534 44158 21586 44210
rect 22206 44158 22258 44210
rect 23662 44158 23714 44210
rect 25006 44158 25058 44210
rect 25678 44158 25730 44210
rect 29262 44158 29314 44210
rect 30606 44158 30658 44210
rect 31166 44158 31218 44210
rect 2606 44046 2658 44098
rect 4622 44046 4674 44098
rect 6974 44046 7026 44098
rect 15150 44046 15202 44098
rect 15598 44046 15650 44098
rect 18174 44046 18226 44098
rect 27918 44046 27970 44098
rect 30382 44046 30434 44098
rect 30718 44046 30770 44098
rect 31502 44046 31554 44098
rect 32846 44046 32898 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 19294 43710 19346 43762
rect 24670 43710 24722 43762
rect 2942 43598 2994 43650
rect 16382 43598 16434 43650
rect 17614 43598 17666 43650
rect 17838 43598 17890 43650
rect 20414 43598 20466 43650
rect 23438 43598 23490 43650
rect 23662 43598 23714 43650
rect 23774 43598 23826 43650
rect 29038 43598 29090 43650
rect 31726 43598 31778 43650
rect 2158 43486 2210 43538
rect 5518 43486 5570 43538
rect 6190 43486 6242 43538
rect 11454 43486 11506 43538
rect 15150 43486 15202 43538
rect 16158 43486 16210 43538
rect 16718 43486 16770 43538
rect 16942 43486 16994 43538
rect 19518 43486 19570 43538
rect 19854 43486 19906 43538
rect 21982 43486 22034 43538
rect 22542 43486 22594 43538
rect 23214 43486 23266 43538
rect 23998 43486 24050 43538
rect 24334 43486 24386 43538
rect 28366 43486 28418 43538
rect 32398 43486 32450 43538
rect 5070 43374 5122 43426
rect 6862 43374 6914 43426
rect 8990 43374 9042 43426
rect 9662 43374 9714 43426
rect 10110 43374 10162 43426
rect 12126 43374 12178 43426
rect 14254 43374 14306 43426
rect 25566 43374 25618 43426
rect 27694 43374 27746 43426
rect 29598 43374 29650 43426
rect 33182 43374 33234 43426
rect 34638 43374 34690 43426
rect 15374 43262 15426 43314
rect 15822 43262 15874 43314
rect 21870 43262 21922 43314
rect 34526 43262 34578 43314
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 6190 42926 6242 42978
rect 30046 42926 30098 42978
rect 30942 42926 30994 42978
rect 5630 42814 5682 42866
rect 7310 42814 7362 42866
rect 9438 42814 9490 42866
rect 16270 42814 16322 42866
rect 20750 42814 20802 42866
rect 27134 42814 27186 42866
rect 27918 42814 27970 42866
rect 29486 42814 29538 42866
rect 5070 42702 5122 42754
rect 5854 42702 5906 42754
rect 6638 42702 6690 42754
rect 10222 42702 10274 42754
rect 21534 42758 21586 42810
rect 31390 42814 31442 42866
rect 32286 42814 32338 42866
rect 33070 42814 33122 42866
rect 36430 42814 36482 42866
rect 38222 42814 38274 42866
rect 10334 42702 10386 42754
rect 12574 42702 12626 42754
rect 15150 42702 15202 42754
rect 18062 42702 18114 42754
rect 20302 42702 20354 42754
rect 21310 42702 21362 42754
rect 21758 42702 21810 42754
rect 24222 42702 24274 42754
rect 26350 42702 26402 42754
rect 27022 42702 27074 42754
rect 28142 42702 28194 42754
rect 29710 42702 29762 42754
rect 30606 42702 30658 42754
rect 35870 42702 35922 42754
rect 9774 42590 9826 42642
rect 9998 42590 10050 42642
rect 11342 42590 11394 42642
rect 12350 42590 12402 42642
rect 15374 42590 15426 42642
rect 15934 42590 15986 42642
rect 17614 42590 17666 42642
rect 19070 42590 19122 42642
rect 22542 42590 22594 42642
rect 25790 42590 25842 42642
rect 26798 42590 26850 42642
rect 30382 42590 30434 42642
rect 35198 42590 35250 42642
rect 36990 42590 37042 42642
rect 10110 42478 10162 42530
rect 11006 42478 11058 42530
rect 14366 42478 14418 42530
rect 14814 42478 14866 42530
rect 16718 42478 16770 42530
rect 22094 42478 22146 42530
rect 26238 42478 26290 42530
rect 31838 42478 31890 42530
rect 32734 42478 32786 42530
rect 37326 42478 37378 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 12574 42142 12626 42194
rect 15486 42142 15538 42194
rect 16382 42142 16434 42194
rect 16830 42142 16882 42194
rect 18958 42142 19010 42194
rect 25454 42142 25506 42194
rect 25678 42142 25730 42194
rect 26462 42142 26514 42194
rect 26686 42142 26738 42194
rect 27358 42142 27410 42194
rect 34862 42142 34914 42194
rect 5630 42030 5682 42082
rect 5854 42030 5906 42082
rect 9550 42030 9602 42082
rect 10894 42030 10946 42082
rect 15934 42030 15986 42082
rect 17502 42030 17554 42082
rect 20638 42030 20690 42082
rect 23326 42030 23378 42082
rect 29486 42030 29538 42082
rect 29934 42030 29986 42082
rect 31278 42030 31330 42082
rect 37438 42030 37490 42082
rect 6078 41918 6130 41970
rect 6302 41918 6354 41970
rect 8094 41918 8146 41970
rect 10558 41918 10610 41970
rect 13134 41918 13186 41970
rect 19182 41918 19234 41970
rect 19518 41918 19570 41970
rect 21646 41918 21698 41970
rect 21870 41918 21922 41970
rect 22094 41918 22146 41970
rect 23550 41918 23602 41970
rect 25230 41918 25282 41970
rect 26238 41918 26290 41970
rect 26798 41918 26850 41970
rect 27022 41918 27074 41970
rect 28926 41918 28978 41970
rect 30494 41918 30546 41970
rect 34638 41918 34690 41970
rect 38222 41918 38274 41970
rect 6190 41806 6242 41858
rect 7198 41806 7250 41858
rect 7646 41806 7698 41858
rect 9774 41806 9826 41858
rect 10110 41806 10162 41858
rect 11342 41806 11394 41858
rect 12350 41806 12402 41858
rect 12910 41806 12962 41858
rect 15038 41806 15090 41858
rect 22990 41806 23042 41858
rect 24446 41806 24498 41858
rect 25454 41806 25506 41858
rect 27806 41806 27858 41858
rect 28254 41806 28306 41858
rect 28814 41806 28866 41858
rect 30942 41806 30994 41858
rect 32286 41806 32338 41858
rect 35310 41806 35362 41858
rect 6638 41694 6690 41746
rect 6974 41694 7026 41746
rect 22430 41694 22482 41746
rect 23886 41694 23938 41746
rect 31502 41694 31554 41746
rect 31838 41694 31890 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 22654 41358 22706 41410
rect 29038 41358 29090 41410
rect 29486 41358 29538 41410
rect 29710 41358 29762 41410
rect 30158 41358 30210 41410
rect 30606 41358 30658 41410
rect 34974 41358 35026 41410
rect 36430 41358 36482 41410
rect 37438 41358 37490 41410
rect 7198 41246 7250 41298
rect 10782 41246 10834 41298
rect 12910 41246 12962 41298
rect 21422 41246 21474 41298
rect 22878 41246 22930 41298
rect 23326 41246 23378 41298
rect 25118 41246 25170 41298
rect 25902 41246 25954 41298
rect 27134 41246 27186 41298
rect 27470 41246 27522 41298
rect 28366 41246 28418 41298
rect 29262 41246 29314 41298
rect 29710 41246 29762 41298
rect 30158 41246 30210 41298
rect 30606 41246 30658 41298
rect 35310 41246 35362 41298
rect 36094 41246 36146 41298
rect 37102 41246 37154 41298
rect 6526 41134 6578 41186
rect 9998 41134 10050 41186
rect 14814 41134 14866 41186
rect 15038 41134 15090 41186
rect 18510 41134 18562 41186
rect 20750 41134 20802 41186
rect 21310 41134 21362 41186
rect 21534 41134 21586 41186
rect 24782 41134 24834 41186
rect 25454 41134 25506 41186
rect 25678 41134 25730 41186
rect 31502 41134 31554 41186
rect 38222 41134 38274 41186
rect 6750 41022 6802 41074
rect 15598 41032 15650 41084
rect 17502 41022 17554 41074
rect 20078 41022 20130 41074
rect 21982 41022 22034 41074
rect 23774 41022 23826 41074
rect 26574 41022 26626 41074
rect 35534 41022 35586 41074
rect 35870 41022 35922 41074
rect 13582 40910 13634 40962
rect 16494 40910 16546 40962
rect 17054 40910 17106 40962
rect 21758 40910 21810 40962
rect 22318 40910 22370 40962
rect 27918 40910 27970 40962
rect 31726 40910 31778 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 6974 40574 7026 40626
rect 13246 40574 13298 40626
rect 16382 40574 16434 40626
rect 16942 40574 16994 40626
rect 17502 40574 17554 40626
rect 22094 40574 22146 40626
rect 22878 40574 22930 40626
rect 23886 40574 23938 40626
rect 24222 40574 24274 40626
rect 24670 40574 24722 40626
rect 25902 40574 25954 40626
rect 26238 40574 26290 40626
rect 26574 40574 26626 40626
rect 27582 40574 27634 40626
rect 28478 40574 28530 40626
rect 29486 40574 29538 40626
rect 30494 40574 30546 40626
rect 35310 40574 35362 40626
rect 35758 40574 35810 40626
rect 38334 40574 38386 40626
rect 4958 40462 5010 40514
rect 5854 40462 5906 40514
rect 13582 40462 13634 40514
rect 14366 40462 14418 40514
rect 15150 40462 15202 40514
rect 17950 40462 18002 40514
rect 20414 40462 20466 40514
rect 20862 40462 20914 40514
rect 21198 40462 21250 40514
rect 29598 40462 29650 40514
rect 3950 40350 4002 40402
rect 4286 40350 4338 40402
rect 4510 40350 4562 40402
rect 5406 40350 5458 40402
rect 5630 40350 5682 40402
rect 5966 40350 6018 40402
rect 6526 40350 6578 40402
rect 9998 40350 10050 40402
rect 17390 40350 17442 40402
rect 19182 40350 19234 40402
rect 29150 40350 29202 40402
rect 30270 40350 30322 40402
rect 5742 40238 5794 40290
rect 10670 40238 10722 40290
rect 12798 40238 12850 40290
rect 15374 40238 15426 40290
rect 22542 40238 22594 40290
rect 23438 40238 23490 40290
rect 25342 40238 25394 40290
rect 27134 40238 27186 40290
rect 28030 40238 28082 40290
rect 37774 40238 37826 40290
rect 15710 40126 15762 40178
rect 23774 40126 23826 40178
rect 24782 40126 24834 40178
rect 25342 40126 25394 40178
rect 25790 40126 25842 40178
rect 26910 40126 26962 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 15598 39790 15650 39842
rect 19518 39790 19570 39842
rect 19966 39790 20018 39842
rect 22766 39790 22818 39842
rect 23774 39790 23826 39842
rect 24110 39790 24162 39842
rect 29822 39790 29874 39842
rect 33630 39790 33682 39842
rect 34078 39790 34130 39842
rect 34302 39790 34354 39842
rect 6190 39678 6242 39730
rect 6750 39678 6802 39730
rect 7198 39678 7250 39730
rect 18510 39678 18562 39730
rect 19966 39678 20018 39730
rect 20302 39678 20354 39730
rect 20862 39678 20914 39730
rect 22206 39678 22258 39730
rect 24446 39678 24498 39730
rect 29262 39678 29314 39730
rect 30382 39678 30434 39730
rect 32510 39678 32562 39730
rect 35758 39678 35810 39730
rect 37886 39678 37938 39730
rect 3166 39566 3218 39618
rect 4398 39566 4450 39618
rect 5070 39566 5122 39618
rect 5630 39566 5682 39618
rect 5854 39566 5906 39618
rect 12910 39566 12962 39618
rect 13806 39566 13858 39618
rect 15150 39566 15202 39618
rect 18174 39566 18226 39618
rect 21870 39566 21922 39618
rect 22654 39566 22706 39618
rect 26462 39566 26514 39618
rect 27022 39566 27074 39618
rect 33182 39566 33234 39618
rect 33742 39566 33794 39618
rect 34526 39566 34578 39618
rect 34974 39566 35026 39618
rect 35310 39566 35362 39618
rect 35870 39566 35922 39618
rect 36094 39566 36146 39618
rect 36206 39566 36258 39618
rect 37214 39566 37266 39618
rect 15038 39454 15090 39506
rect 17726 39454 17778 39506
rect 21646 39454 21698 39506
rect 23662 39454 23714 39506
rect 24334 39454 24386 39506
rect 24894 39454 24946 39506
rect 27470 39454 27522 39506
rect 29934 39454 29986 39506
rect 35198 39454 35250 39506
rect 2942 39342 2994 39394
rect 4622 39342 4674 39394
rect 4734 39342 4786 39394
rect 4846 39342 4898 39394
rect 6078 39342 6130 39394
rect 6190 39342 6242 39394
rect 12462 39342 12514 39394
rect 14030 39342 14082 39394
rect 14926 39342 14978 39394
rect 16382 39342 16434 39394
rect 18174 39342 18226 39394
rect 22094 39342 22146 39394
rect 22206 39342 22258 39394
rect 22766 39342 22818 39394
rect 23326 39342 23378 39394
rect 28478 39342 28530 39394
rect 35758 39342 35810 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 5182 39006 5234 39058
rect 5518 39006 5570 39058
rect 10446 39006 10498 39058
rect 13022 39006 13074 39058
rect 18398 39006 18450 39058
rect 22990 39006 23042 39058
rect 24110 39006 24162 39058
rect 24222 39006 24274 39058
rect 31390 39006 31442 39058
rect 33630 39006 33682 39058
rect 2494 38894 2546 38946
rect 5966 38894 6018 38946
rect 6302 38894 6354 38946
rect 6862 38894 6914 38946
rect 17390 38894 17442 38946
rect 17726 38894 17778 38946
rect 21646 38894 21698 38946
rect 23326 38894 23378 38946
rect 24334 38894 24386 38946
rect 25230 38894 25282 38946
rect 26014 38894 26066 38946
rect 30606 38894 30658 38946
rect 32398 38894 32450 38946
rect 1822 38782 1874 38834
rect 5854 38782 5906 38834
rect 6414 38782 6466 38834
rect 10110 38782 10162 38834
rect 16270 38782 16322 38834
rect 19182 38782 19234 38834
rect 22318 38770 22370 38822
rect 23998 38782 24050 38834
rect 24558 38782 24610 38834
rect 25790 38782 25842 38834
rect 26238 38782 26290 38834
rect 26462 38782 26514 38834
rect 27246 38782 27298 38834
rect 31838 38782 31890 38834
rect 32174 38782 32226 38834
rect 38110 38782 38162 38834
rect 4622 38670 4674 38722
rect 13358 38670 13410 38722
rect 15486 38670 15538 38722
rect 16830 38670 16882 38722
rect 18622 38670 18674 38722
rect 18958 38670 19010 38722
rect 19518 38670 19570 38722
rect 28030 38670 28082 38722
rect 30158 38670 30210 38722
rect 32510 38670 32562 38722
rect 33070 38670 33122 38722
rect 35310 38670 35362 38722
rect 37438 38670 37490 38722
rect 17950 38558 18002 38610
rect 18398 38558 18450 38610
rect 33294 38558 33346 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 26462 38222 26514 38274
rect 26910 38222 26962 38274
rect 4846 38110 4898 38162
rect 5742 38110 5794 38162
rect 7422 38110 7474 38162
rect 14814 38110 14866 38162
rect 15934 38110 15986 38162
rect 16382 38110 16434 38162
rect 18398 38110 18450 38162
rect 20526 38110 20578 38162
rect 22206 38110 22258 38162
rect 23102 38110 23154 38162
rect 25230 38110 25282 38162
rect 26462 38110 26514 38162
rect 30494 38110 30546 38162
rect 35534 38110 35586 38162
rect 38222 38110 38274 38162
rect 4622 37998 4674 38050
rect 10222 37998 10274 38050
rect 11454 37998 11506 38050
rect 14590 37998 14642 38050
rect 15822 37998 15874 38050
rect 17054 37998 17106 38050
rect 17726 37998 17778 38050
rect 22318 37998 22370 38050
rect 26014 37998 26066 38050
rect 33406 37998 33458 38050
rect 36430 37998 36482 38050
rect 37774 37998 37826 38050
rect 3278 37886 3330 37938
rect 9550 37886 9602 37938
rect 10670 37886 10722 37938
rect 11006 37886 11058 37938
rect 15374 37886 15426 37938
rect 16606 37886 16658 37938
rect 16830 37886 16882 37938
rect 21646 37886 21698 37938
rect 21870 37886 21922 37938
rect 32622 37886 32674 37938
rect 36990 37886 37042 37938
rect 37326 37886 37378 37938
rect 2942 37774 2994 37826
rect 4286 37774 4338 37826
rect 13918 37774 13970 37826
rect 14254 37774 14306 37826
rect 15598 37774 15650 37826
rect 15934 37774 15986 37826
rect 17390 37774 17442 37826
rect 22094 37774 22146 37826
rect 22766 37774 22818 37826
rect 26910 37774 26962 37826
rect 33854 37774 33906 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 5070 37438 5122 37490
rect 10110 37438 10162 37490
rect 10558 37438 10610 37490
rect 15374 37438 15426 37490
rect 15710 37438 15762 37490
rect 16606 37438 16658 37490
rect 18286 37438 18338 37490
rect 19518 37438 19570 37490
rect 20750 37438 20802 37490
rect 21870 37438 21922 37490
rect 23438 37438 23490 37490
rect 23886 37438 23938 37490
rect 24334 37438 24386 37490
rect 25790 37438 25842 37490
rect 28254 37438 28306 37490
rect 28926 37438 28978 37490
rect 2494 37326 2546 37378
rect 13470 37326 13522 37378
rect 13806 37326 13858 37378
rect 16046 37326 16098 37378
rect 22430 37326 22482 37378
rect 27806 37326 27858 37378
rect 28142 37326 28194 37378
rect 1822 37214 1874 37266
rect 5518 37214 5570 37266
rect 5630 37214 5682 37266
rect 5742 37214 5794 37266
rect 5966 37214 6018 37266
rect 9774 37214 9826 37266
rect 12574 37214 12626 37266
rect 22654 37214 22706 37266
rect 28478 37214 28530 37266
rect 38222 37214 38274 37266
rect 4622 37102 4674 37154
rect 6750 37102 6802 37154
rect 9550 37102 9602 37154
rect 11678 37102 11730 37154
rect 13022 37102 13074 37154
rect 17726 37102 17778 37154
rect 19966 37102 20018 37154
rect 20526 37102 20578 37154
rect 21310 37102 21362 37154
rect 25342 37102 25394 37154
rect 31614 37102 31666 37154
rect 35310 37102 35362 37154
rect 37438 37102 37490 37154
rect 6414 36990 6466 37042
rect 12014 36990 12066 37042
rect 12350 36990 12402 37042
rect 21086 36990 21138 37042
rect 22990 36990 23042 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 22654 36654 22706 36706
rect 23326 36654 23378 36706
rect 37550 36654 37602 36706
rect 5182 36542 5234 36594
rect 5966 36542 6018 36594
rect 6750 36542 6802 36594
rect 8542 36542 8594 36594
rect 15150 36542 15202 36594
rect 16606 36542 16658 36594
rect 17278 36542 17330 36594
rect 18510 36542 18562 36594
rect 22766 36542 22818 36594
rect 23102 36542 23154 36594
rect 28142 36542 28194 36594
rect 38222 36542 38274 36594
rect 5854 36430 5906 36482
rect 6078 36430 6130 36482
rect 8990 36430 9042 36482
rect 9102 36430 9154 36482
rect 9438 36430 9490 36482
rect 11678 36430 11730 36482
rect 23998 36430 24050 36482
rect 25230 36430 25282 36482
rect 29150 36430 29202 36482
rect 30158 36430 30210 36482
rect 31054 36430 31106 36482
rect 31838 36430 31890 36482
rect 36206 36430 36258 36482
rect 36990 36430 37042 36482
rect 37214 36430 37266 36482
rect 5630 36318 5682 36370
rect 9214 36318 9266 36370
rect 24334 36318 24386 36370
rect 26014 36318 26066 36370
rect 36430 36318 36482 36370
rect 6190 36206 6242 36258
rect 7198 36206 7250 36258
rect 9886 36206 9938 36258
rect 11454 36206 11506 36258
rect 21534 36206 21586 36258
rect 22206 36206 22258 36258
rect 23550 36206 23602 36258
rect 28590 36206 28642 36258
rect 30942 36206 30994 36258
rect 32846 36206 32898 36258
rect 35758 36206 35810 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 9774 35870 9826 35922
rect 9886 35870 9938 35922
rect 10670 35870 10722 35922
rect 15710 35870 15762 35922
rect 20526 35870 20578 35922
rect 20862 35870 20914 35922
rect 23326 35870 23378 35922
rect 28702 35870 28754 35922
rect 31054 35870 31106 35922
rect 31166 35870 31218 35922
rect 35086 35870 35138 35922
rect 36430 35870 36482 35922
rect 4174 35758 4226 35810
rect 7310 35758 7362 35810
rect 9550 35758 9602 35810
rect 12798 35758 12850 35810
rect 17502 35758 17554 35810
rect 17838 35758 17890 35810
rect 19742 35758 19794 35810
rect 19966 35758 20018 35810
rect 26686 35758 26738 35810
rect 28926 35758 28978 35810
rect 30606 35758 30658 35810
rect 3950 35646 4002 35698
rect 4510 35646 4562 35698
rect 4734 35646 4786 35698
rect 5518 35646 5570 35698
rect 6974 35646 7026 35698
rect 9998 35646 10050 35698
rect 10110 35646 10162 35698
rect 11118 35646 11170 35698
rect 12014 35646 12066 35698
rect 15598 35646 15650 35698
rect 15934 35646 15986 35698
rect 16158 35646 16210 35698
rect 17950 35646 18002 35698
rect 19518 35646 19570 35698
rect 20078 35646 20130 35698
rect 27022 35646 27074 35698
rect 28254 35646 28306 35698
rect 29150 35646 29202 35698
rect 30830 35646 30882 35698
rect 32398 35646 32450 35698
rect 6638 35534 6690 35586
rect 14926 35534 14978 35586
rect 15822 35534 15874 35586
rect 17390 35534 17442 35586
rect 18734 35534 18786 35586
rect 19294 35534 19346 35586
rect 30942 35534 30994 35586
rect 33182 35534 33234 35586
rect 35534 35534 35586 35586
rect 36094 35534 36146 35586
rect 36766 35534 36818 35586
rect 36990 35534 37042 35586
rect 3614 35422 3666 35474
rect 5070 35422 5122 35474
rect 10782 35422 10834 35474
rect 11230 35422 11282 35474
rect 18398 35422 18450 35474
rect 18622 35422 18674 35474
rect 19294 35422 19346 35474
rect 31838 35422 31890 35474
rect 32174 35422 32226 35474
rect 35534 35422 35586 35474
rect 36206 35422 36258 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 28478 35086 28530 35138
rect 4398 34974 4450 35026
rect 7534 34974 7586 35026
rect 9662 34974 9714 35026
rect 10782 34974 10834 35026
rect 12910 34974 12962 35026
rect 15374 34974 15426 35026
rect 19630 34974 19682 35026
rect 22206 34974 22258 35026
rect 34862 34974 34914 35026
rect 35646 34974 35698 35026
rect 3278 34862 3330 34914
rect 5854 34862 5906 34914
rect 5966 34862 6018 34914
rect 6302 34862 6354 34914
rect 6750 34862 6802 34914
rect 10110 34862 10162 34914
rect 15150 34862 15202 34914
rect 17838 34862 17890 34914
rect 18622 34862 18674 34914
rect 25118 34862 25170 34914
rect 25566 34862 25618 34914
rect 30270 34862 30322 34914
rect 31390 34862 31442 34914
rect 31950 34862 32002 34914
rect 35870 34862 35922 34914
rect 35982 34862 36034 34914
rect 18062 34750 18114 34802
rect 18174 34750 18226 34802
rect 24334 34750 24386 34802
rect 28590 34750 28642 34802
rect 31614 34750 31666 34802
rect 32734 34750 32786 34802
rect 35534 34750 35586 34802
rect 2942 34638 2994 34690
rect 6078 34638 6130 34690
rect 6190 34638 6242 34690
rect 13582 34638 13634 34690
rect 14814 34638 14866 34690
rect 15822 34638 15874 34690
rect 18846 34638 18898 34690
rect 19182 34638 19234 34690
rect 35646 34638 35698 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 6974 34302 7026 34354
rect 7422 34302 7474 34354
rect 17726 34302 17778 34354
rect 19630 34302 19682 34354
rect 22990 34302 23042 34354
rect 24558 34302 24610 34354
rect 27022 34302 27074 34354
rect 29374 34302 29426 34354
rect 31950 34302 32002 34354
rect 33406 34302 33458 34354
rect 33742 34302 33794 34354
rect 34078 34302 34130 34354
rect 34526 34302 34578 34354
rect 2494 34190 2546 34242
rect 4958 34190 5010 34242
rect 15038 34190 15090 34242
rect 15374 34190 15426 34242
rect 18622 34190 18674 34242
rect 27358 34190 27410 34242
rect 31054 34190 31106 34242
rect 31278 34190 31330 34242
rect 35198 34190 35250 34242
rect 35422 34190 35474 34242
rect 1822 34078 1874 34130
rect 5182 34078 5234 34130
rect 6078 34078 6130 34130
rect 6190 34078 6242 34130
rect 6302 34078 6354 34130
rect 6526 34078 6578 34130
rect 7758 34078 7810 34130
rect 13134 34078 13186 34130
rect 17390 34078 17442 34130
rect 17614 34078 17666 34130
rect 17838 34078 17890 34130
rect 17950 34078 18002 34130
rect 18846 34078 18898 34130
rect 19294 34078 19346 34130
rect 19518 34078 19570 34130
rect 19742 34078 19794 34130
rect 19854 34078 19906 34130
rect 23550 34078 23602 34130
rect 23886 34078 23938 34130
rect 24222 34078 24274 34130
rect 28478 34078 28530 34130
rect 29150 34078 29202 34130
rect 29486 34078 29538 34130
rect 31502 34078 31554 34130
rect 33854 34078 33906 34130
rect 34302 34078 34354 34130
rect 34750 34078 34802 34130
rect 4622 33966 4674 34018
rect 9886 33966 9938 34018
rect 12238 33966 12290 34018
rect 20974 33966 21026 34018
rect 23326 33966 23378 34018
rect 30942 33966 30994 34018
rect 33966 33966 34018 34018
rect 35534 33966 35586 34018
rect 12574 33854 12626 33906
rect 12910 33854 12962 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 4734 33518 4786 33570
rect 4958 33518 5010 33570
rect 6526 33518 6578 33570
rect 26350 33518 26402 33570
rect 26798 33518 26850 33570
rect 27022 33518 27074 33570
rect 27694 33518 27746 33570
rect 29262 33518 29314 33570
rect 33070 33518 33122 33570
rect 5966 33406 6018 33458
rect 7422 33406 7474 33458
rect 15262 33406 15314 33458
rect 17390 33406 17442 33458
rect 18622 33406 18674 33458
rect 20750 33406 20802 33458
rect 21870 33406 21922 33458
rect 26350 33406 26402 33458
rect 26798 33406 26850 33458
rect 31278 33406 31330 33458
rect 35310 33406 35362 33458
rect 6190 33294 6242 33346
rect 6974 33294 7026 33346
rect 12574 33294 12626 33346
rect 14590 33294 14642 33346
rect 17838 33294 17890 33346
rect 21646 33294 21698 33346
rect 27358 33294 27410 33346
rect 28030 33294 28082 33346
rect 31502 33294 31554 33346
rect 33294 33294 33346 33346
rect 33742 33294 33794 33346
rect 34078 33294 34130 33346
rect 34974 33294 35026 33346
rect 35534 33294 35586 33346
rect 28478 33182 28530 33234
rect 29150 33182 29202 33234
rect 32174 33182 32226 33234
rect 32510 33182 32562 33234
rect 33966 33182 34018 33234
rect 35870 33182 35922 33234
rect 36990 33182 37042 33234
rect 4846 33070 4898 33122
rect 12798 33070 12850 33122
rect 21310 33070 21362 33122
rect 24110 33070 24162 33122
rect 27134 33070 27186 33122
rect 27806 33070 27858 33122
rect 30942 33070 30994 33122
rect 31838 33070 31890 33122
rect 37326 33070 37378 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 16830 32734 16882 32786
rect 17502 32734 17554 32786
rect 18398 32734 18450 32786
rect 4622 32622 4674 32674
rect 8094 32622 8146 32674
rect 12574 32622 12626 32674
rect 21422 32622 21474 32674
rect 27582 32622 27634 32674
rect 33070 32622 33122 32674
rect 33406 32622 33458 32674
rect 37438 32622 37490 32674
rect 3950 32510 4002 32562
rect 7310 32510 7362 32562
rect 11790 32510 11842 32562
rect 15150 32510 15202 32562
rect 17838 32510 17890 32562
rect 21198 32510 21250 32562
rect 26910 32510 26962 32562
rect 38222 32510 38274 32562
rect 6750 32398 6802 32450
rect 7086 32398 7138 32450
rect 14702 32398 14754 32450
rect 29710 32398 29762 32450
rect 30158 32398 30210 32450
rect 35310 32398 35362 32450
rect 7646 32286 7698 32338
rect 18062 32286 18114 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 35870 31950 35922 32002
rect 10110 31838 10162 31890
rect 10558 31838 10610 31890
rect 15598 31838 15650 31890
rect 17614 31838 17666 31890
rect 21310 31838 21362 31890
rect 23438 31838 23490 31890
rect 26462 31838 26514 31890
rect 28590 31838 28642 31890
rect 29262 31838 29314 31890
rect 35422 31838 35474 31890
rect 35646 31838 35698 31890
rect 7310 31726 7362 31778
rect 15822 31726 15874 31778
rect 24222 31726 24274 31778
rect 24670 31726 24722 31778
rect 25678 31726 25730 31778
rect 7982 31614 8034 31666
rect 15262 31614 15314 31666
rect 36206 31614 36258 31666
rect 36990 31614 37042 31666
rect 16158 31502 16210 31554
rect 37326 31502 37378 31554
rect 38222 31502 38274 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 5742 31166 5794 31218
rect 7982 31166 8034 31218
rect 8990 31166 9042 31218
rect 24222 31166 24274 31218
rect 31950 31166 32002 31218
rect 7646 31054 7698 31106
rect 16270 31054 16322 31106
rect 16606 31054 16658 31106
rect 19966 31054 20018 31106
rect 33854 31054 33906 31106
rect 2494 30942 2546 30994
rect 9886 30942 9938 30994
rect 10110 30942 10162 30994
rect 19854 30942 19906 30994
rect 33182 30942 33234 30994
rect 3166 30830 3218 30882
rect 5294 30830 5346 30882
rect 19070 30830 19122 30882
rect 19518 30830 19570 30882
rect 22878 30830 22930 30882
rect 23214 30830 23266 30882
rect 30494 30830 30546 30882
rect 31278 30830 31330 30882
rect 32398 30830 32450 30882
rect 35982 30830 36034 30882
rect 36430 30830 36482 30882
rect 10446 30718 10498 30770
rect 19966 30718 20018 30770
rect 23438 30718 23490 30770
rect 23774 30718 23826 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 19406 30382 19458 30434
rect 31838 30382 31890 30434
rect 16718 30270 16770 30322
rect 18846 30270 18898 30322
rect 19182 30270 19234 30322
rect 4734 30158 4786 30210
rect 10670 30158 10722 30210
rect 12686 30158 12738 30210
rect 15934 30158 15986 30210
rect 22206 30158 22258 30210
rect 22430 30158 22482 30210
rect 24110 30158 24162 30210
rect 26910 30158 26962 30210
rect 31614 30158 31666 30210
rect 32174 30158 32226 30210
rect 32734 30158 32786 30210
rect 3502 30046 3554 30098
rect 3838 30046 3890 30098
rect 20078 30046 20130 30098
rect 29822 30046 29874 30098
rect 30494 30046 30546 30098
rect 30830 30046 30882 30098
rect 32510 30046 32562 30098
rect 32958 30046 33010 30098
rect 11006 29934 11058 29986
rect 12910 29934 12962 29986
rect 19742 29934 19794 29986
rect 20414 29934 20466 29986
rect 22766 29934 22818 29986
rect 23214 29934 23266 29986
rect 24446 29934 24498 29986
rect 30158 29934 30210 29986
rect 31054 29934 31106 29986
rect 31278 29934 31330 29986
rect 31390 29934 31442 29986
rect 33070 29934 33122 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 4958 29598 5010 29650
rect 9886 29598 9938 29650
rect 15710 29598 15762 29650
rect 16606 29598 16658 29650
rect 17502 29598 17554 29650
rect 23438 29598 23490 29650
rect 25902 29598 25954 29650
rect 27246 29598 27298 29650
rect 28142 29598 28194 29650
rect 33630 29598 33682 29650
rect 10782 29486 10834 29538
rect 13470 29486 13522 29538
rect 15486 29486 15538 29538
rect 20526 29486 20578 29538
rect 22430 29486 22482 29538
rect 22766 29486 22818 29538
rect 30382 29486 30434 29538
rect 37438 29486 37490 29538
rect 1710 29374 1762 29426
rect 5518 29374 5570 29426
rect 10558 29374 10610 29426
rect 14142 29374 14194 29426
rect 14702 29374 14754 29426
rect 15822 29374 15874 29426
rect 16270 29374 16322 29426
rect 21198 29374 21250 29426
rect 21758 29374 21810 29426
rect 24110 29374 24162 29426
rect 24334 29374 24386 29426
rect 26686 29374 26738 29426
rect 27022 29374 27074 29426
rect 29710 29374 29762 29426
rect 33070 29374 33122 29426
rect 38222 29374 38274 29426
rect 2494 29262 2546 29314
rect 4622 29262 4674 29314
rect 7086 29262 7138 29314
rect 11342 29262 11394 29314
rect 18398 29262 18450 29314
rect 26238 29262 26290 29314
rect 27358 29262 27410 29314
rect 27582 29262 27634 29314
rect 32510 29262 32562 29314
rect 35310 29262 35362 29314
rect 5294 29150 5346 29202
rect 10222 29150 10274 29202
rect 23774 29150 23826 29202
rect 27806 29150 27858 29202
rect 33294 29150 33346 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 13470 28814 13522 28866
rect 13806 28814 13858 28866
rect 19182 28814 19234 28866
rect 20302 28814 20354 28866
rect 27470 28814 27522 28866
rect 30382 28814 30434 28866
rect 30718 28814 30770 28866
rect 32398 28814 32450 28866
rect 4398 28702 4450 28754
rect 4846 28702 4898 28754
rect 6526 28702 6578 28754
rect 7310 28702 7362 28754
rect 9214 28702 9266 28754
rect 10782 28702 10834 28754
rect 12910 28702 12962 28754
rect 14030 28702 14082 28754
rect 17054 28702 17106 28754
rect 24782 28702 24834 28754
rect 26910 28702 26962 28754
rect 27246 28702 27298 28754
rect 30046 28702 30098 28754
rect 30942 28702 30994 28754
rect 31838 28702 31890 28754
rect 32846 28702 32898 28754
rect 3390 28590 3442 28642
rect 3838 28590 3890 28642
rect 4174 28590 4226 28642
rect 6302 28590 6354 28642
rect 6750 28590 6802 28642
rect 8206 28590 8258 28642
rect 10110 28590 10162 28642
rect 18622 28590 18674 28642
rect 23998 28590 24050 28642
rect 27806 28590 27858 28642
rect 28366 28590 28418 28642
rect 29262 28590 29314 28642
rect 32062 28590 32114 28642
rect 3054 28478 3106 28530
rect 6414 28478 6466 28530
rect 6638 28478 6690 28530
rect 7982 28478 8034 28530
rect 20190 28478 20242 28530
rect 20302 28366 20354 28418
rect 28142 28366 28194 28418
rect 38222 28366 38274 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 13246 28030 13298 28082
rect 13582 28030 13634 28082
rect 17614 28030 17666 28082
rect 17838 28030 17890 28082
rect 17950 28030 18002 28082
rect 18510 28030 18562 28082
rect 20526 28030 20578 28082
rect 25342 28030 25394 28082
rect 26798 28030 26850 28082
rect 30718 28030 30770 28082
rect 32622 28030 32674 28082
rect 36878 28030 36930 28082
rect 8206 27918 8258 27970
rect 16830 27918 16882 27970
rect 17726 27918 17778 27970
rect 22318 27918 22370 27970
rect 25566 27918 25618 27970
rect 28142 27918 28194 27970
rect 32062 27918 32114 27970
rect 32510 27918 32562 27970
rect 8990 27806 9042 27858
rect 9886 27806 9938 27858
rect 10558 27806 10610 27858
rect 16606 27806 16658 27858
rect 17390 27806 17442 27858
rect 20078 27806 20130 27858
rect 21646 27806 21698 27858
rect 25678 27806 25730 27858
rect 26350 27806 26402 27858
rect 26574 27806 26626 27858
rect 27470 27806 27522 27858
rect 32286 27806 32338 27858
rect 36990 27806 37042 27858
rect 4622 27694 4674 27746
rect 6078 27694 6130 27746
rect 10110 27694 10162 27746
rect 24446 27694 24498 27746
rect 26686 27694 26738 27746
rect 30270 27694 30322 27746
rect 31502 27694 31554 27746
rect 9550 27582 9602 27634
rect 30494 27582 30546 27634
rect 30830 27582 30882 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 5518 27246 5570 27298
rect 6078 27246 6130 27298
rect 29934 27246 29986 27298
rect 30718 27246 30770 27298
rect 31502 27246 31554 27298
rect 4734 27134 4786 27186
rect 5742 27134 5794 27186
rect 6302 27134 6354 27186
rect 13470 27134 13522 27186
rect 17726 27134 17778 27186
rect 19854 27134 19906 27186
rect 24670 27134 24722 27186
rect 26910 27134 26962 27186
rect 29934 27134 29986 27186
rect 31838 27134 31890 27186
rect 32398 27134 32450 27186
rect 36206 27134 36258 27186
rect 1822 27022 1874 27074
rect 9102 27022 9154 27074
rect 9662 27022 9714 27074
rect 16270 27022 16322 27074
rect 16942 27022 16994 27074
rect 20302 27022 20354 27074
rect 26462 27022 26514 27074
rect 30830 27022 30882 27074
rect 32062 27022 32114 27074
rect 2606 26910 2658 26962
rect 8430 26910 8482 26962
rect 15598 26910 15650 26962
rect 24222 26910 24274 26962
rect 25902 26910 25954 26962
rect 26350 26910 26402 26962
rect 30382 26910 30434 26962
rect 31390 26910 31442 26962
rect 32622 26910 32674 26962
rect 34974 26910 35026 26962
rect 35198 26910 35250 26962
rect 36990 26910 37042 26962
rect 38222 26910 38274 26962
rect 25454 26798 25506 26850
rect 31166 26798 31218 26850
rect 32398 26798 32450 26850
rect 37326 26798 37378 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 8318 26462 8370 26514
rect 15038 26462 15090 26514
rect 16830 26462 16882 26514
rect 17390 26462 17442 26514
rect 23438 26462 23490 26514
rect 24334 26462 24386 26514
rect 25902 26462 25954 26514
rect 26014 26462 26066 26514
rect 31726 26462 31778 26514
rect 32062 26462 32114 26514
rect 22094 26350 22146 26402
rect 22654 26350 22706 26402
rect 23774 26350 23826 26402
rect 37438 26350 37490 26402
rect 5406 26238 5458 26290
rect 8094 26238 8146 26290
rect 14814 26238 14866 26290
rect 15822 26238 15874 26290
rect 17950 26238 18002 26290
rect 22878 26238 22930 26290
rect 24782 26238 24834 26290
rect 25454 26238 25506 26290
rect 25678 26238 25730 26290
rect 38222 26238 38274 26290
rect 4510 26126 4562 26178
rect 15486 26126 15538 26178
rect 16382 26126 16434 26178
rect 22990 26126 23042 26178
rect 26350 26126 26402 26178
rect 35310 26126 35362 26178
rect 4846 26014 4898 26066
rect 5182 26014 5234 26066
rect 16158 26014 16210 26066
rect 17726 26014 17778 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 25230 25678 25282 25730
rect 36990 25678 37042 25730
rect 6190 25566 6242 25618
rect 6638 25566 6690 25618
rect 17054 25566 17106 25618
rect 25902 25566 25954 25618
rect 26350 25566 26402 25618
rect 37326 25566 37378 25618
rect 5966 25454 6018 25506
rect 22094 25454 22146 25506
rect 25118 25454 25170 25506
rect 3726 25342 3778 25394
rect 4062 25342 4114 25394
rect 12686 25342 12738 25394
rect 23550 25342 23602 25394
rect 24446 25342 24498 25394
rect 26126 25342 26178 25394
rect 27022 25342 27074 25394
rect 35422 25342 35474 25394
rect 36094 25342 36146 25394
rect 37550 25342 37602 25394
rect 37886 25342 37938 25394
rect 38222 25342 38274 25394
rect 5630 25230 5682 25282
rect 26686 25230 26738 25282
rect 27358 25230 27410 25282
rect 27806 25230 27858 25282
rect 30158 25230 30210 25282
rect 31054 25230 31106 25282
rect 31502 25230 31554 25282
rect 35758 25230 35810 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 14030 24894 14082 24946
rect 24670 24894 24722 24946
rect 25678 24894 25730 24946
rect 31166 24894 31218 24946
rect 3278 24782 3330 24834
rect 3614 24782 3666 24834
rect 3950 24782 4002 24834
rect 4286 24782 4338 24834
rect 27806 24782 27858 24834
rect 30270 24782 30322 24834
rect 31838 24782 31890 24834
rect 33406 24782 33458 24834
rect 35758 24782 35810 24834
rect 9662 24670 9714 24722
rect 13022 24670 13074 24722
rect 21422 24670 21474 24722
rect 27022 24670 27074 24722
rect 31390 24670 31442 24722
rect 32062 24670 32114 24722
rect 33070 24670 33122 24722
rect 34974 24670 35026 24722
rect 10334 24558 10386 24610
rect 12462 24558 12514 24610
rect 22094 24558 22146 24610
rect 24222 24558 24274 24610
rect 29934 24558 29986 24610
rect 30830 24558 30882 24610
rect 32398 24558 32450 24610
rect 34638 24558 34690 24610
rect 37886 24558 37938 24610
rect 13246 24446 13298 24498
rect 13582 24446 13634 24498
rect 30494 24446 30546 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 5630 24110 5682 24162
rect 12798 24110 12850 24162
rect 19630 24110 19682 24162
rect 16942 23998 16994 24050
rect 26126 23998 26178 24050
rect 32622 23998 32674 24050
rect 32958 23998 33010 24050
rect 35086 23998 35138 24050
rect 38334 23998 38386 24050
rect 5966 23886 6018 23938
rect 6190 23886 6242 23938
rect 9774 23886 9826 23938
rect 13582 23886 13634 23938
rect 16270 23886 16322 23938
rect 18510 23886 18562 23938
rect 21870 23886 21922 23938
rect 25566 23886 25618 23938
rect 25902 23886 25954 23938
rect 29710 23886 29762 23938
rect 35758 23886 35810 23938
rect 9998 23774 10050 23826
rect 12686 23774 12738 23826
rect 16382 23774 16434 23826
rect 18286 23774 18338 23826
rect 19518 23774 19570 23826
rect 20414 23774 20466 23826
rect 20750 23774 20802 23826
rect 25230 23774 25282 23826
rect 27918 23774 27970 23826
rect 30494 23774 30546 23826
rect 5070 23662 5122 23714
rect 9214 23662 9266 23714
rect 12350 23662 12402 23714
rect 12798 23662 12850 23714
rect 13918 23662 13970 23714
rect 18846 23662 18898 23714
rect 19630 23662 19682 23714
rect 22094 23662 22146 23714
rect 27582 23662 27634 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 5518 23326 5570 23378
rect 6750 23326 6802 23378
rect 8654 23326 8706 23378
rect 10110 23326 10162 23378
rect 10558 23326 10610 23378
rect 16718 23326 16770 23378
rect 19070 23326 19122 23378
rect 19966 23326 20018 23378
rect 29262 23326 29314 23378
rect 33182 23326 33234 23378
rect 33630 23326 33682 23378
rect 34750 23326 34802 23378
rect 34862 23326 34914 23378
rect 36094 23326 36146 23378
rect 2606 23214 2658 23266
rect 11566 23214 11618 23266
rect 14142 23214 14194 23266
rect 22654 23214 22706 23266
rect 24670 23214 24722 23266
rect 27358 23214 27410 23266
rect 28590 23214 28642 23266
rect 1822 23102 1874 23154
rect 5294 23102 5346 23154
rect 5406 23102 5458 23154
rect 5630 23102 5682 23154
rect 5854 23102 5906 23154
rect 6302 23102 6354 23154
rect 8318 23102 8370 23154
rect 8542 23102 8594 23154
rect 8766 23102 8818 23154
rect 8878 23102 8930 23154
rect 9774 23102 9826 23154
rect 11790 23102 11842 23154
rect 13470 23102 13522 23154
rect 17950 23102 18002 23154
rect 23438 23102 23490 23154
rect 24446 23102 24498 23154
rect 28030 23102 28082 23154
rect 29822 23102 29874 23154
rect 34526 23102 34578 23154
rect 34974 23102 35026 23154
rect 35198 23102 35250 23154
rect 35534 23102 35586 23154
rect 4734 22990 4786 23042
rect 9550 22990 9602 23042
rect 11006 22990 11058 23042
rect 12350 22990 12402 23042
rect 16270 22990 16322 23042
rect 17614 22990 17666 23042
rect 18174 22990 18226 23042
rect 20526 22990 20578 23042
rect 23886 22990 23938 23042
rect 25230 22990 25282 23042
rect 34078 22990 34130 23042
rect 18510 22878 18562 22930
rect 29598 22878 29650 22930
rect 33742 22878 33794 22930
rect 34302 22878 34354 22930
rect 35758 22878 35810 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 11790 22542 11842 22594
rect 21870 22542 21922 22594
rect 2494 22430 2546 22482
rect 4622 22430 4674 22482
rect 5070 22430 5122 22482
rect 6302 22430 6354 22482
rect 6862 22430 6914 22482
rect 7310 22430 7362 22482
rect 11454 22430 11506 22482
rect 12350 22430 12402 22482
rect 12798 22430 12850 22482
rect 15598 22430 15650 22482
rect 16382 22430 16434 22482
rect 21534 22430 21586 22482
rect 22206 22430 22258 22482
rect 25006 22430 25058 22482
rect 27134 22430 27186 22482
rect 27694 22430 27746 22482
rect 32734 22430 32786 22482
rect 1822 22318 1874 22370
rect 5966 22318 6018 22370
rect 8654 22318 8706 22370
rect 12126 22318 12178 22370
rect 14926 22318 14978 22370
rect 15262 22318 15314 22370
rect 15934 22318 15986 22370
rect 19182 22318 19234 22370
rect 19966 22318 20018 22370
rect 20414 22318 20466 22370
rect 22430 22318 22482 22370
rect 24222 22318 24274 22370
rect 5742 22206 5794 22258
rect 9326 22206 9378 22258
rect 18510 22206 18562 22258
rect 19630 22206 19682 22258
rect 6190 22094 6242 22146
rect 6302 22094 6354 22146
rect 15486 22094 15538 22146
rect 15710 22094 15762 22146
rect 29262 22094 29314 22146
rect 34190 22094 34242 22146
rect 35198 22094 35250 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 9550 21758 9602 21810
rect 15934 21758 15986 21810
rect 16046 21758 16098 21810
rect 16158 21758 16210 21810
rect 16830 21758 16882 21810
rect 21422 21758 21474 21810
rect 4734 21646 4786 21698
rect 11566 21646 11618 21698
rect 21982 21646 22034 21698
rect 5294 21534 5346 21586
rect 5966 21534 6018 21586
rect 9774 21534 9826 21586
rect 10894 21534 10946 21586
rect 14142 21534 14194 21586
rect 15710 21534 15762 21586
rect 16382 21534 16434 21586
rect 17390 21534 17442 21586
rect 32510 21534 32562 21586
rect 34526 21534 34578 21586
rect 37774 21534 37826 21586
rect 4398 21422 4450 21474
rect 6750 21422 6802 21474
rect 8878 21422 8930 21474
rect 13694 21422 13746 21474
rect 18174 21422 18226 21474
rect 20302 21422 20354 21474
rect 21086 21422 21138 21474
rect 29598 21422 29650 21474
rect 31726 21422 31778 21474
rect 33630 21422 33682 21474
rect 34862 21422 34914 21474
rect 36990 21422 37042 21474
rect 5070 21310 5122 21362
rect 21758 21310 21810 21362
rect 33070 21310 33122 21362
rect 33406 21310 33458 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 8990 20974 9042 21026
rect 5742 20862 5794 20914
rect 9550 20862 9602 20914
rect 16382 20862 16434 20914
rect 16830 20862 16882 20914
rect 17726 20862 17778 20914
rect 18286 20862 18338 20914
rect 20526 20862 20578 20914
rect 21534 20862 21586 20914
rect 27022 20862 27074 20914
rect 34974 20862 35026 20914
rect 4174 20750 4226 20802
rect 5070 20750 5122 20802
rect 5966 20750 6018 20802
rect 7422 20750 7474 20802
rect 8430 20750 8482 20802
rect 8654 20750 8706 20802
rect 17390 20750 17442 20802
rect 27246 20750 27298 20802
rect 31838 20750 31890 20802
rect 35870 20750 35922 20802
rect 6302 20638 6354 20690
rect 6638 20638 6690 20690
rect 6974 20638 7026 20690
rect 31502 20638 31554 20690
rect 36094 20638 36146 20690
rect 3838 20526 3890 20578
rect 8094 20526 8146 20578
rect 26686 20526 26738 20578
rect 27582 20526 27634 20578
rect 32734 20526 32786 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 18174 20190 18226 20242
rect 3278 20078 3330 20130
rect 20638 20078 20690 20130
rect 20974 20078 21026 20130
rect 24558 20078 24610 20130
rect 27806 20078 27858 20130
rect 28142 20078 28194 20130
rect 34638 20078 34690 20130
rect 2606 19966 2658 20018
rect 12014 19966 12066 20018
rect 17838 19966 17890 20018
rect 23886 19966 23938 20018
rect 24110 19966 24162 20018
rect 34414 19966 34466 20018
rect 34526 19966 34578 20018
rect 34750 19966 34802 20018
rect 34974 19966 35026 20018
rect 38110 19966 38162 20018
rect 5406 19854 5458 19906
rect 5966 19854 6018 19906
rect 11118 19854 11170 19906
rect 23214 19854 23266 19906
rect 33294 19854 33346 19906
rect 33742 19854 33794 19906
rect 35310 19854 35362 19906
rect 37438 19854 37490 19906
rect 11454 19742 11506 19794
rect 11790 19742 11842 19794
rect 23550 19742 23602 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 4174 19406 4226 19458
rect 36094 19406 36146 19458
rect 4398 19294 4450 19346
rect 14254 19294 14306 19346
rect 16382 19294 16434 19346
rect 17278 19294 17330 19346
rect 23774 19294 23826 19346
rect 29262 19294 29314 19346
rect 29710 19294 29762 19346
rect 30718 19294 30770 19346
rect 32398 19294 32450 19346
rect 32846 19294 32898 19346
rect 33966 19294 34018 19346
rect 35534 19294 35586 19346
rect 13470 19182 13522 19234
rect 16830 19182 16882 19234
rect 17166 19182 17218 19234
rect 23214 19182 23266 19234
rect 26686 19182 26738 19234
rect 30382 19182 30434 19234
rect 30494 19182 30546 19234
rect 30830 19182 30882 19234
rect 33630 19182 33682 19234
rect 34078 19182 34130 19234
rect 34862 19182 34914 19234
rect 35758 19182 35810 19234
rect 25902 19070 25954 19122
rect 33406 19070 33458 19122
rect 34638 19070 34690 19122
rect 36990 19070 37042 19122
rect 37326 19070 37378 19122
rect 3838 18958 3890 19010
rect 4846 18958 4898 19010
rect 17166 18958 17218 19010
rect 23438 18958 23490 19010
rect 27134 18958 27186 19010
rect 30718 18958 30770 19010
rect 31390 18958 31442 19010
rect 33854 18958 33906 19010
rect 35198 18958 35250 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 17726 18622 17778 18674
rect 34302 18622 34354 18674
rect 9550 18510 9602 18562
rect 10334 18510 10386 18562
rect 10670 18510 10722 18562
rect 19854 18510 19906 18562
rect 19966 18510 20018 18562
rect 28366 18510 28418 18562
rect 31726 18510 31778 18562
rect 33742 18510 33794 18562
rect 2270 18398 2322 18450
rect 9886 18398 9938 18450
rect 16830 18398 16882 18450
rect 20414 18398 20466 18450
rect 27694 18398 27746 18450
rect 31054 18398 31106 18450
rect 32062 18398 32114 18450
rect 33518 18398 33570 18450
rect 38110 18398 38162 18450
rect 2942 18286 2994 18338
rect 5070 18286 5122 18338
rect 5518 18286 5570 18338
rect 18286 18286 18338 18338
rect 20974 18286 21026 18338
rect 30494 18286 30546 18338
rect 30830 18286 30882 18338
rect 31390 18286 31442 18338
rect 32510 18286 32562 18338
rect 34974 18286 35026 18338
rect 35310 18286 35362 18338
rect 37438 18286 37490 18338
rect 5294 18174 5346 18226
rect 5630 18174 5682 18226
rect 18062 18174 18114 18226
rect 19854 18174 19906 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 5854 17838 5906 17890
rect 33630 17838 33682 17890
rect 5070 17726 5122 17778
rect 5630 17726 5682 17778
rect 7982 17726 8034 17778
rect 10110 17726 10162 17778
rect 17838 17726 17890 17778
rect 19966 17726 20018 17778
rect 23438 17726 23490 17778
rect 25566 17726 25618 17778
rect 30046 17726 30098 17778
rect 31166 17726 31218 17778
rect 33294 17726 33346 17778
rect 34190 17726 34242 17778
rect 3614 17614 3666 17666
rect 6190 17614 6242 17666
rect 6750 17614 6802 17666
rect 10782 17614 10834 17666
rect 13694 17614 13746 17666
rect 20750 17614 20802 17666
rect 22654 17614 22706 17666
rect 26126 17614 26178 17666
rect 30494 17614 30546 17666
rect 33966 17614 34018 17666
rect 35086 17614 35138 17666
rect 3278 17502 3330 17554
rect 14478 17502 14530 17554
rect 21310 17502 21362 17554
rect 25902 17502 25954 17554
rect 34638 17502 34690 17554
rect 6526 17390 6578 17442
rect 11342 17390 11394 17442
rect 13470 17390 13522 17442
rect 14142 17390 14194 17442
rect 14926 17390 14978 17442
rect 21646 17390 21698 17442
rect 26686 17390 26738 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 8654 17054 8706 17106
rect 15038 17054 15090 17106
rect 16270 17054 16322 17106
rect 17502 17054 17554 17106
rect 25902 17054 25954 17106
rect 26910 17054 26962 17106
rect 29262 17054 29314 17106
rect 32510 17054 32562 17106
rect 36654 17054 36706 17106
rect 6078 16942 6130 16994
rect 12574 16942 12626 16994
rect 17950 16942 18002 16994
rect 21870 16942 21922 16994
rect 23102 16942 23154 16994
rect 33854 16942 33906 16994
rect 5406 16830 5458 16882
rect 11790 16830 11842 16882
rect 15598 16830 15650 16882
rect 16158 16830 16210 16882
rect 16494 16830 16546 16882
rect 16718 16830 16770 16882
rect 22654 16830 22706 16882
rect 26238 16830 26290 16882
rect 33182 16830 33234 16882
rect 36318 16830 36370 16882
rect 8206 16718 8258 16770
rect 14702 16718 14754 16770
rect 16382 16718 16434 16770
rect 19070 16718 19122 16770
rect 19742 16718 19794 16770
rect 26462 16718 26514 16770
rect 28814 16718 28866 16770
rect 35982 16718 36034 16770
rect 15374 16606 15426 16658
rect 28814 16606 28866 16658
rect 29374 16606 29426 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 13470 16270 13522 16322
rect 22094 16270 22146 16322
rect 29486 16270 29538 16322
rect 35534 16270 35586 16322
rect 9326 16158 9378 16210
rect 11454 16158 11506 16210
rect 12910 16158 12962 16210
rect 13806 16158 13858 16210
rect 15934 16158 15986 16210
rect 21870 16158 21922 16210
rect 22878 16158 22930 16210
rect 23438 16158 23490 16210
rect 25678 16158 25730 16210
rect 34974 16158 35026 16210
rect 8654 16046 8706 16098
rect 12014 16046 12066 16098
rect 12462 16046 12514 16098
rect 14030 16046 14082 16098
rect 14478 16046 14530 16098
rect 18734 16046 18786 16098
rect 19294 16046 19346 16098
rect 20750 16046 20802 16098
rect 21422 16046 21474 16098
rect 28590 16046 28642 16098
rect 29710 16046 29762 16098
rect 35198 16046 35250 16098
rect 11790 15934 11842 15986
rect 18062 15934 18114 15986
rect 19406 15934 19458 15986
rect 20526 15934 20578 15986
rect 27806 15934 27858 15986
rect 12126 15822 12178 15874
rect 12238 15822 12290 15874
rect 14926 15822 14978 15874
rect 20414 15822 20466 15874
rect 22430 15822 22482 15874
rect 29150 15822 29202 15874
rect 34638 15822 34690 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 7534 15486 7586 15538
rect 8990 15486 9042 15538
rect 11678 15486 11730 15538
rect 12686 15486 12738 15538
rect 16494 15486 16546 15538
rect 17278 15486 17330 15538
rect 18958 15486 19010 15538
rect 21310 15486 21362 15538
rect 23102 15486 23154 15538
rect 23886 15486 23938 15538
rect 23998 15486 24050 15538
rect 25342 15486 25394 15538
rect 26238 15486 26290 15538
rect 27358 15486 27410 15538
rect 28702 15486 28754 15538
rect 32286 15486 32338 15538
rect 13918 15374 13970 15426
rect 17838 15374 17890 15426
rect 18174 15374 18226 15426
rect 19294 15374 19346 15426
rect 19630 15374 19682 15426
rect 22654 15374 22706 15426
rect 24222 15374 24274 15426
rect 26462 15374 26514 15426
rect 6862 15262 6914 15314
rect 7086 15262 7138 15314
rect 10222 15262 10274 15314
rect 10446 15262 10498 15314
rect 13134 15262 13186 15314
rect 17502 15262 17554 15314
rect 19742 15262 19794 15314
rect 20302 15262 20354 15314
rect 21646 15262 21698 15314
rect 22430 15262 22482 15314
rect 24110 15262 24162 15314
rect 24446 15262 24498 15314
rect 26014 15262 26066 15314
rect 26686 15262 26738 15314
rect 27134 15262 27186 15314
rect 29038 15262 29090 15314
rect 16046 15150 16098 15202
rect 18286 15150 18338 15202
rect 19406 15150 19458 15202
rect 21870 15150 21922 15202
rect 26350 15150 26402 15202
rect 29710 15150 29762 15202
rect 31838 15150 31890 15202
rect 6526 15038 6578 15090
rect 9886 15038 9938 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 25902 14702 25954 14754
rect 26350 14702 26402 14754
rect 27358 14702 27410 14754
rect 14702 14590 14754 14642
rect 18958 14590 19010 14642
rect 22542 14590 22594 14642
rect 24670 14590 24722 14642
rect 25454 14590 25506 14642
rect 25902 14590 25954 14642
rect 26462 14590 26514 14642
rect 30606 14590 30658 14642
rect 30942 14590 30994 14642
rect 31166 14590 31218 14642
rect 34750 14590 34802 14642
rect 6302 14478 6354 14530
rect 14478 14478 14530 14530
rect 17502 14478 17554 14530
rect 21870 14478 21922 14530
rect 26798 14478 26850 14530
rect 27022 14478 27074 14530
rect 29262 14478 29314 14530
rect 31950 14478 32002 14530
rect 17726 14366 17778 14418
rect 29598 14366 29650 14418
rect 32622 14366 32674 14418
rect 5966 14254 6018 14306
rect 14142 14254 14194 14306
rect 15150 14254 15202 14306
rect 31502 14254 31554 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 17614 13918 17666 13970
rect 33070 13918 33122 13970
rect 5406 13806 5458 13858
rect 9550 13806 9602 13858
rect 9886 13806 9938 13858
rect 4734 13694 4786 13746
rect 7982 13694 8034 13746
rect 33294 13694 33346 13746
rect 7534 13582 7586 13634
rect 17950 13582 18002 13634
rect 18174 13582 18226 13634
rect 18622 13582 18674 13634
rect 25342 13582 25394 13634
rect 31502 13582 31554 13634
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 24558 13134 24610 13186
rect 31166 13134 31218 13186
rect 7198 13022 7250 13074
rect 8318 13022 8370 13074
rect 10446 13022 10498 13074
rect 17054 13022 17106 13074
rect 17502 13022 17554 13074
rect 18286 13022 18338 13074
rect 24782 13022 24834 13074
rect 25230 13022 25282 13074
rect 30270 13022 30322 13074
rect 7646 12910 7698 12962
rect 13806 12910 13858 12962
rect 30718 12910 30770 12962
rect 10894 12686 10946 12738
rect 13470 12686 13522 12738
rect 18958 12686 19010 12738
rect 24222 12686 24274 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 6638 12350 6690 12402
rect 8094 12350 8146 12402
rect 12238 12350 12290 12402
rect 13358 12350 13410 12402
rect 13806 12350 13858 12402
rect 15038 12350 15090 12402
rect 15486 12350 15538 12402
rect 16158 12350 16210 12402
rect 17278 12350 17330 12402
rect 18846 12350 18898 12402
rect 6302 12238 6354 12290
rect 12014 12238 12066 12290
rect 19070 12238 19122 12290
rect 24222 12238 24274 12290
rect 6078 12126 6130 12178
rect 6974 12126 7026 12178
rect 8430 12126 8482 12178
rect 9886 12126 9938 12178
rect 12462 12126 12514 12178
rect 12686 12126 12738 12178
rect 15934 12126 15986 12178
rect 16270 12126 16322 12178
rect 16382 12126 16434 12178
rect 16606 12126 16658 12178
rect 17502 12126 17554 12178
rect 17950 12126 18002 12178
rect 18062 12126 18114 12178
rect 18622 12126 18674 12178
rect 19294 12126 19346 12178
rect 23774 12126 23826 12178
rect 29710 12126 29762 12178
rect 7198 12014 7250 12066
rect 7646 12014 7698 12066
rect 8990 12014 9042 12066
rect 10110 12014 10162 12066
rect 12350 12014 12402 12066
rect 18286 12014 18338 12066
rect 18958 12014 19010 12066
rect 19742 12014 19794 12066
rect 20862 12014 20914 12066
rect 22990 12014 23042 12066
rect 26798 12014 26850 12066
rect 28926 12014 28978 12066
rect 30158 12014 30210 12066
rect 9550 11902 9602 11954
rect 29934 11902 29986 11954
rect 30158 11902 30210 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 14478 11566 14530 11618
rect 6974 11454 7026 11506
rect 12014 11454 12066 11506
rect 12910 11454 12962 11506
rect 14814 11454 14866 11506
rect 18734 11454 18786 11506
rect 19182 11454 19234 11506
rect 20750 11454 20802 11506
rect 25902 11454 25954 11506
rect 26350 11454 26402 11506
rect 27134 11454 27186 11506
rect 30270 11454 30322 11506
rect 5630 11342 5682 11394
rect 9102 11342 9154 11394
rect 15374 11342 15426 11394
rect 15822 11342 15874 11394
rect 19630 11342 19682 11394
rect 20190 11342 20242 11394
rect 21422 11342 21474 11394
rect 21758 11342 21810 11394
rect 22318 11342 22370 11394
rect 24334 11342 24386 11394
rect 33070 11342 33122 11394
rect 9886 11230 9938 11282
rect 14254 11230 14306 11282
rect 16606 11230 16658 11282
rect 19742 11230 19794 11282
rect 19966 11230 20018 11282
rect 21310 11230 21362 11282
rect 21646 11230 21698 11282
rect 22542 11230 22594 11282
rect 27694 11230 27746 11282
rect 28030 11230 28082 11282
rect 32398 11230 32450 11282
rect 12462 11118 12514 11170
rect 15150 11118 15202 11170
rect 24110 11118 24162 11170
rect 29934 11118 29986 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 8990 10782 9042 10834
rect 9886 10782 9938 10834
rect 10670 10782 10722 10834
rect 10782 10782 10834 10834
rect 11342 10782 11394 10834
rect 11790 10782 11842 10834
rect 16158 10782 16210 10834
rect 17838 10782 17890 10834
rect 20638 10782 20690 10834
rect 21534 10782 21586 10834
rect 22430 10782 22482 10834
rect 22878 10782 22930 10834
rect 24222 10782 24274 10834
rect 25342 10782 25394 10834
rect 25454 10782 25506 10834
rect 26798 10782 26850 10834
rect 27470 10782 27522 10834
rect 31390 10782 31442 10834
rect 5294 10670 5346 10722
rect 6414 10670 6466 10722
rect 9550 10670 9602 10722
rect 12910 10670 12962 10722
rect 19742 10670 19794 10722
rect 20526 10670 20578 10722
rect 5742 10558 5794 10610
rect 10222 10558 10274 10610
rect 10446 10558 10498 10610
rect 12126 10558 12178 10610
rect 15822 10558 15874 10610
rect 18062 10558 18114 10610
rect 18510 10558 18562 10610
rect 18622 10558 18674 10610
rect 18846 10558 18898 10610
rect 19294 10558 19346 10610
rect 19630 10558 19682 10610
rect 19966 10558 20018 10610
rect 20190 10558 20242 10610
rect 20750 10558 20802 10610
rect 20974 10558 21026 10610
rect 22094 10558 22146 10610
rect 24670 10558 24722 10610
rect 25678 10558 25730 10610
rect 25790 10558 25842 10610
rect 26462 10558 26514 10610
rect 26686 10558 26738 10610
rect 26910 10558 26962 10610
rect 27134 10558 27186 10610
rect 31166 10558 31218 10610
rect 4286 10446 4338 10498
rect 8542 10446 8594 10498
rect 10670 10446 10722 10498
rect 15038 10446 15090 10498
rect 17502 10446 17554 10498
rect 21870 10446 21922 10498
rect 25342 10446 25394 10498
rect 28030 10446 28082 10498
rect 11342 10334 11394 10386
rect 11566 10334 11618 10386
rect 27806 10334 27858 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 11342 9998 11394 10050
rect 12014 9998 12066 10050
rect 27246 9998 27298 10050
rect 28030 9998 28082 10050
rect 31166 9998 31218 10050
rect 4734 9886 4786 9938
rect 11006 9886 11058 9938
rect 11566 9886 11618 9938
rect 12014 9886 12066 9938
rect 14254 9886 14306 9938
rect 16382 9886 16434 9938
rect 16830 9886 16882 9938
rect 17614 9886 17666 9938
rect 18286 9886 18338 9938
rect 18958 9886 19010 9938
rect 19406 9886 19458 9938
rect 19854 9886 19906 9938
rect 20078 9886 20130 9938
rect 23886 9886 23938 9938
rect 26014 9886 26066 9938
rect 26462 9886 26514 9938
rect 27470 9886 27522 9938
rect 27918 9886 27970 9938
rect 30046 9886 30098 9938
rect 31726 9886 31778 9938
rect 5630 9774 5682 9826
rect 10446 9774 10498 9826
rect 10670 9774 10722 9826
rect 11118 9774 11170 9826
rect 13470 9774 13522 9826
rect 17166 9774 17218 9826
rect 17726 9774 17778 9826
rect 20302 9774 20354 9826
rect 23102 9774 23154 9826
rect 26350 9774 26402 9826
rect 26798 9774 26850 9826
rect 29710 9774 29762 9826
rect 31502 9774 31554 9826
rect 32174 9774 32226 9826
rect 5070 9662 5122 9714
rect 7422 9662 7474 9714
rect 27022 9662 27074 9714
rect 30830 9662 30882 9714
rect 10894 9550 10946 9602
rect 17390 9550 17442 9602
rect 17614 9550 17666 9602
rect 20638 9550 20690 9602
rect 26574 9550 26626 9602
rect 28366 9550 28418 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 8990 9214 9042 9266
rect 15710 9214 15762 9266
rect 18174 9214 18226 9266
rect 20526 9102 20578 9154
rect 9886 8990 9938 9042
rect 10110 8990 10162 9042
rect 15486 8990 15538 9042
rect 16830 8990 16882 9042
rect 20302 8990 20354 9042
rect 25454 8990 25506 9042
rect 31950 8990 32002 9042
rect 32510 8990 32562 9042
rect 38222 8990 38274 9042
rect 5294 8878 5346 8930
rect 16270 8878 16322 8930
rect 19742 8878 19794 8930
rect 26126 8878 26178 8930
rect 28254 8878 28306 8930
rect 28702 8878 28754 8930
rect 29150 8878 29202 8930
rect 31278 8878 31330 8930
rect 37214 8878 37266 8930
rect 9550 8766 9602 8818
rect 16606 8766 16658 8818
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 29934 8430 29986 8482
rect 26126 8318 26178 8370
rect 27582 8318 27634 8370
rect 38334 8318 38386 8370
rect 8878 8206 8930 8258
rect 25566 8206 25618 8258
rect 26350 8206 26402 8258
rect 27022 8206 27074 8258
rect 27358 8206 27410 8258
rect 29598 8206 29650 8258
rect 31278 8206 31330 8258
rect 31502 8206 31554 8258
rect 25790 8094 25842 8146
rect 8542 7982 8594 8034
rect 15934 7982 15986 8034
rect 25118 7982 25170 8034
rect 26686 7982 26738 8034
rect 28030 7982 28082 8034
rect 30942 7982 30994 8034
rect 31950 7982 32002 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 10670 7646 10722 7698
rect 14478 7646 14530 7698
rect 30830 7646 30882 7698
rect 31390 7646 31442 7698
rect 10222 7534 10274 7586
rect 21198 7534 21250 7586
rect 26910 7534 26962 7586
rect 28030 7534 28082 7586
rect 5966 7422 6018 7474
rect 9998 7422 10050 7474
rect 11118 7422 11170 7474
rect 21982 7422 22034 7474
rect 26686 7422 26738 7474
rect 27246 7422 27298 7474
rect 30606 7422 30658 7474
rect 6638 7310 6690 7362
rect 7422 7310 7474 7362
rect 11902 7310 11954 7362
rect 14030 7310 14082 7362
rect 19070 7310 19122 7362
rect 22430 7310 22482 7362
rect 30158 7310 30210 7362
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 10782 6862 10834 6914
rect 12126 6862 12178 6914
rect 14366 6862 14418 6914
rect 10110 6750 10162 6802
rect 11006 6750 11058 6802
rect 11454 6750 11506 6802
rect 13694 6750 13746 6802
rect 14590 6750 14642 6802
rect 17838 6750 17890 6802
rect 7310 6638 7362 6690
rect 7982 6638 8034 6690
rect 10446 6638 10498 6690
rect 12350 6638 12402 6690
rect 15038 6638 15090 6690
rect 18286 6638 18338 6690
rect 23550 6638 23602 6690
rect 30382 6638 30434 6690
rect 15710 6526 15762 6578
rect 11790 6414 11842 6466
rect 14030 6414 14082 6466
rect 21870 6414 21922 6466
rect 22318 6414 22370 6466
rect 24894 6414 24946 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 16270 6078 16322 6130
rect 17390 5966 17442 6018
rect 9662 5854 9714 5906
rect 13022 5854 13074 5906
rect 17614 5854 17666 5906
rect 18958 5854 19010 5906
rect 22206 5854 22258 5906
rect 24222 5854 24274 5906
rect 24446 5854 24498 5906
rect 25566 5854 25618 5906
rect 25790 5854 25842 5906
rect 10334 5742 10386 5794
rect 12462 5742 12514 5794
rect 13694 5742 13746 5794
rect 15822 5742 15874 5794
rect 19630 5742 19682 5794
rect 21758 5742 21810 5794
rect 23214 5742 23266 5794
rect 23886 5630 23938 5682
rect 25230 5630 25282 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 20414 5294 20466 5346
rect 21534 5294 21586 5346
rect 9326 5182 9378 5234
rect 10110 5182 10162 5234
rect 12798 5182 12850 5234
rect 15934 5182 15986 5234
rect 17054 5182 17106 5234
rect 19182 5182 19234 5234
rect 19742 5182 19794 5234
rect 20638 5182 20690 5234
rect 21310 5182 21362 5234
rect 23102 5182 23154 5234
rect 27022 5182 27074 5234
rect 8654 5070 8706 5122
rect 12126 5070 12178 5122
rect 14478 5070 14530 5122
rect 15038 5070 15090 5122
rect 15710 5070 15762 5122
rect 16382 5070 16434 5122
rect 21870 5070 21922 5122
rect 22430 5070 22482 5122
rect 23550 5070 23602 5122
rect 24222 5070 24274 5122
rect 8318 4958 8370 5010
rect 14254 4958 14306 5010
rect 24894 4958 24946 5010
rect 27470 4958 27522 5010
rect 7982 4846 8034 4898
rect 8766 4846 8818 4898
rect 8990 4846 9042 4898
rect 11902 4846 11954 4898
rect 14030 4846 14082 4898
rect 15374 4846 15426 4898
rect 20078 4846 20130 4898
rect 22206 4846 22258 4898
rect 23774 4846 23826 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 8990 4510 9042 4562
rect 9774 4510 9826 4562
rect 11342 4510 11394 4562
rect 15822 4510 15874 4562
rect 16830 4510 16882 4562
rect 17390 4510 17442 4562
rect 19070 4510 19122 4562
rect 19630 4510 19682 4562
rect 23326 4510 23378 4562
rect 24670 4510 24722 4562
rect 7758 4398 7810 4450
rect 10222 4398 10274 4450
rect 10894 4398 10946 4450
rect 14030 4398 14082 4450
rect 22094 4398 22146 4450
rect 25230 4398 25282 4450
rect 25566 4398 25618 4450
rect 8542 4286 8594 4338
rect 10110 4286 10162 4338
rect 10446 4286 10498 4338
rect 10782 4286 10834 4338
rect 14590 4286 14642 4338
rect 16046 4286 16098 4338
rect 17726 4286 17778 4338
rect 17950 4286 18002 4338
rect 19406 4286 19458 4338
rect 22878 4286 22930 4338
rect 24446 4286 24498 4338
rect 25902 4286 25954 4338
rect 34414 4286 34466 4338
rect 34750 4286 34802 4338
rect 5630 4174 5682 4226
rect 15038 4174 15090 4226
rect 15486 4174 15538 4226
rect 18398 4174 18450 4226
rect 19966 4174 20018 4226
rect 26462 4174 26514 4226
rect 34526 4174 34578 4226
rect 33966 4062 34018 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 8094 3614 8146 3666
rect 10446 3614 10498 3666
rect 12574 3614 12626 3666
rect 23886 3614 23938 3666
rect 26014 3614 26066 3666
rect 26574 3614 26626 3666
rect 8318 3502 8370 3554
rect 8542 3502 8594 3554
rect 10110 3502 10162 3554
rect 10334 3502 10386 3554
rect 14814 3502 14866 3554
rect 15486 3502 15538 3554
rect 16046 3502 16098 3554
rect 18174 3502 18226 3554
rect 23214 3502 23266 3554
rect 27470 3502 27522 3554
rect 27918 3502 27970 3554
rect 31054 3502 31106 3554
rect 33182 3502 33234 3554
rect 6190 3390 6242 3442
rect 6302 3390 6354 3442
rect 7422 3390 7474 3442
rect 11118 3390 11170 3442
rect 13694 3390 13746 3442
rect 13918 3390 13970 3442
rect 14254 3390 14306 3442
rect 15038 3390 15090 3442
rect 15710 3390 15762 3442
rect 17166 3390 17218 3442
rect 18622 3390 18674 3442
rect 26910 3390 26962 3442
rect 28478 3390 28530 3442
rect 31166 3390 31218 3442
rect 33630 3390 33682 3442
rect 11454 3278 11506 3330
rect 12126 3278 12178 3330
rect 16158 3278 16210 3330
rect 20862 3278 20914 3330
rect 22654 3278 22706 3330
rect 27022 3278 27074 3330
rect 33070 3278 33122 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 10558 2942 10610 2994
rect 13694 2942 13746 2994
rect 17390 2942 17442 2994
rect 19854 2942 19906 2994
rect 25902 2942 25954 2994
rect 6414 2830 6466 2882
rect 10110 2830 10162 2882
rect 11566 2830 11618 2882
rect 12798 2830 12850 2882
rect 15262 2830 15314 2882
rect 20302 2830 20354 2882
rect 22318 2830 22370 2882
rect 25342 2830 25394 2882
rect 26798 2830 26850 2882
rect 33966 2830 34018 2882
rect 4622 2718 4674 2770
rect 10558 2718 10610 2770
rect 11118 2718 11170 2770
rect 12686 2718 12738 2770
rect 14814 2718 14866 2770
rect 17614 2718 17666 2770
rect 18174 2718 18226 2770
rect 19742 2718 19794 2770
rect 21870 2718 21922 2770
rect 25230 2718 25282 2770
rect 26350 2718 26402 2770
rect 33070 2718 33122 2770
rect 34750 2718 34802 2770
rect 7646 2606 7698 2658
rect 8542 2606 8594 2658
rect 9102 2606 9154 2658
rect 9774 2606 9826 2658
rect 12462 2606 12514 2658
rect 19070 2606 19122 2658
rect 19518 2606 19570 2658
rect 24334 2606 24386 2658
rect 24782 2606 24834 2658
rect 27358 2606 27410 2658
rect 27806 2606 27858 2658
rect 28366 2606 28418 2658
rect 28926 2606 28978 2658
rect 29822 2606 29874 2658
rect 30718 2606 30770 2658
rect 31950 2606 32002 2658
rect 32622 2606 32674 2658
rect 36094 2606 36146 2658
rect 36542 2606 36594 2658
rect 33182 2494 33234 2546
rect 4478 2326 4530 2378
rect 4582 2326 4634 2378
rect 4686 2326 4738 2378
rect 35198 2326 35250 2378
rect 35302 2326 35354 2378
rect 35406 2326 35458 2378
rect 13246 2158 13298 2210
rect 8542 1934 8594 1986
rect 10446 1934 10498 1986
rect 11230 1934 11282 1986
rect 11678 1934 11730 1986
rect 12350 1934 12402 1986
rect 13470 1934 13522 1986
rect 16270 1934 16322 1986
rect 17614 1934 17666 1986
rect 21086 1934 21138 1986
rect 21982 1934 22034 1986
rect 22878 1934 22930 1986
rect 23662 1934 23714 1986
rect 26014 1934 26066 1986
rect 27582 1934 27634 1986
rect 29374 1934 29426 1986
rect 32174 1934 32226 1986
rect 33742 1934 33794 1986
rect 34862 1934 34914 1986
rect 35310 1934 35362 1986
rect 36206 1934 36258 1986
rect 36878 1934 36930 1986
rect 3838 1822 3890 1874
rect 4062 1822 4114 1874
rect 4398 1822 4450 1874
rect 5854 1822 5906 1874
rect 6190 1822 6242 1874
rect 7086 1822 7138 1874
rect 7646 1822 7698 1874
rect 7982 1822 8034 1874
rect 8766 1822 8818 1874
rect 9438 1822 9490 1874
rect 9774 1822 9826 1874
rect 10222 1822 10274 1874
rect 10894 1822 10946 1874
rect 11902 1822 11954 1874
rect 12574 1822 12626 1874
rect 13694 1822 13746 1874
rect 14926 1822 14978 1874
rect 17838 1822 17890 1874
rect 18398 1822 18450 1874
rect 18734 1822 18786 1874
rect 19182 1822 19234 1874
rect 19518 1822 19570 1874
rect 19854 1822 19906 1874
rect 20190 1822 20242 1874
rect 21422 1822 21474 1874
rect 22318 1822 22370 1874
rect 23214 1822 23266 1874
rect 24558 1822 24610 1874
rect 24894 1822 24946 1874
rect 25230 1822 25282 1874
rect 25566 1822 25618 1874
rect 26238 1822 26290 1874
rect 26574 1822 26626 1874
rect 27358 1822 27410 1874
rect 28366 1822 28418 1874
rect 28702 1822 28754 1874
rect 30046 1822 30098 1874
rect 30382 1822 30434 1874
rect 30942 1822 30994 1874
rect 31278 1822 31330 1874
rect 32510 1822 32562 1874
rect 32846 1822 32898 1874
rect 33182 1822 33234 1874
rect 34526 1822 34578 1874
rect 35982 1822 36034 1874
rect 36654 1822 36706 1874
rect 3390 1710 3442 1762
rect 5070 1710 5122 1762
rect 6750 1710 6802 1762
rect 17278 1710 17330 1762
rect 26910 1710 26962 1762
rect 29150 1710 29202 1762
rect 33966 1710 34018 1762
rect 37438 1710 37490 1762
rect 19838 1542 19890 1594
rect 19942 1542 19994 1594
rect 20046 1542 20098 1594
<< metal2 >>
rect 1344 99600 1456 100000
rect 3808 99600 3920 100000
rect 6272 99600 6384 100000
rect 8736 99600 8848 100000
rect 8988 99708 9380 99764
rect 1372 97524 1428 99600
rect 3836 97524 3892 99600
rect 4476 98028 4740 98038
rect 4532 97972 4580 98028
rect 4636 97972 4684 98028
rect 4476 97962 4740 97972
rect 6300 97524 6356 99600
rect 8764 99540 8820 99600
rect 8988 99540 9044 99708
rect 8764 99484 9044 99540
rect 1372 97468 1652 97524
rect 3836 97468 4116 97524
rect 6300 97468 6580 97524
rect 1596 97412 1652 97468
rect 1708 97412 1764 97422
rect 1596 97410 1764 97412
rect 1596 97358 1710 97410
rect 1762 97358 1764 97410
rect 1596 97356 1764 97358
rect 1708 97346 1764 97356
rect 4060 97410 4116 97468
rect 4060 97358 4062 97410
rect 4114 97358 4116 97410
rect 4060 97346 4116 97358
rect 6524 97410 6580 97468
rect 6524 97358 6526 97410
rect 6578 97358 6580 97410
rect 6524 97346 6580 97358
rect 9324 97410 9380 99708
rect 11200 99600 11312 100000
rect 13664 99600 13776 100000
rect 16128 99600 16240 100000
rect 18592 99600 18704 100000
rect 21056 99600 21168 100000
rect 23520 99600 23632 100000
rect 25984 99600 26096 100000
rect 28448 99600 28560 100000
rect 30912 99600 31024 100000
rect 33376 99600 33488 100000
rect 35840 99600 35952 100000
rect 38304 99600 38416 100000
rect 11228 97524 11284 99600
rect 13020 97524 13076 97534
rect 11228 97468 11508 97524
rect 9324 97358 9326 97410
rect 9378 97358 9380 97410
rect 9324 97346 9380 97358
rect 11452 97410 11508 97468
rect 13020 97430 13076 97468
rect 11452 97358 11454 97410
rect 11506 97358 11508 97410
rect 11452 97346 11508 97358
rect 13692 97412 13748 99600
rect 13692 97346 13748 97356
rect 14476 97634 14532 97646
rect 14476 97582 14478 97634
rect 14530 97582 14532 97634
rect 14476 97524 14532 97582
rect 7980 96852 8036 96862
rect 7644 96850 8372 96852
rect 7644 96798 7982 96850
rect 8034 96798 8372 96850
rect 7644 96796 8372 96798
rect 6188 96628 6244 96638
rect 4476 96460 4740 96470
rect 4532 96404 4580 96460
rect 4636 96404 4684 96460
rect 4476 96394 4740 96404
rect 2940 96066 2996 96078
rect 2940 96014 2942 96066
rect 2994 96014 2996 96066
rect 2940 94498 2996 96014
rect 2940 94446 2942 94498
rect 2994 94446 2996 94498
rect 1708 94388 1764 94398
rect 1708 94294 1764 94332
rect 2940 93716 2996 94446
rect 3836 96066 3892 96078
rect 3836 96014 3838 96066
rect 3890 96014 3892 96066
rect 3836 94498 3892 96014
rect 5180 95844 5236 95854
rect 5740 95844 5796 95854
rect 6188 95844 6244 96572
rect 6860 96628 6916 96638
rect 6860 96534 6916 96572
rect 7644 96628 7700 96796
rect 7980 96786 8036 96796
rect 4844 95842 6244 95844
rect 4844 95790 5182 95842
rect 5234 95790 5742 95842
rect 5794 95790 6244 95842
rect 4844 95788 6244 95790
rect 3836 94446 3838 94498
rect 3890 94446 3892 94498
rect 2044 93492 2100 93502
rect 2044 93398 2100 93436
rect 2940 92930 2996 93660
rect 3388 93716 3444 93726
rect 3836 93716 3892 94446
rect 3388 93714 3892 93716
rect 3388 93662 3390 93714
rect 3442 93662 3892 93714
rect 3388 93660 3892 93662
rect 3948 95282 4004 95294
rect 3948 95230 3950 95282
rect 4002 95230 4004 95282
rect 3948 93716 4004 95230
rect 4844 95284 4900 95788
rect 5180 95778 5236 95788
rect 4844 95282 5012 95284
rect 4844 95230 4846 95282
rect 4898 95230 5012 95282
rect 4844 95228 5012 95230
rect 4844 95218 4900 95228
rect 4476 94892 4740 94902
rect 4532 94836 4580 94892
rect 4636 94836 4684 94892
rect 4476 94826 4740 94836
rect 4956 94724 5012 95228
rect 4620 94722 5012 94724
rect 4620 94670 4958 94722
rect 5010 94670 5012 94722
rect 4620 94668 5012 94670
rect 4620 93938 4676 94668
rect 4620 93886 4622 93938
rect 4674 93886 4676 93938
rect 4620 93874 4676 93886
rect 4172 93716 4228 93726
rect 3948 93660 4172 93716
rect 3388 93492 3444 93660
rect 3388 93426 3444 93436
rect 2940 92878 2942 92930
rect 2994 92878 2996 92930
rect 2940 92146 2996 92878
rect 2940 92094 2942 92146
rect 2994 92094 2996 92146
rect 2940 91362 2996 92094
rect 2940 91310 2942 91362
rect 2994 91310 2996 91362
rect 2940 90748 2996 91310
rect 3836 92930 3892 93660
rect 4172 93622 4228 93660
rect 4476 93324 4740 93334
rect 4532 93268 4580 93324
rect 4636 93268 4684 93324
rect 4476 93258 4740 93268
rect 3836 92878 3838 92930
rect 3890 92878 3892 92930
rect 3836 92148 3892 92878
rect 4956 93154 5012 94668
rect 4956 93102 4958 93154
rect 5010 93102 5012 93154
rect 4844 92260 4900 92270
rect 4956 92260 5012 93102
rect 5740 94610 5796 95788
rect 6188 95508 6244 95788
rect 6748 96068 6804 96078
rect 6188 95506 6356 95508
rect 6188 95454 6190 95506
rect 6242 95454 6356 95506
rect 6188 95452 6356 95454
rect 6188 95442 6244 95452
rect 5740 94558 5742 94610
rect 5794 94558 5796 94610
rect 5740 93044 5796 94558
rect 6300 94610 6356 95452
rect 6300 94558 6302 94610
rect 6354 94558 6356 94610
rect 6300 94546 6356 94558
rect 6748 95282 6804 96012
rect 6748 95230 6750 95282
rect 6802 95230 6804 95282
rect 6748 93716 6804 95230
rect 7644 96066 7700 96572
rect 7644 96014 7646 96066
rect 7698 96014 7700 96066
rect 7644 95282 7700 96014
rect 8316 95956 8372 96796
rect 8876 96850 8932 96862
rect 8876 96798 8878 96850
rect 8930 96798 8932 96850
rect 8876 96068 8932 96798
rect 13916 96850 13972 96862
rect 13916 96798 13918 96850
rect 13970 96798 13972 96850
rect 9660 96738 9716 96750
rect 9660 96686 9662 96738
rect 9714 96686 9716 96738
rect 8876 96002 8932 96012
rect 9324 96068 9380 96078
rect 9324 95974 9380 96012
rect 8652 95956 8708 95966
rect 8316 95954 8708 95956
rect 8316 95902 8654 95954
rect 8706 95902 8708 95954
rect 8316 95900 8708 95902
rect 8652 95844 8708 95900
rect 8652 95778 8708 95788
rect 9660 95844 9716 96686
rect 10108 96738 10164 96750
rect 10108 96686 10110 96738
rect 10162 96686 10164 96738
rect 10108 96068 10164 96686
rect 12348 96738 12404 96750
rect 12348 96686 12350 96738
rect 12402 96686 12404 96738
rect 10332 96068 10388 96078
rect 10108 96066 10388 96068
rect 10108 96014 10334 96066
rect 10386 96014 10388 96066
rect 10108 96012 10388 96014
rect 9660 95508 9716 95788
rect 10332 95844 10388 96012
rect 10332 95778 10388 95788
rect 11676 95844 11732 95854
rect 12012 95844 12068 95854
rect 12348 95844 12404 96686
rect 11732 95842 12404 95844
rect 11732 95790 12014 95842
rect 12066 95790 12404 95842
rect 11732 95788 12404 95790
rect 11676 95750 11732 95788
rect 12012 95778 12068 95788
rect 7644 95230 7646 95282
rect 7698 95230 7700 95282
rect 7644 93716 7700 95230
rect 9324 95506 9716 95508
rect 9324 95454 9662 95506
rect 9714 95454 9716 95506
rect 9324 95452 9716 95454
rect 9100 95172 9156 95182
rect 9324 95172 9380 95452
rect 9660 95442 9716 95452
rect 12348 95508 12404 95788
rect 13580 96066 13636 96078
rect 13580 96014 13582 96066
rect 13634 96014 13636 96066
rect 13580 95732 13636 96014
rect 13580 95666 13636 95676
rect 12348 95414 12404 95452
rect 13916 95508 13972 96798
rect 13916 95282 13972 95452
rect 14476 96066 14532 97468
rect 15260 97634 15316 97646
rect 15260 97582 15262 97634
rect 15314 97582 15316 97634
rect 15260 96964 15316 97582
rect 15708 97412 15764 97422
rect 15708 97318 15764 97356
rect 16156 97412 16212 99600
rect 18620 97524 18676 99600
rect 18620 97468 18900 97524
rect 21084 97468 21140 99600
rect 16156 97346 16212 97356
rect 16268 97410 16324 97422
rect 16268 97358 16270 97410
rect 16322 97358 16324 97410
rect 15036 96908 15316 96964
rect 14476 96014 14478 96066
rect 14530 96014 14532 96066
rect 14476 95508 14532 96014
rect 14476 95442 14532 95452
rect 14700 96852 14756 96862
rect 15036 96852 15092 96908
rect 14700 96850 15092 96852
rect 14700 96798 14702 96850
rect 14754 96798 15092 96850
rect 14700 96796 15092 96798
rect 14700 95732 14756 96796
rect 13916 95230 13918 95282
rect 13970 95230 13972 95282
rect 13916 95218 13972 95230
rect 14700 95282 14756 95676
rect 15148 96740 15204 96750
rect 15148 96738 15652 96740
rect 15148 96686 15150 96738
rect 15202 96686 15652 96738
rect 15148 96684 15652 96686
rect 15148 95508 15204 96684
rect 15596 96292 15652 96684
rect 16268 96292 16324 97358
rect 16940 97412 16996 97422
rect 16940 97318 16996 97356
rect 18844 97410 18900 97468
rect 18844 97358 18846 97410
rect 18898 97358 18900 97410
rect 18844 97346 18900 97358
rect 20860 97412 21140 97468
rect 19836 97244 20100 97254
rect 19892 97188 19940 97244
rect 19996 97188 20044 97244
rect 19836 97178 20100 97188
rect 15596 96290 16324 96292
rect 15596 96238 15598 96290
rect 15650 96238 16324 96290
rect 15596 96236 16324 96238
rect 15596 96226 15652 96236
rect 16156 96178 16212 96236
rect 16156 96126 16158 96178
rect 16210 96126 16212 96178
rect 16156 96114 16212 96126
rect 16268 95732 16324 96236
rect 19516 96290 19572 96302
rect 19516 96238 19518 96290
rect 19570 96238 19572 96290
rect 16268 95666 16324 95676
rect 17500 96066 17556 96078
rect 17500 96014 17502 96066
rect 17554 96014 17556 96066
rect 14700 95230 14702 95282
rect 14754 95230 14756 95282
rect 9100 95170 9380 95172
rect 9100 95118 9102 95170
rect 9154 95118 9380 95170
rect 9100 95116 9380 95118
rect 9100 95106 9156 95116
rect 9100 93940 9156 93950
rect 9324 93940 9380 95116
rect 14700 94724 14756 95230
rect 14700 94658 14756 94668
rect 14812 95452 15148 95508
rect 9100 93938 9380 93940
rect 9100 93886 9102 93938
rect 9154 93886 9380 93938
rect 9100 93884 9380 93886
rect 9100 93874 9156 93884
rect 6804 93660 7028 93716
rect 6748 93622 6804 93660
rect 5628 93042 5796 93044
rect 5628 92990 5742 93042
rect 5794 92990 5796 93042
rect 5628 92988 5796 92990
rect 5628 92370 5684 92988
rect 5740 92978 5796 92988
rect 6972 92930 7028 93660
rect 7644 93714 7812 93716
rect 7644 93662 7646 93714
rect 7698 93662 7812 93714
rect 7644 93660 7812 93662
rect 7644 93650 7700 93660
rect 6972 92878 6974 92930
rect 7026 92878 7028 92930
rect 5628 92318 5630 92370
rect 5682 92318 5684 92370
rect 5628 92306 5684 92318
rect 6524 92596 6580 92606
rect 4844 92258 5012 92260
rect 4844 92206 4846 92258
rect 4898 92206 5012 92258
rect 4844 92204 5012 92206
rect 4844 92194 4900 92204
rect 3836 91362 3892 92092
rect 4956 92148 5012 92204
rect 4476 91756 4740 91766
rect 4532 91700 4580 91756
rect 4636 91700 4684 91756
rect 4476 91690 4740 91700
rect 4956 91586 5012 92092
rect 6524 92146 6580 92540
rect 6972 92596 7028 92878
rect 6972 92530 7028 92540
rect 7756 92930 7812 93660
rect 9324 93044 9380 93884
rect 13244 93828 13300 93838
rect 12124 93826 13300 93828
rect 12124 93774 13246 93826
rect 13298 93774 13300 93826
rect 12124 93772 13300 93774
rect 10332 93716 10388 93726
rect 7756 92878 7758 92930
rect 7810 92878 7812 92930
rect 6524 92094 6526 92146
rect 6578 92094 6580 92146
rect 6524 92082 6580 92094
rect 7308 92484 7364 92494
rect 7308 92146 7364 92428
rect 7756 92484 7812 92878
rect 7756 92418 7812 92428
rect 8876 93042 9380 93044
rect 8876 92990 9326 93042
rect 9378 92990 9380 93042
rect 8876 92988 9380 92990
rect 8764 92372 8820 92382
rect 8876 92372 8932 92988
rect 9324 92978 9380 92988
rect 9660 93602 9716 93614
rect 9660 93550 9662 93602
rect 9714 93550 9716 93602
rect 9660 92820 9716 93550
rect 9660 92484 9716 92764
rect 10332 92818 10388 93660
rect 12012 93716 12068 93726
rect 12012 93622 12068 93660
rect 10332 92766 10334 92818
rect 10386 92766 10388 92818
rect 10332 92754 10388 92766
rect 10780 93154 10836 93166
rect 10780 93102 10782 93154
rect 10834 93102 10836 93154
rect 10780 92820 10836 93102
rect 12124 92930 12180 93772
rect 13244 93762 13300 93772
rect 13356 93716 13412 93726
rect 13356 93622 13412 93660
rect 14140 93716 14196 93726
rect 12684 93604 12740 93614
rect 12684 93510 12740 93548
rect 12124 92878 12126 92930
rect 12178 92878 12180 92930
rect 12124 92866 12180 92878
rect 12348 93490 12404 93502
rect 12348 93438 12350 93490
rect 12402 93438 12404 93490
rect 10836 92764 11060 92820
rect 10780 92754 10836 92764
rect 9660 92418 9716 92428
rect 10780 92596 10836 92606
rect 8764 92370 8932 92372
rect 8764 92318 8766 92370
rect 8818 92318 8932 92370
rect 8764 92316 8932 92318
rect 8764 92306 8820 92316
rect 7308 92094 7310 92146
rect 7362 92094 7364 92146
rect 7308 92082 7364 92094
rect 4956 91534 4958 91586
rect 5010 91534 5012 91586
rect 4956 91522 5012 91534
rect 8876 91474 8932 92316
rect 10780 92370 10836 92540
rect 10780 92318 10782 92370
rect 10834 92318 10836 92370
rect 10780 92306 10836 92318
rect 9996 92260 10052 92270
rect 10220 92260 10276 92270
rect 9996 92258 10220 92260
rect 9996 92206 9998 92258
rect 10050 92206 10220 92258
rect 9996 92204 10220 92206
rect 9996 92194 10052 92204
rect 10220 92166 10276 92204
rect 10892 92148 10948 92158
rect 10780 92146 10948 92148
rect 10780 92094 10894 92146
rect 10946 92094 10948 92146
rect 10780 92092 10948 92094
rect 10332 91924 10388 91934
rect 10780 91924 10836 92092
rect 10892 92082 10948 92092
rect 10332 91922 10836 91924
rect 10332 91870 10334 91922
rect 10386 91870 10836 91922
rect 10332 91868 10836 91870
rect 10332 91858 10388 91868
rect 8876 91422 8878 91474
rect 8930 91422 8932 91474
rect 8876 91410 8932 91422
rect 3836 91310 3838 91362
rect 3890 91310 3892 91362
rect 2940 90692 3220 90748
rect 3164 90578 3220 90692
rect 3164 90526 3166 90578
rect 3218 90526 3220 90578
rect 3164 89796 3220 90526
rect 3836 90578 3892 91310
rect 3836 90526 3838 90578
rect 3890 90526 3892 90578
rect 3388 89796 3444 89806
rect 3836 89796 3892 90526
rect 5740 91138 5796 91150
rect 5740 91086 5742 91138
rect 5794 91086 5796 91138
rect 5740 90466 5796 91086
rect 11004 90748 11060 92764
rect 12348 92372 12404 93438
rect 12908 92932 12964 92942
rect 12908 92930 13524 92932
rect 12908 92878 12910 92930
rect 12962 92878 13524 92930
rect 12908 92876 13524 92878
rect 12908 92866 12964 92876
rect 12236 92316 12404 92372
rect 12572 92820 12628 92830
rect 12236 91586 12292 92316
rect 12348 92148 12404 92158
rect 12348 92054 12404 92092
rect 12236 91534 12238 91586
rect 12290 91534 12292 91586
rect 11564 91364 11620 91374
rect 11564 91270 11620 91308
rect 12012 91364 12068 91374
rect 12012 91270 12068 91308
rect 5740 90414 5742 90466
rect 5794 90414 5796 90466
rect 5180 90354 5236 90366
rect 5180 90302 5182 90354
rect 5234 90302 5236 90354
rect 4476 90188 4740 90198
rect 4532 90132 4580 90188
rect 4636 90132 4684 90188
rect 4476 90122 4740 90132
rect 3164 89730 3220 89740
rect 3276 89794 3892 89796
rect 3276 89742 3390 89794
rect 3442 89742 3892 89794
rect 3276 89740 3892 89742
rect 4284 89796 4340 89806
rect 2044 89572 2100 89582
rect 2044 89570 2212 89572
rect 2044 89518 2046 89570
rect 2098 89518 2212 89570
rect 2044 89516 2212 89518
rect 2044 89506 2100 89516
rect 2156 88450 2212 89516
rect 2156 88398 2158 88450
rect 2210 88398 2212 88450
rect 2156 87218 2212 88398
rect 2156 87166 2158 87218
rect 2210 87166 2212 87218
rect 2156 86882 2212 87166
rect 2156 86830 2158 86882
rect 2210 86830 2212 86882
rect 2156 85650 2212 86830
rect 2156 85598 2158 85650
rect 2210 85598 2212 85650
rect 2156 85314 2212 85598
rect 2156 85262 2158 85314
rect 2210 85262 2212 85314
rect 2156 84082 2212 85262
rect 2156 84030 2158 84082
rect 2210 84030 2212 84082
rect 2156 83748 2212 84030
rect 3276 88226 3332 89740
rect 3388 89730 3444 89740
rect 4284 89702 4340 89740
rect 4844 89572 4900 89582
rect 5180 89572 5236 90302
rect 5740 89572 5796 90414
rect 10780 90692 11060 90748
rect 11676 91138 11732 91150
rect 11676 91086 11678 91138
rect 11730 91086 11732 91138
rect 11676 90692 11732 91086
rect 10780 89906 10836 90692
rect 11676 90626 11732 90636
rect 12236 90356 12292 91534
rect 12572 91586 12628 92764
rect 13468 92818 13524 92876
rect 13468 92766 13470 92818
rect 13522 92766 13524 92818
rect 13468 92754 13524 92766
rect 13804 92820 13860 92830
rect 13804 92726 13860 92764
rect 14140 92818 14196 93660
rect 14588 93604 14644 93614
rect 14140 92766 14142 92818
rect 14194 92766 14196 92818
rect 14140 92754 14196 92766
rect 14252 93044 14308 93054
rect 13580 92372 13636 92382
rect 13468 92316 13580 92372
rect 12908 92260 12964 92270
rect 12572 91534 12574 91586
rect 12626 91534 12628 91586
rect 12572 91522 12628 91534
rect 12684 92146 12740 92158
rect 12684 92094 12686 92146
rect 12738 92094 12740 92146
rect 12572 90804 12628 90814
rect 12684 90804 12740 92094
rect 12572 90802 12740 90804
rect 12572 90750 12574 90802
rect 12626 90750 12740 90802
rect 12572 90748 12740 90750
rect 12572 90738 12628 90748
rect 12348 90692 12404 90702
rect 12348 90578 12404 90636
rect 12348 90526 12350 90578
rect 12402 90526 12404 90578
rect 12348 90514 12404 90526
rect 12684 90356 12740 90366
rect 12236 90354 12740 90356
rect 12236 90302 12686 90354
rect 12738 90302 12740 90354
rect 12236 90300 12740 90302
rect 12684 90290 12740 90300
rect 10780 89854 10782 89906
rect 10834 89854 10836 89906
rect 10780 89842 10836 89854
rect 7308 89796 7364 89806
rect 7980 89796 8036 89806
rect 8428 89796 8484 89806
rect 7308 89794 7588 89796
rect 7308 89742 7310 89794
rect 7362 89742 7588 89794
rect 7308 89740 7588 89742
rect 7308 89730 7364 89740
rect 4844 89570 5796 89572
rect 4844 89518 4846 89570
rect 4898 89518 5742 89570
rect 5794 89518 5796 89570
rect 4844 89516 5796 89518
rect 4476 88620 4740 88630
rect 4532 88564 4580 88620
rect 4636 88564 4684 88620
rect 4476 88554 4740 88564
rect 3276 88174 3278 88226
rect 3330 88174 3332 88226
rect 3276 87442 3332 88174
rect 3276 87390 3278 87442
rect 3330 87390 3332 87442
rect 3276 86658 3332 87390
rect 3276 86606 3278 86658
rect 3330 86606 3332 86658
rect 3276 85874 3332 86606
rect 3276 85822 3278 85874
rect 3330 85822 3332 85874
rect 3276 85090 3332 85822
rect 3276 85038 3278 85090
rect 3330 85038 3332 85090
rect 3276 84306 3332 85038
rect 3276 84254 3278 84306
rect 3330 84254 3332 84306
rect 3276 83748 3332 84254
rect 2156 83746 3332 83748
rect 2156 83694 2158 83746
rect 2210 83694 3332 83746
rect 2156 83692 3332 83694
rect 2156 83682 2212 83692
rect 3276 83522 3332 83692
rect 3276 83470 3278 83522
rect 3330 83470 3332 83522
rect 3276 83412 3332 83470
rect 4284 88226 4340 88238
rect 4284 88174 4286 88226
rect 4338 88174 4340 88226
rect 4284 87442 4340 88174
rect 4284 87390 4286 87442
rect 4338 87390 4340 87442
rect 4284 86658 4340 87390
rect 4732 88004 4788 88014
rect 4844 88004 4900 89516
rect 5740 89506 5796 89516
rect 6860 89012 6916 89022
rect 6860 88228 6916 88956
rect 7532 89012 7588 89740
rect 7980 89794 8484 89796
rect 7980 89742 7982 89794
rect 8034 89742 8430 89794
rect 8482 89742 8484 89794
rect 7980 89740 8484 89742
rect 7980 89012 8036 89740
rect 8428 89730 8484 89740
rect 9324 89794 9380 89806
rect 9324 89742 9326 89794
rect 9378 89742 9380 89794
rect 7532 89010 7924 89012
rect 7532 88958 7534 89010
rect 7586 88958 7924 89010
rect 7532 88956 7924 88958
rect 7532 88946 7588 88956
rect 7084 88228 7140 88238
rect 7868 88228 7924 88956
rect 6860 88226 7140 88228
rect 6860 88174 7086 88226
rect 7138 88174 7140 88226
rect 6860 88172 7140 88174
rect 4732 88002 4900 88004
rect 4732 87950 4734 88002
rect 4786 87950 4900 88002
rect 4732 87948 4900 87950
rect 4732 87332 4788 87948
rect 6860 87444 6916 87454
rect 7084 87444 7140 88172
rect 6860 87442 7140 87444
rect 6860 87390 6862 87442
rect 6914 87390 7140 87442
rect 6860 87388 7140 87390
rect 7756 88226 7924 88228
rect 7756 88174 7870 88226
rect 7922 88174 7924 88226
rect 7756 88172 7924 88174
rect 7756 88004 7812 88172
rect 7868 88162 7924 88172
rect 7980 88228 8036 88956
rect 7980 88162 8036 88172
rect 9100 88898 9156 88910
rect 9100 88846 9102 88898
rect 9154 88846 9156 88898
rect 7756 87442 7812 87948
rect 7756 87390 7758 87442
rect 7810 87390 7812 87442
rect 6860 87378 6916 87388
rect 7756 87378 7812 87390
rect 8428 88004 8484 88014
rect 5180 87332 5236 87342
rect 4732 87330 5236 87332
rect 4732 87278 4734 87330
rect 4786 87278 5182 87330
rect 5234 87278 5236 87330
rect 4732 87276 5236 87278
rect 4732 87266 4788 87276
rect 4476 87052 4740 87062
rect 4532 86996 4580 87052
rect 4636 86996 4684 87052
rect 4476 86986 4740 86996
rect 4284 86606 4286 86658
rect 4338 86606 4340 86658
rect 4284 86548 4340 86606
rect 4284 85876 4340 86492
rect 4732 86436 4788 86446
rect 4844 86436 4900 87276
rect 5180 87266 5236 87276
rect 4732 86434 4900 86436
rect 4732 86382 4734 86434
rect 4786 86382 4900 86434
rect 4732 86380 4900 86382
rect 4732 86370 4788 86380
rect 4620 85876 4676 85886
rect 4284 85874 4676 85876
rect 4284 85822 4286 85874
rect 4338 85822 4622 85874
rect 4674 85822 4676 85874
rect 4284 85820 4676 85822
rect 4284 85090 4340 85820
rect 4620 85810 4676 85820
rect 4844 85876 4900 86380
rect 6972 87220 7028 87230
rect 6972 86434 7028 87164
rect 8428 86658 8484 87948
rect 9100 87892 9156 88846
rect 9324 88116 9380 89742
rect 12908 89012 12964 92204
rect 13468 92258 13524 92316
rect 13580 92306 13636 92316
rect 13468 92206 13470 92258
rect 13522 92206 13524 92258
rect 13468 92194 13524 92206
rect 14028 91588 14084 91598
rect 13804 91586 14084 91588
rect 13804 91534 14030 91586
rect 14082 91534 14084 91586
rect 13804 91532 14084 91534
rect 13580 91364 13636 91374
rect 13580 91270 13636 91308
rect 13804 91362 13860 91532
rect 14028 91522 14084 91532
rect 13804 91310 13806 91362
rect 13858 91310 13860 91362
rect 13804 91298 13860 91310
rect 14252 91474 14308 92988
rect 14588 92818 14644 93548
rect 14588 92766 14590 92818
rect 14642 92766 14644 92818
rect 14588 92754 14644 92766
rect 14812 92484 14868 95452
rect 15148 95414 15204 95452
rect 16828 95396 16884 95406
rect 16828 95302 16884 95340
rect 17500 95396 17556 96014
rect 16492 95284 16548 95294
rect 16044 95282 16548 95284
rect 16044 95230 16494 95282
rect 16546 95230 16548 95282
rect 16044 95228 16548 95230
rect 15596 94724 15652 94734
rect 15596 94610 15652 94668
rect 15596 94558 15598 94610
rect 15650 94558 15652 94610
rect 15596 94546 15652 94558
rect 15932 94610 15988 94622
rect 15932 94558 15934 94610
rect 15986 94558 15988 94610
rect 15932 93716 15988 94558
rect 16044 94052 16100 95228
rect 16492 95218 16548 95228
rect 17500 95282 17556 95340
rect 17500 95230 17502 95282
rect 17554 95230 17556 95282
rect 16156 94500 16212 94510
rect 16716 94500 16772 94510
rect 16156 94498 16772 94500
rect 16156 94446 16158 94498
rect 16210 94446 16718 94498
rect 16770 94446 16772 94498
rect 16156 94444 16772 94446
rect 16156 94434 16212 94444
rect 16716 94434 16772 94444
rect 17500 94500 17556 95230
rect 16828 94386 16884 94398
rect 16828 94334 16830 94386
rect 16882 94334 16884 94386
rect 16828 94052 16884 94334
rect 17276 94274 17332 94286
rect 17276 94222 17278 94274
rect 17330 94222 17332 94274
rect 17276 94052 17332 94222
rect 16044 93996 16324 94052
rect 16268 93938 16324 93996
rect 16268 93886 16270 93938
rect 16322 93886 16324 93938
rect 16268 93874 16324 93886
rect 16828 93996 17276 94052
rect 15932 93650 15988 93660
rect 16604 93716 16660 93726
rect 16604 93622 16660 93660
rect 16828 93714 16884 93996
rect 17276 93986 17332 93996
rect 16828 93662 16830 93714
rect 16882 93662 16884 93714
rect 14364 92428 14868 92484
rect 14364 92372 14420 92428
rect 14364 92146 14420 92316
rect 14700 92260 14756 92270
rect 14700 92166 14756 92204
rect 14364 92094 14366 92146
rect 14418 92094 14420 92146
rect 14364 92082 14420 92094
rect 14588 91922 14644 91934
rect 14588 91870 14590 91922
rect 14642 91870 14644 91922
rect 14588 91586 14644 91870
rect 14588 91534 14590 91586
rect 14642 91534 14644 91586
rect 14588 91522 14644 91534
rect 14252 91422 14254 91474
rect 14306 91422 14308 91474
rect 13468 91250 13524 91262
rect 13468 91198 13470 91250
rect 13522 91198 13524 91250
rect 13468 91140 13524 91198
rect 14252 91140 14308 91422
rect 14700 91476 14756 91486
rect 14812 91476 14868 92428
rect 15148 92260 15204 92270
rect 15148 92166 15204 92204
rect 16828 92260 16884 93662
rect 17052 93716 17108 93726
rect 17052 92930 17108 93660
rect 17500 93714 17556 94444
rect 18396 96066 18452 96078
rect 18396 96014 18398 96066
rect 18450 96014 18452 96066
rect 18396 95282 18452 96014
rect 18396 95230 18398 95282
rect 18450 95230 18452 95282
rect 17500 93662 17502 93714
rect 17554 93662 17556 93714
rect 17500 93650 17556 93662
rect 17724 94274 17780 94286
rect 17724 94222 17726 94274
rect 17778 94222 17780 94274
rect 17724 94052 17780 94222
rect 17724 93380 17780 93996
rect 18396 93716 18452 95230
rect 19516 95844 19572 96238
rect 20076 95844 20132 95854
rect 20748 95844 20804 95854
rect 19516 95842 20804 95844
rect 19516 95790 20078 95842
rect 20130 95790 20750 95842
rect 20802 95790 20804 95842
rect 19516 95788 20804 95790
rect 19516 95732 19572 95788
rect 20076 95778 20132 95788
rect 19516 95172 19572 95676
rect 19836 95676 20100 95686
rect 19892 95620 19940 95676
rect 19996 95620 20044 95676
rect 19836 95610 20100 95620
rect 20636 95284 20692 95788
rect 20748 95778 20804 95788
rect 19852 95172 19908 95182
rect 19516 95170 19908 95172
rect 19516 95118 19854 95170
rect 19906 95118 19908 95170
rect 19516 95116 19908 95118
rect 19516 95058 19572 95116
rect 19852 95106 19908 95116
rect 19516 95006 19518 95058
rect 19570 95006 19572 95058
rect 18508 94500 18564 94510
rect 18508 94406 18564 94444
rect 19292 94498 19348 94510
rect 19292 94446 19294 94498
rect 19346 94446 19348 94498
rect 18396 93622 18452 93660
rect 19292 93716 19348 94446
rect 17724 93314 17780 93324
rect 19292 93154 19348 93660
rect 19516 93490 19572 95006
rect 20636 94722 20692 95228
rect 20636 94670 20638 94722
rect 20690 94670 20692 94722
rect 20636 94658 20692 94670
rect 20300 94388 20356 94398
rect 19836 94108 20100 94118
rect 19892 94052 19940 94108
rect 19996 94052 20044 94108
rect 19836 94042 20100 94052
rect 20300 93716 20356 94332
rect 20636 93940 20692 93950
rect 20636 93846 20692 93884
rect 20300 93714 20692 93716
rect 20300 93662 20302 93714
rect 20354 93662 20692 93714
rect 20300 93660 20692 93662
rect 20300 93650 20356 93660
rect 19516 93438 19518 93490
rect 19570 93438 19572 93490
rect 19516 93426 19572 93438
rect 20076 93602 20132 93614
rect 20076 93550 20078 93602
rect 20130 93550 20132 93602
rect 20076 93380 20132 93550
rect 20076 93314 20132 93324
rect 19292 93102 19294 93154
rect 19346 93102 19348 93154
rect 19292 93090 19348 93102
rect 17276 93044 17332 93054
rect 17276 92950 17332 92988
rect 18620 93044 18676 93054
rect 18620 92950 18676 92988
rect 17052 92878 17054 92930
rect 17106 92878 17108 92930
rect 17052 92866 17108 92878
rect 17948 92930 18004 92942
rect 17948 92878 17950 92930
rect 18002 92878 18004 92930
rect 17948 92708 18004 92878
rect 17948 92642 18004 92652
rect 19404 92818 19460 92830
rect 19404 92766 19406 92818
rect 19458 92766 19460 92818
rect 19404 92708 19460 92766
rect 19404 92642 19460 92652
rect 19836 92540 20100 92550
rect 19892 92484 19940 92540
rect 19996 92484 20044 92540
rect 19836 92474 20100 92484
rect 20636 92260 20692 93660
rect 20748 93380 20804 93390
rect 20748 93042 20804 93324
rect 20748 92990 20750 93042
rect 20802 92990 20804 93042
rect 20748 92978 20804 92990
rect 20748 92260 20804 92270
rect 20636 92258 20804 92260
rect 20636 92206 20750 92258
rect 20802 92206 20804 92258
rect 20636 92204 20804 92206
rect 16828 92194 16884 92204
rect 20748 92194 20804 92204
rect 14700 91474 14868 91476
rect 14700 91422 14702 91474
rect 14754 91422 14868 91474
rect 14700 91420 14868 91422
rect 14700 91410 14756 91420
rect 13468 91084 14308 91140
rect 14252 90748 14308 91084
rect 19836 90972 20100 90982
rect 19892 90916 19940 90972
rect 19996 90916 20044 90972
rect 19836 90906 20100 90916
rect 14140 90692 14308 90748
rect 12796 89010 12964 89012
rect 12796 88958 12910 89010
rect 12962 88958 12964 89010
rect 12796 88956 12964 88958
rect 12796 88338 12852 88956
rect 12908 88946 12964 88956
rect 13356 89012 13412 89022
rect 13356 88918 13412 88956
rect 12796 88286 12798 88338
rect 12850 88286 12852 88338
rect 9324 88050 9380 88060
rect 9660 88228 9716 88238
rect 9436 88002 9492 88014
rect 9436 87950 9438 88002
rect 9490 87950 9492 88002
rect 9436 87892 9492 87950
rect 9548 87892 9604 87902
rect 9100 87836 9548 87892
rect 9100 87666 9156 87836
rect 9548 87826 9604 87836
rect 9100 87614 9102 87666
rect 9154 87614 9156 87666
rect 9100 87220 9156 87614
rect 9660 87444 9716 88172
rect 9100 87154 9156 87164
rect 9324 87442 9716 87444
rect 9324 87390 9662 87442
rect 9714 87390 9716 87442
rect 9324 87388 9716 87390
rect 8428 86606 8430 86658
rect 8482 86606 8484 86658
rect 8428 86594 8484 86606
rect 9324 86660 9380 87388
rect 9660 87378 9716 87388
rect 10556 88226 10612 88238
rect 10556 88174 10558 88226
rect 10610 88174 10612 88226
rect 10556 88116 10612 88174
rect 10556 87556 10612 88060
rect 12572 88226 12628 88238
rect 12572 88174 12574 88226
rect 12626 88174 12628 88226
rect 10556 87442 10612 87500
rect 10556 87390 10558 87442
rect 10610 87390 10612 87442
rect 10556 87378 10612 87390
rect 10668 88004 10724 88014
rect 9324 86566 9380 86604
rect 10108 86660 10164 86670
rect 10108 86566 10164 86604
rect 10668 86658 10724 87948
rect 12012 88002 12068 88014
rect 12012 87950 12014 88002
rect 12066 87950 12068 88002
rect 12012 87892 12068 87950
rect 12236 88004 12292 88014
rect 12236 87910 12292 87948
rect 11900 87668 11956 87678
rect 12012 87668 12068 87836
rect 11900 87666 12068 87668
rect 11900 87614 11902 87666
rect 11954 87614 12068 87666
rect 11900 87612 12068 87614
rect 12460 87780 12516 87790
rect 11900 87602 11956 87612
rect 12348 87444 12404 87454
rect 12460 87444 12516 87724
rect 12348 87442 12516 87444
rect 12348 87390 12350 87442
rect 12402 87390 12516 87442
rect 12348 87388 12516 87390
rect 12348 87378 12404 87388
rect 12572 87218 12628 88174
rect 12572 87166 12574 87218
rect 12626 87166 12628 87218
rect 10668 86606 10670 86658
rect 10722 86606 10724 86658
rect 10668 86594 10724 86606
rect 11676 86658 11732 86670
rect 11676 86606 11678 86658
rect 11730 86606 11732 86658
rect 10892 86548 10948 86558
rect 10892 86454 10948 86492
rect 6972 86382 6974 86434
rect 7026 86382 7028 86434
rect 6972 86100 7028 86382
rect 7308 86100 7364 86110
rect 6972 86098 7364 86100
rect 6972 86046 7310 86098
rect 7362 86046 7364 86098
rect 6972 86044 7364 86046
rect 5404 85876 5460 85886
rect 4844 85820 5404 85876
rect 4476 85484 4740 85494
rect 4532 85428 4580 85484
rect 4636 85428 4684 85484
rect 4476 85418 4740 85428
rect 4284 85038 4286 85090
rect 4338 85038 4340 85090
rect 4284 84306 4340 85038
rect 4284 84254 4286 84306
rect 4338 84254 4340 84306
rect 4284 83522 4340 84254
rect 4732 84868 4788 84878
rect 4844 84868 4900 85820
rect 5404 85782 5460 85820
rect 6972 85876 7028 86044
rect 7308 86034 7364 86044
rect 11564 86100 11620 86110
rect 11564 85986 11620 86044
rect 11676 86098 11732 86606
rect 12572 86546 12628 87166
rect 12572 86494 12574 86546
rect 12626 86494 12628 86546
rect 12572 86482 12628 86494
rect 11676 86046 11678 86098
rect 11730 86046 11732 86098
rect 11676 86034 11732 86046
rect 12124 86100 12180 86110
rect 12124 86006 12180 86044
rect 12796 86100 12852 88286
rect 14028 88898 14084 88910
rect 14028 88846 14030 88898
rect 14082 88846 14084 88898
rect 14028 88226 14084 88846
rect 14028 88174 14030 88226
rect 14082 88174 14084 88226
rect 14028 88162 14084 88174
rect 13804 88004 13860 88014
rect 13580 87556 13636 87566
rect 13580 87462 13636 87500
rect 13020 87444 13076 87454
rect 13020 87350 13076 87388
rect 12796 86034 12852 86044
rect 13804 85988 13860 87948
rect 14140 87780 14196 90692
rect 19964 89796 20020 89806
rect 19628 89740 19964 89796
rect 15932 89570 15988 89582
rect 15932 89518 15934 89570
rect 15986 89518 15988 89570
rect 14252 89124 14308 89134
rect 14252 88004 14308 89068
rect 15932 89124 15988 89518
rect 16492 89572 16548 89582
rect 17276 89572 17332 89582
rect 17500 89572 17556 89582
rect 16492 89570 17500 89572
rect 16492 89518 16494 89570
rect 16546 89518 17278 89570
rect 17330 89518 17500 89570
rect 16492 89516 17500 89518
rect 16492 89124 16548 89516
rect 17276 89506 17332 89516
rect 15932 89058 15988 89068
rect 16044 89068 16548 89124
rect 16716 89124 16772 89134
rect 16044 89012 16100 89068
rect 16716 89030 16772 89068
rect 15484 88338 15540 88350
rect 15484 88286 15486 88338
rect 15538 88286 15540 88338
rect 15260 88226 15316 88238
rect 15260 88174 15262 88226
rect 15314 88174 15316 88226
rect 14364 88114 14420 88126
rect 14700 88116 14756 88126
rect 14364 88062 14366 88114
rect 14418 88062 14420 88114
rect 14364 88004 14420 88062
rect 14588 88114 14756 88116
rect 14588 88062 14702 88114
rect 14754 88062 14756 88114
rect 14588 88060 14756 88062
rect 14588 88004 14644 88060
rect 14700 88050 14756 88060
rect 14364 87948 14644 88004
rect 14252 87910 14308 87948
rect 14196 87724 14420 87780
rect 14140 87686 14196 87724
rect 14364 87666 14420 87724
rect 14364 87614 14366 87666
rect 14418 87614 14420 87666
rect 14364 87602 14420 87614
rect 15260 87668 15316 88174
rect 15260 87574 15316 87612
rect 13916 87444 13972 87454
rect 13916 87350 13972 87388
rect 15484 87444 15540 88286
rect 16044 88228 16100 88956
rect 16828 89010 16884 89022
rect 16828 88958 16830 89010
rect 16882 88958 16884 89010
rect 16156 88900 16212 88910
rect 16156 88898 16324 88900
rect 16156 88846 16158 88898
rect 16210 88846 16324 88898
rect 16156 88844 16324 88846
rect 16156 88834 16212 88844
rect 16156 88228 16212 88238
rect 15932 88226 16212 88228
rect 15932 88174 16158 88226
rect 16210 88174 16212 88226
rect 15932 88172 16212 88174
rect 15708 87668 15764 87678
rect 15708 87574 15764 87612
rect 15596 87444 15652 87454
rect 15484 87388 15596 87444
rect 11564 85934 11566 85986
rect 11618 85934 11620 85986
rect 11564 85922 11620 85934
rect 13580 85932 13860 85988
rect 14140 86548 14196 86558
rect 6972 85782 7028 85820
rect 4732 84866 4900 84868
rect 4732 84814 4734 84866
rect 4786 84814 4900 84866
rect 4732 84812 4900 84814
rect 12908 84868 12964 84878
rect 4732 84196 4788 84812
rect 12908 84774 12964 84812
rect 4956 84532 5012 84542
rect 4732 84194 4900 84196
rect 4732 84142 4734 84194
rect 4786 84142 4900 84194
rect 4732 84140 4900 84142
rect 4732 84130 4788 84140
rect 4476 83916 4740 83926
rect 4532 83860 4580 83916
rect 4636 83860 4684 83916
rect 4476 83850 4740 83860
rect 4284 83470 4286 83522
rect 4338 83470 4340 83522
rect 4284 83458 4340 83470
rect 3276 83346 3332 83356
rect 4396 83412 4452 83422
rect 4732 83412 4788 83422
rect 4844 83412 4900 84140
rect 4452 83410 4900 83412
rect 4452 83358 4734 83410
rect 4786 83358 4900 83410
rect 4452 83356 4900 83358
rect 4396 83346 4452 83356
rect 4732 83346 4788 83356
rect 4956 82628 5012 84476
rect 8764 84194 8820 84206
rect 8764 84142 8766 84194
rect 8818 84142 8820 84194
rect 8092 83524 8148 83534
rect 7980 83522 8148 83524
rect 7980 83470 8094 83522
rect 8146 83470 8148 83522
rect 7980 83468 8148 83470
rect 4956 82562 5012 82572
rect 6076 82628 6132 82638
rect 6076 82534 6132 82572
rect 7196 82516 7252 82526
rect 4476 82348 4740 82358
rect 4532 82292 4580 82348
rect 4636 82292 4684 82348
rect 4476 82282 4740 82292
rect 5180 82012 6356 82068
rect 5180 81954 5236 82012
rect 5180 81902 5182 81954
rect 5234 81902 5236 81954
rect 5180 81890 5236 81902
rect 6300 81954 6356 82012
rect 6300 81902 6302 81954
rect 6354 81902 6356 81954
rect 6300 81890 6356 81902
rect 6636 81956 6692 81966
rect 6636 81862 6692 81900
rect 4844 81842 4900 81854
rect 4844 81790 4846 81842
rect 4898 81790 4900 81842
rect 4620 81732 4676 81742
rect 4844 81732 4900 81790
rect 6076 81842 6132 81854
rect 6076 81790 6078 81842
rect 6130 81790 6132 81842
rect 4620 81730 4900 81732
rect 4620 81678 4622 81730
rect 4674 81678 4900 81730
rect 4620 81676 4900 81678
rect 4620 81666 4676 81676
rect 4844 81284 4900 81676
rect 4844 81218 4900 81228
rect 4956 81730 5012 81742
rect 4956 81678 4958 81730
rect 5010 81678 5012 81730
rect 3724 81060 3780 81070
rect 4956 81060 5012 81678
rect 5852 81732 5908 81742
rect 6076 81732 6132 81790
rect 6412 81732 6468 81742
rect 5908 81676 6132 81732
rect 6188 81730 6468 81732
rect 6188 81678 6414 81730
rect 6466 81678 6468 81730
rect 6188 81676 6468 81678
rect 5852 81638 5908 81676
rect 6188 81396 6244 81676
rect 6412 81666 6468 81676
rect 7196 81732 7252 82460
rect 7980 82516 8036 83468
rect 8092 83458 8148 83468
rect 8428 83410 8484 83422
rect 8428 83358 8430 83410
rect 8482 83358 8484 83410
rect 8316 83298 8372 83310
rect 8316 83246 8318 83298
rect 8370 83246 8372 83298
rect 8204 82852 8260 82862
rect 8316 82852 8372 83246
rect 8428 82964 8484 83358
rect 8428 82898 8484 82908
rect 8204 82850 8372 82852
rect 8204 82798 8206 82850
rect 8258 82798 8372 82850
rect 8204 82796 8372 82798
rect 8204 82786 8260 82796
rect 7980 82450 8036 82460
rect 8764 82516 8820 84142
rect 12572 84196 12628 84206
rect 9100 83746 9156 83758
rect 9100 83694 9102 83746
rect 9154 83694 9156 83746
rect 8764 82450 8820 82460
rect 8988 82740 9044 82750
rect 9100 82740 9156 83694
rect 9772 83746 9828 83758
rect 9772 83694 9774 83746
rect 9826 83694 9828 83746
rect 9772 83634 9828 83694
rect 9772 83582 9774 83634
rect 9826 83582 9828 83634
rect 9772 83570 9828 83582
rect 9324 83298 9380 83310
rect 9324 83246 9326 83298
rect 9378 83246 9380 83298
rect 9324 83188 9380 83246
rect 9324 83132 9604 83188
rect 8988 82738 9156 82740
rect 8988 82686 8990 82738
rect 9042 82686 9156 82738
rect 8988 82684 9156 82686
rect 9548 82738 9604 83132
rect 9548 82686 9550 82738
rect 9602 82686 9604 82738
rect 5852 81340 6244 81396
rect 6524 81396 6580 81406
rect 7084 81396 7140 81406
rect 3724 81058 5012 81060
rect 3724 81006 3726 81058
rect 3778 81006 5012 81058
rect 3724 81004 5012 81006
rect 3724 80994 3780 81004
rect 4476 80780 4740 80790
rect 4532 80724 4580 80780
rect 4636 80724 4684 80780
rect 4476 80714 4740 80724
rect 4476 79212 4740 79222
rect 4532 79156 4580 79212
rect 4636 79156 4684 79212
rect 4476 79146 4740 79156
rect 3612 78484 3668 78494
rect 3612 77922 3668 78428
rect 3612 77870 3614 77922
rect 3666 77870 3668 77922
rect 2156 74228 2212 74238
rect 2156 74134 2212 74172
rect 2156 69410 2212 69422
rect 2156 69358 2158 69410
rect 2210 69358 2212 69410
rect 1820 67060 1876 67070
rect 2156 67060 2212 69358
rect 2940 69300 2996 69310
rect 2940 69298 3332 69300
rect 2940 69246 2942 69298
rect 2994 69246 3332 69298
rect 2940 69244 3332 69246
rect 2940 69234 2996 69244
rect 3276 68852 3332 69244
rect 3500 68852 3556 68862
rect 3276 68850 3556 68852
rect 3276 68798 3502 68850
rect 3554 68798 3556 68850
rect 3276 68796 3556 68798
rect 3500 68786 3556 68796
rect 3612 67844 3668 77870
rect 4476 77644 4740 77654
rect 4532 77588 4580 77644
rect 4636 77588 4684 77644
rect 4476 77578 4740 77588
rect 4476 76076 4740 76086
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4476 76010 4740 76020
rect 4844 75796 4900 75806
rect 4284 75684 4340 75694
rect 4172 74788 4228 74798
rect 4172 74116 4228 74732
rect 4284 74226 4340 75628
rect 4396 74788 4452 74798
rect 4396 74694 4452 74732
rect 4844 74676 4900 75740
rect 4844 74610 4900 74620
rect 4476 74508 4740 74518
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4476 74442 4740 74452
rect 4284 74174 4286 74226
rect 4338 74174 4340 74226
rect 4284 74162 4340 74174
rect 3500 67788 3668 67844
rect 3724 74004 3780 74014
rect 3164 67730 3220 67742
rect 3164 67678 3166 67730
rect 3218 67678 3220 67730
rect 2828 67618 2884 67630
rect 2828 67566 2830 67618
rect 2882 67566 2884 67618
rect 2828 67228 2884 67566
rect 2492 67172 2884 67228
rect 3164 67228 3220 67678
rect 3164 67172 3444 67228
rect 2492 67170 2548 67172
rect 2492 67118 2494 67170
rect 2546 67118 2548 67170
rect 2492 67106 2548 67118
rect 1820 67058 2212 67060
rect 1820 67006 1822 67058
rect 1874 67006 2212 67058
rect 1820 67004 2212 67006
rect 1820 66994 1876 67004
rect 2156 65492 2212 67004
rect 3388 66498 3444 67172
rect 3388 66446 3390 66498
rect 3442 66446 3444 66498
rect 3388 66434 3444 66446
rect 2940 65492 2996 65502
rect 2156 65490 2996 65492
rect 2156 65438 2942 65490
rect 2994 65438 2996 65490
rect 2156 65436 2996 65438
rect 1708 62354 1764 62366
rect 1708 62302 1710 62354
rect 1762 62302 1764 62354
rect 1708 62244 1764 62302
rect 1708 62178 1764 62188
rect 2492 62244 2548 62254
rect 2940 62244 2996 65436
rect 2492 62242 2884 62244
rect 2492 62190 2494 62242
rect 2546 62190 2884 62242
rect 2492 62188 2884 62190
rect 2492 62178 2548 62188
rect 2828 61458 2884 62188
rect 2940 62178 2996 62188
rect 2828 61406 2830 61458
rect 2882 61406 2884 61458
rect 2828 61394 2884 61406
rect 3164 61460 3220 61470
rect 3164 61458 3444 61460
rect 3164 61406 3166 61458
rect 3218 61406 3444 61458
rect 3164 61404 3444 61406
rect 3164 61394 3220 61404
rect 3388 61010 3444 61404
rect 3388 60958 3390 61010
rect 3442 60958 3444 61010
rect 3388 60946 3444 60958
rect 3388 60564 3444 60574
rect 1820 60002 1876 60014
rect 1820 59950 1822 60002
rect 1874 59950 1876 60002
rect 1820 59220 1876 59950
rect 2492 59892 2548 59902
rect 2492 59890 2884 59892
rect 2492 59838 2494 59890
rect 2546 59838 2884 59890
rect 2492 59836 2884 59838
rect 2492 59826 2548 59836
rect 1820 57650 1876 59164
rect 1820 57598 1822 57650
rect 1874 57598 1876 57650
rect 1820 57586 1876 57598
rect 2492 57540 2548 57550
rect 2492 57538 2772 57540
rect 2492 57486 2494 57538
rect 2546 57486 2772 57538
rect 2492 57484 2772 57486
rect 2492 57474 2548 57484
rect 2716 56308 2772 57484
rect 2828 56754 2884 59836
rect 2828 56702 2830 56754
rect 2882 56702 2884 56754
rect 2828 56690 2884 56702
rect 3052 56866 3108 56878
rect 3052 56814 3054 56866
rect 3106 56814 3108 56866
rect 2828 56308 2884 56318
rect 2716 56306 2884 56308
rect 2716 56254 2830 56306
rect 2882 56254 2884 56306
rect 2716 56252 2884 56254
rect 2828 56242 2884 56252
rect 3052 55412 3108 56814
rect 3052 55346 3108 55356
rect 3164 56082 3220 56094
rect 3164 56030 3166 56082
rect 3218 56030 3220 56082
rect 3164 54740 3220 56030
rect 3388 55972 3444 60508
rect 3388 55906 3444 55916
rect 3500 55748 3556 67788
rect 3724 66500 3780 73948
rect 4172 70588 4228 74060
rect 4476 72940 4740 72950
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4476 72874 4740 72884
rect 4476 71372 4740 71382
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4476 71306 4740 71316
rect 4060 70532 4228 70588
rect 3836 68626 3892 68638
rect 3836 68574 3838 68626
rect 3890 68574 3892 68626
rect 3836 68516 3892 68574
rect 3836 68450 3892 68460
rect 3724 66444 3892 66500
rect 3612 66388 3668 66398
rect 3668 66332 3780 66388
rect 3612 66322 3668 66332
rect 3724 66274 3780 66332
rect 3724 66222 3726 66274
rect 3778 66222 3780 66274
rect 3724 66210 3780 66222
rect 3724 66052 3780 66062
rect 3612 65996 3724 66052
rect 3612 65602 3668 65996
rect 3724 65986 3780 65996
rect 3612 65550 3614 65602
rect 3666 65550 3668 65602
rect 3612 65538 3668 65550
rect 3836 65492 3892 66444
rect 3724 65436 3892 65492
rect 3948 66274 4004 66286
rect 3948 66222 3950 66274
rect 4002 66222 4004 66274
rect 3724 65380 3780 65436
rect 3164 54674 3220 54684
rect 3388 55692 3556 55748
rect 3612 65324 3780 65380
rect 3388 53732 3444 55692
rect 3612 55636 3668 65324
rect 3836 65268 3892 65278
rect 3836 64930 3892 65212
rect 3836 64878 3838 64930
rect 3890 64878 3892 64930
rect 3836 64866 3892 64878
rect 3948 61684 4004 66222
rect 3948 61618 4004 61628
rect 4060 61460 4116 70532
rect 4476 69804 4740 69814
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4476 69738 4740 69748
rect 4508 68628 4564 68638
rect 4508 68534 4564 68572
rect 4476 68236 4740 68246
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4476 68170 4740 68180
rect 4620 66948 4676 66958
rect 4620 66946 4900 66948
rect 4620 66894 4622 66946
rect 4674 66894 4900 66946
rect 4620 66892 4900 66894
rect 4620 66882 4676 66892
rect 4476 66668 4740 66678
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4476 66602 4740 66612
rect 4396 66388 4452 66398
rect 4284 66052 4340 66062
rect 4284 65958 4340 65996
rect 4396 65268 4452 66332
rect 4172 65212 4452 65268
rect 4508 66274 4564 66286
rect 4508 66222 4510 66274
rect 4562 66222 4564 66274
rect 4508 65268 4564 66222
rect 4172 64818 4228 65212
rect 4508 65202 4564 65212
rect 4476 65100 4740 65110
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4476 65034 4740 65044
rect 4172 64766 4174 64818
rect 4226 64766 4228 64818
rect 4172 64596 4228 64766
rect 4396 64820 4452 64830
rect 4844 64820 4900 66892
rect 4396 64818 4900 64820
rect 4396 64766 4398 64818
rect 4450 64766 4900 64818
rect 4396 64764 4900 64766
rect 4396 64754 4452 64764
rect 4172 64530 4228 64540
rect 4620 63812 4676 64764
rect 4844 64596 4900 64606
rect 4844 64502 4900 64540
rect 4620 63746 4676 63756
rect 4476 63532 4740 63542
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4476 63466 4740 63476
rect 4620 62242 4676 62254
rect 4620 62190 4622 62242
rect 4674 62190 4676 62242
rect 4620 62188 4676 62190
rect 3724 61404 4116 61460
rect 4284 62132 4676 62188
rect 3724 60788 3780 61404
rect 4172 61348 4228 61358
rect 4172 61254 4228 61292
rect 4284 60900 4340 62132
rect 4476 61964 4740 61974
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4476 61898 4740 61908
rect 3724 60732 3892 60788
rect 3724 60564 3780 60574
rect 3724 60470 3780 60508
rect 3836 60340 3892 60732
rect 4284 60786 4340 60844
rect 4284 60734 4286 60786
rect 4338 60734 4340 60786
rect 4284 60722 4340 60734
rect 4396 61684 4452 61694
rect 3500 55580 3668 55636
rect 3724 60284 3892 60340
rect 3948 60674 4004 60686
rect 3948 60622 3950 60674
rect 4002 60622 4004 60674
rect 3500 54964 3556 55580
rect 3612 55412 3668 55422
rect 3612 55318 3668 55356
rect 3500 54898 3556 54908
rect 3612 54740 3668 54750
rect 3612 54646 3668 54684
rect 3724 53844 3780 60284
rect 3836 59218 3892 59230
rect 3836 59166 3838 59218
rect 3890 59166 3892 59218
rect 3836 59108 3892 59166
rect 3836 59042 3892 59052
rect 3948 58212 4004 60622
rect 4396 60564 4452 61628
rect 4284 60508 4452 60564
rect 4508 61348 4564 61358
rect 4508 60564 4564 61292
rect 4284 60228 4340 60508
rect 4508 60498 4564 60508
rect 4844 60562 4900 60574
rect 4844 60510 4846 60562
rect 4898 60510 4900 60562
rect 4476 60396 4740 60406
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4476 60330 4740 60340
rect 4284 60172 4676 60228
rect 4284 58436 4340 60172
rect 4620 60114 4676 60172
rect 4620 60062 4622 60114
rect 4674 60062 4676 60114
rect 4620 60050 4676 60062
rect 4844 60004 4900 60510
rect 4844 59938 4900 59948
rect 4620 59780 4676 59790
rect 4620 59330 4676 59724
rect 4620 59278 4622 59330
rect 4674 59278 4676 59330
rect 4620 59266 4676 59278
rect 4476 58828 4740 58838
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4476 58762 4740 58772
rect 4396 58436 4452 58446
rect 4844 58436 4900 58446
rect 4284 58434 4452 58436
rect 4284 58382 4398 58434
rect 4450 58382 4452 58434
rect 4284 58380 4452 58382
rect 4396 58370 4452 58380
rect 4508 58434 4900 58436
rect 4508 58382 4846 58434
rect 4898 58382 4900 58434
rect 4508 58380 4900 58382
rect 4508 58212 4564 58380
rect 4844 58370 4900 58380
rect 3948 58156 4564 58212
rect 4508 57540 4564 58156
rect 4620 58212 4676 58222
rect 4620 58118 4676 58156
rect 4732 58212 4788 58222
rect 4732 58210 4900 58212
rect 4732 58158 4734 58210
rect 4786 58158 4900 58210
rect 4732 58156 4900 58158
rect 4732 58146 4788 58156
rect 4620 57540 4676 57550
rect 4508 57538 4676 57540
rect 4508 57486 4622 57538
rect 4674 57486 4676 57538
rect 4508 57484 4676 57486
rect 4620 57474 4676 57484
rect 4476 57260 4740 57270
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4476 57194 4740 57204
rect 4476 55692 4740 55702
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4476 55626 4740 55636
rect 4844 55524 4900 58156
rect 3612 53788 3780 53844
rect 3836 55468 4900 55524
rect 3388 53676 3556 53732
rect 3388 53508 3444 53518
rect 2492 53506 3444 53508
rect 2492 53454 3390 53506
rect 3442 53454 3444 53506
rect 2492 53452 3444 53454
rect 2492 53058 2548 53452
rect 3388 53442 3444 53452
rect 2492 53006 2494 53058
rect 2546 53006 2548 53058
rect 2492 52994 2548 53006
rect 1820 52946 1876 52958
rect 3500 52948 3556 53676
rect 1820 52894 1822 52946
rect 1874 52894 1876 52946
rect 1820 52164 1876 52894
rect 3388 52892 3556 52948
rect 2044 52164 2100 52174
rect 1820 52108 2044 52164
rect 2044 52070 2100 52108
rect 2716 52052 2772 52062
rect 2716 51958 2772 51996
rect 3388 51828 3444 52892
rect 3276 51772 3444 51828
rect 3500 52724 3556 52734
rect 3164 51492 3220 51502
rect 2492 51490 3220 51492
rect 2492 51438 3166 51490
rect 3218 51438 3220 51490
rect 2492 51436 3220 51438
rect 2492 49922 2548 51436
rect 3164 51426 3220 51436
rect 3276 51156 3332 51772
rect 3500 51490 3556 52668
rect 3500 51438 3502 51490
rect 3554 51438 3556 51490
rect 3500 51426 3556 51438
rect 3276 51100 3444 51156
rect 2492 49870 2494 49922
rect 2546 49870 2548 49922
rect 2492 49858 2548 49870
rect 1820 49810 1876 49822
rect 1820 49758 1822 49810
rect 1874 49758 1876 49810
rect 1820 47068 1876 49758
rect 2940 48356 2996 48366
rect 2940 47570 2996 48300
rect 2940 47518 2942 47570
rect 2994 47518 2996 47570
rect 2940 47506 2996 47518
rect 2268 47458 2324 47470
rect 2268 47406 2270 47458
rect 2322 47406 2324 47458
rect 2268 47124 2324 47406
rect 1820 47012 2324 47068
rect 1820 45106 1876 47012
rect 1820 45054 1822 45106
rect 1874 45054 1876 45106
rect 1820 43540 1876 45054
rect 3276 45668 3332 45678
rect 2492 44996 2548 45006
rect 2492 44994 2996 44996
rect 2492 44942 2494 44994
rect 2546 44942 2996 44994
rect 2492 44940 2996 44942
rect 2492 44930 2548 44940
rect 2268 44324 2324 44334
rect 2268 44230 2324 44268
rect 2940 44210 2996 44940
rect 3276 44322 3332 45612
rect 3276 44270 3278 44322
rect 3330 44270 3332 44322
rect 3276 44258 3332 44270
rect 2940 44158 2942 44210
rect 2994 44158 2996 44210
rect 2940 44146 2996 44158
rect 2604 44098 2660 44110
rect 2604 44046 2606 44098
rect 2658 44046 2660 44098
rect 2604 43708 2660 44046
rect 2604 43652 2996 43708
rect 2940 43650 2996 43652
rect 2940 43598 2942 43650
rect 2994 43598 2996 43650
rect 2940 43586 2996 43598
rect 2156 43540 2212 43550
rect 1820 43538 2212 43540
rect 1820 43486 2158 43538
rect 2210 43486 2212 43538
rect 1820 43484 2212 43486
rect 1820 38834 1876 43484
rect 2156 43474 2212 43484
rect 3164 40404 3220 40414
rect 3164 39618 3220 40348
rect 3164 39566 3166 39618
rect 3218 39566 3220 39618
rect 3164 39554 3220 39566
rect 2940 39396 2996 39406
rect 2492 39394 2996 39396
rect 2492 39342 2942 39394
rect 2994 39342 2996 39394
rect 2492 39340 2996 39342
rect 2492 38946 2548 39340
rect 2940 39330 2996 39340
rect 2492 38894 2494 38946
rect 2546 38894 2548 38946
rect 2492 38882 2548 38894
rect 1820 38782 1822 38834
rect 1874 38782 1876 38834
rect 1820 38724 1876 38782
rect 1932 38724 1988 38734
rect 1820 38668 1932 38724
rect 1932 38658 1988 38668
rect 3276 37938 3332 37950
rect 3276 37886 3278 37938
rect 3330 37886 3332 37938
rect 2940 37828 2996 37838
rect 2492 37826 2996 37828
rect 2492 37774 2942 37826
rect 2994 37774 2996 37826
rect 2492 37772 2996 37774
rect 2492 37378 2548 37772
rect 2940 37762 2996 37772
rect 3276 37828 3332 37886
rect 3276 37762 3332 37772
rect 2492 37326 2494 37378
rect 2546 37326 2548 37378
rect 2492 37314 2548 37326
rect 1820 37266 1876 37278
rect 1820 37214 1822 37266
rect 1874 37214 1876 37266
rect 1820 34130 1876 37214
rect 3388 35588 3444 51100
rect 3612 50428 3668 53788
rect 3724 53620 3780 53630
rect 3724 53526 3780 53564
rect 3836 52276 3892 55468
rect 3948 55298 4004 55310
rect 4172 55300 4228 55310
rect 3948 55246 3950 55298
rect 4002 55246 4004 55298
rect 3948 54404 4004 55246
rect 3948 54310 4004 54348
rect 4060 55298 4228 55300
rect 4060 55246 4174 55298
rect 4226 55246 4228 55298
rect 4060 55244 4228 55246
rect 3500 50372 3668 50428
rect 3724 52220 3892 52276
rect 3948 54068 4004 54078
rect 3724 50428 3780 52220
rect 3836 52052 3892 52062
rect 3836 51602 3892 51996
rect 3836 51550 3838 51602
rect 3890 51550 3892 51602
rect 3836 51538 3892 51550
rect 3724 50372 3892 50428
rect 3500 45108 3556 50372
rect 3724 48356 3780 48366
rect 3724 48262 3780 48300
rect 3612 45668 3668 45678
rect 3612 45574 3668 45612
rect 3500 45042 3556 45052
rect 3612 44324 3668 44334
rect 3612 44230 3668 44268
rect 3612 40516 3668 40526
rect 3612 35700 3668 40460
rect 3612 35634 3668 35644
rect 3724 39396 3780 39406
rect 3164 35532 3444 35588
rect 3164 35252 3220 35532
rect 3612 35476 3668 35486
rect 3164 35186 3220 35196
rect 3276 35474 3668 35476
rect 3276 35422 3614 35474
rect 3666 35422 3668 35474
rect 3276 35420 3668 35422
rect 3276 34914 3332 35420
rect 3612 35410 3668 35420
rect 3276 34862 3278 34914
rect 3330 34862 3332 34914
rect 3276 34850 3332 34862
rect 3612 35252 3668 35262
rect 2940 34692 2996 34702
rect 2492 34690 2996 34692
rect 2492 34638 2942 34690
rect 2994 34638 2996 34690
rect 2492 34636 2996 34638
rect 2492 34242 2548 34636
rect 2940 34626 2996 34636
rect 2492 34190 2494 34242
rect 2546 34190 2548 34242
rect 2492 34178 2548 34190
rect 1820 34078 1822 34130
rect 1874 34078 1876 34130
rect 1820 31948 1876 34078
rect 2492 32452 2548 32462
rect 2492 31948 2548 32396
rect 1708 31892 2548 31948
rect 1708 29426 1764 31892
rect 2492 30994 2548 31892
rect 2492 30942 2494 30994
rect 2546 30942 2548 30994
rect 2492 30930 2548 30942
rect 3164 30884 3220 30894
rect 3164 30882 3556 30884
rect 3164 30830 3166 30882
rect 3218 30830 3556 30882
rect 3164 30828 3556 30830
rect 3164 30818 3220 30828
rect 3500 30098 3556 30828
rect 3500 30046 3502 30098
rect 3554 30046 3556 30098
rect 3500 30034 3556 30046
rect 1708 29374 1710 29426
rect 1762 29374 1764 29426
rect 1708 27076 1764 29374
rect 2492 29316 2548 29326
rect 2492 29314 3108 29316
rect 2492 29262 2494 29314
rect 2546 29262 3108 29314
rect 2492 29260 3108 29262
rect 2492 29250 2548 29260
rect 3052 28530 3108 29260
rect 3612 29204 3668 35196
rect 3724 29316 3780 39340
rect 3836 37268 3892 50372
rect 3948 45892 4004 54012
rect 4060 53060 4116 55244
rect 4172 55234 4228 55244
rect 4620 55074 4676 55086
rect 4620 55022 4622 55074
rect 4674 55022 4676 55074
rect 4172 54404 4228 54414
rect 4620 54404 4676 55022
rect 4172 54402 4340 54404
rect 4172 54350 4174 54402
rect 4226 54350 4340 54402
rect 4172 54348 4340 54350
rect 4172 54338 4228 54348
rect 4284 53396 4340 54348
rect 4620 54310 4676 54348
rect 4476 54124 4740 54134
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4476 54058 4740 54068
rect 4844 53844 4900 53854
rect 4844 53750 4900 53788
rect 4284 53340 4676 53396
rect 4060 52994 4116 53004
rect 4620 53172 4676 53340
rect 4956 53284 5012 81004
rect 5628 81284 5684 81294
rect 5628 79492 5684 81228
rect 5852 81282 5908 81340
rect 5852 81230 5854 81282
rect 5906 81230 5908 81282
rect 5852 81218 5908 81230
rect 6524 81170 6580 81340
rect 6524 81118 6526 81170
rect 6578 81118 6580 81170
rect 6524 81106 6580 81118
rect 6972 81340 7084 81396
rect 6076 79714 6132 79726
rect 6076 79662 6078 79714
rect 6130 79662 6132 79714
rect 5964 79602 6020 79614
rect 5964 79550 5966 79602
rect 6018 79550 6020 79602
rect 5964 79492 6020 79550
rect 5628 79490 5964 79492
rect 5628 79438 5630 79490
rect 5682 79438 5964 79490
rect 5628 79436 5964 79438
rect 5628 79426 5684 79436
rect 5964 79426 6020 79436
rect 5964 78932 6020 78942
rect 5964 78706 6020 78876
rect 5964 78654 5966 78706
rect 6018 78654 6020 78706
rect 5964 78596 6020 78654
rect 5628 78540 6020 78596
rect 5628 76020 5684 78540
rect 6076 78484 6132 79662
rect 6300 79602 6356 79614
rect 6300 79550 6302 79602
rect 6354 79550 6356 79602
rect 6300 78818 6356 79550
rect 6300 78766 6302 78818
rect 6354 78766 6356 78818
rect 6300 78754 6356 78766
rect 6860 79490 6916 79502
rect 6860 79438 6862 79490
rect 6914 79438 6916 79490
rect 6860 78820 6916 79438
rect 6860 78754 6916 78764
rect 6524 78708 6580 78718
rect 6524 78614 6580 78652
rect 6300 78596 6356 78606
rect 6076 78418 6132 78428
rect 6188 78594 6356 78596
rect 6188 78542 6302 78594
rect 6354 78542 6356 78594
rect 6188 78540 6356 78542
rect 5740 77924 5796 77934
rect 6188 77924 6244 78540
rect 6300 78530 6356 78540
rect 6972 78260 7028 81340
rect 7084 81302 7140 81340
rect 7196 79490 7252 81676
rect 7196 79438 7198 79490
rect 7250 79438 7252 79490
rect 7084 78932 7140 78942
rect 7196 78932 7252 79438
rect 7140 78876 7252 78932
rect 7420 81730 7476 81742
rect 7420 81678 7422 81730
rect 7474 81678 7476 81730
rect 7420 81172 7476 81678
rect 8988 81396 9044 82684
rect 8988 81330 9044 81340
rect 9548 81172 9604 82686
rect 9660 82964 9716 82974
rect 9660 82626 9716 82908
rect 10220 82852 10276 82862
rect 10220 82758 10276 82796
rect 9660 82574 9662 82626
rect 9714 82574 9716 82626
rect 9660 82562 9716 82574
rect 9772 82738 9828 82750
rect 9772 82686 9774 82738
rect 9826 82686 9828 82738
rect 9772 82628 9828 82686
rect 9772 82562 9828 82572
rect 9996 82738 10052 82750
rect 9996 82686 9998 82738
rect 10050 82686 10052 82738
rect 9660 81844 9716 81854
rect 9660 81750 9716 81788
rect 9884 81396 9940 81406
rect 9884 81302 9940 81340
rect 9660 81172 9716 81182
rect 9548 81170 9716 81172
rect 9548 81118 9662 81170
rect 9714 81118 9716 81170
rect 9548 81116 9716 81118
rect 7084 78866 7140 78876
rect 6524 78258 7028 78260
rect 6524 78206 6974 78258
rect 7026 78206 7028 78258
rect 6524 78204 7028 78206
rect 6524 78034 6580 78204
rect 6524 77982 6526 78034
rect 6578 77982 6580 78034
rect 6524 77970 6580 77982
rect 5740 77922 6244 77924
rect 5740 77870 5742 77922
rect 5794 77870 6244 77922
rect 5740 77868 6244 77870
rect 5740 77858 5796 77868
rect 6860 77476 6916 77486
rect 6860 76132 6916 77420
rect 6972 77364 7028 78204
rect 7308 78596 7364 78606
rect 7308 77476 7364 78540
rect 7028 77308 7252 77364
rect 6972 77298 7028 77308
rect 6860 76076 7028 76132
rect 5964 76020 6020 76030
rect 5628 75964 5964 76020
rect 5964 75682 6020 75964
rect 6860 75908 6916 75918
rect 6860 75796 6916 75852
rect 6524 75794 6916 75796
rect 6524 75742 6862 75794
rect 6914 75742 6916 75794
rect 6524 75740 6916 75742
rect 5964 75630 5966 75682
rect 6018 75630 6020 75682
rect 5964 75618 6020 75630
rect 6300 75684 6356 75694
rect 6300 75590 6356 75628
rect 6524 75682 6580 75740
rect 6860 75730 6916 75740
rect 6524 75630 6526 75682
rect 6578 75630 6580 75682
rect 6524 75618 6580 75630
rect 6076 75570 6132 75582
rect 6972 75572 7028 76076
rect 6076 75518 6078 75570
rect 6130 75518 6132 75570
rect 5292 74340 5348 74350
rect 5068 74116 5124 74126
rect 5292 74116 5348 74284
rect 5068 74114 5348 74116
rect 5068 74062 5070 74114
rect 5122 74062 5348 74114
rect 5068 74060 5348 74062
rect 5068 74050 5124 74060
rect 5292 73554 5348 74060
rect 5740 74114 5796 74126
rect 5740 74062 5742 74114
rect 5794 74062 5796 74114
rect 5740 73892 5796 74062
rect 6076 74114 6132 75518
rect 6860 75516 7028 75572
rect 6524 74788 6580 74798
rect 6524 74694 6580 74732
rect 6076 74062 6078 74114
rect 6130 74062 6132 74114
rect 6076 74050 6132 74062
rect 6636 74114 6692 74126
rect 6636 74062 6638 74114
rect 6690 74062 6692 74114
rect 5852 74004 5908 74042
rect 5852 73938 5908 73948
rect 5740 73826 5796 73836
rect 6188 73892 6244 73902
rect 5292 73502 5294 73554
rect 5346 73502 5348 73554
rect 5292 73490 5348 73502
rect 6188 73554 6244 73836
rect 6636 73892 6692 74062
rect 6748 74116 6804 74126
rect 6748 74002 6804 74060
rect 6748 73950 6750 74002
rect 6802 73950 6804 74002
rect 6748 73938 6804 73950
rect 6636 73826 6692 73836
rect 6188 73502 6190 73554
rect 6242 73502 6244 73554
rect 6188 73490 6244 73502
rect 6748 70978 6804 70990
rect 6748 70926 6750 70978
rect 6802 70926 6804 70978
rect 5628 70866 5684 70878
rect 5628 70814 5630 70866
rect 5682 70814 5684 70866
rect 5516 70194 5572 70206
rect 5516 70142 5518 70194
rect 5570 70142 5572 70194
rect 5068 69522 5124 69534
rect 5068 69470 5070 69522
rect 5122 69470 5124 69522
rect 5068 68852 5124 69470
rect 5068 68786 5124 68796
rect 5292 69188 5348 69198
rect 5292 68402 5348 69132
rect 5516 68964 5572 70142
rect 5628 69634 5684 70814
rect 5964 70756 6020 70766
rect 5964 70754 6244 70756
rect 5964 70702 5966 70754
rect 6018 70702 6244 70754
rect 5964 70700 6244 70702
rect 5964 70690 6020 70700
rect 6188 70306 6244 70700
rect 6188 70254 6190 70306
rect 6242 70254 6244 70306
rect 6188 70242 6244 70254
rect 5628 69582 5630 69634
rect 5682 69582 5684 69634
rect 5628 69570 5684 69582
rect 6748 70084 6804 70926
rect 6748 69634 6804 70028
rect 6748 69582 6750 69634
rect 6802 69582 6804 69634
rect 6748 69570 6804 69582
rect 5964 69410 6020 69422
rect 5964 69358 5966 69410
rect 6018 69358 6020 69410
rect 5964 69188 6020 69358
rect 5964 69122 6020 69132
rect 6188 69410 6244 69422
rect 6188 69358 6190 69410
rect 6242 69358 6244 69410
rect 5516 68898 5572 68908
rect 6076 68964 6132 68974
rect 5292 68350 5294 68402
rect 5346 68350 5348 68402
rect 5068 66948 5124 66958
rect 5068 66854 5124 66892
rect 5068 66388 5124 66398
rect 5068 66294 5124 66332
rect 5292 64484 5348 68350
rect 5068 62244 5124 62282
rect 5068 59778 5124 62188
rect 5292 60674 5348 64428
rect 5292 60622 5294 60674
rect 5346 60622 5348 60674
rect 5292 60564 5348 60622
rect 5628 68628 5684 68638
rect 5628 67620 5684 68572
rect 6076 68626 6132 68908
rect 6076 68574 6078 68626
rect 6130 68574 6132 68626
rect 5740 67620 5796 67630
rect 5628 67618 5796 67620
rect 5628 67566 5742 67618
rect 5794 67566 5796 67618
rect 5628 67564 5796 67566
rect 5628 60676 5684 67564
rect 5740 67554 5796 67564
rect 5852 66948 5908 66958
rect 6076 66948 6132 68574
rect 6188 68852 6244 69358
rect 6636 69188 6692 69198
rect 6636 69094 6692 69132
rect 6860 68964 6916 75516
rect 7196 74898 7252 77308
rect 7308 77362 7364 77420
rect 7308 77310 7310 77362
rect 7362 77310 7364 77362
rect 7308 77298 7364 77310
rect 7196 74846 7198 74898
rect 7250 74846 7252 74898
rect 7084 74452 7140 74462
rect 6972 74396 7084 74452
rect 6972 74114 7028 74396
rect 7084 74386 7140 74396
rect 7196 74340 7252 74846
rect 7308 76020 7364 76030
rect 7308 75458 7364 75964
rect 7308 75406 7310 75458
rect 7362 75406 7364 75458
rect 7308 74900 7364 75406
rect 7308 74834 7364 74844
rect 7196 74246 7252 74284
rect 6972 74062 6974 74114
rect 7026 74062 7028 74114
rect 6972 74050 7028 74062
rect 7308 74114 7364 74126
rect 7308 74062 7310 74114
rect 7362 74062 7364 74114
rect 7196 74004 7252 74014
rect 7308 74004 7364 74062
rect 7252 73948 7364 74004
rect 7196 73938 7252 73948
rect 7420 72324 7476 81116
rect 8988 81058 9044 81070
rect 8988 81006 8990 81058
rect 9042 81006 9044 81058
rect 8988 79492 9044 81006
rect 8988 79426 9044 79436
rect 9660 79492 9716 81116
rect 9772 81172 9828 81182
rect 9772 81078 9828 81116
rect 9996 81170 10052 82686
rect 12012 82738 12068 82750
rect 12012 82686 12014 82738
rect 12066 82686 12068 82738
rect 10668 82626 10724 82638
rect 10668 82574 10670 82626
rect 10722 82574 10724 82626
rect 10668 82516 10724 82574
rect 11116 82626 11172 82638
rect 11116 82574 11118 82626
rect 11170 82574 11172 82626
rect 10668 82450 10724 82460
rect 11004 82516 11060 82526
rect 10444 82404 10500 82414
rect 10444 81954 10500 82348
rect 10444 81902 10446 81954
rect 10498 81902 10500 81954
rect 10220 81284 10276 81294
rect 10220 81190 10276 81228
rect 9996 81118 9998 81170
rect 10050 81118 10052 81170
rect 9996 81060 10052 81118
rect 9996 80994 10052 81004
rect 10444 79604 10500 81902
rect 10780 81842 10836 81854
rect 10780 81790 10782 81842
rect 10834 81790 10836 81842
rect 10780 81396 10836 81790
rect 10892 81844 10948 81854
rect 10892 81750 10948 81788
rect 11004 81842 11060 82460
rect 11004 81790 11006 81842
rect 11058 81790 11060 81842
rect 11004 81778 11060 81790
rect 10780 81330 10836 81340
rect 10668 81060 10724 81070
rect 11116 81060 11172 82574
rect 11564 82404 11620 82414
rect 11564 82066 11620 82348
rect 12012 82404 12068 82686
rect 12572 82404 12628 84140
rect 12684 83300 12740 83310
rect 12684 82850 12740 83244
rect 12684 82798 12686 82850
rect 12738 82798 12740 82850
rect 12684 82786 12740 82798
rect 13020 83298 13076 83310
rect 13020 83246 13022 83298
rect 13074 83246 13076 83298
rect 12572 82348 12740 82404
rect 12012 82338 12068 82348
rect 11564 82014 11566 82066
rect 11618 82014 11620 82066
rect 11564 82002 11620 82014
rect 12572 81060 12628 81070
rect 10724 81004 11172 81060
rect 12236 81058 12628 81060
rect 12236 81006 12574 81058
rect 12626 81006 12628 81058
rect 12236 81004 12628 81006
rect 10668 80966 10724 81004
rect 10556 79604 10612 79614
rect 10444 79548 10556 79604
rect 10556 79510 10612 79548
rect 7532 78820 7588 78830
rect 7532 74676 7588 78764
rect 8876 78706 8932 78718
rect 8876 78654 8878 78706
rect 8930 78654 8932 78706
rect 8876 77924 8932 78654
rect 9548 78036 9604 78046
rect 9436 78034 9604 78036
rect 9436 77982 9550 78034
rect 9602 77982 9604 78034
rect 9436 77980 9604 77982
rect 8988 77924 9044 77934
rect 9436 77924 9492 77980
rect 9548 77970 9604 77980
rect 8876 77922 9492 77924
rect 8876 77870 8990 77922
rect 9042 77870 9492 77922
rect 8876 77868 9492 77870
rect 9660 77924 9716 79436
rect 10108 78932 10164 78942
rect 9884 78930 10164 78932
rect 9884 78878 10110 78930
rect 10162 78878 10164 78930
rect 9884 78876 10164 78878
rect 9884 78146 9940 78876
rect 10108 78866 10164 78876
rect 10668 78932 10724 78942
rect 10668 78818 10724 78876
rect 10668 78766 10670 78818
rect 10722 78766 10724 78818
rect 10668 78754 10724 78766
rect 10108 78596 10164 78606
rect 9884 78094 9886 78146
rect 9938 78094 9940 78146
rect 9884 78082 9940 78094
rect 9996 78594 10164 78596
rect 9996 78542 10110 78594
rect 10162 78542 10164 78594
rect 9996 78540 10164 78542
rect 9996 77924 10052 78540
rect 10108 78530 10164 78540
rect 10220 78596 10276 78606
rect 10220 78502 10276 78540
rect 10444 78594 10500 78606
rect 10444 78542 10446 78594
rect 10498 78542 10500 78594
rect 10444 78484 10500 78542
rect 10780 78484 10836 81004
rect 11900 80274 11956 80286
rect 11900 80222 11902 80274
rect 11954 80222 11956 80274
rect 11564 80164 11620 80174
rect 11340 80162 11620 80164
rect 11340 80110 11566 80162
rect 11618 80110 11620 80162
rect 11340 80108 11620 80110
rect 11340 79714 11396 80108
rect 11564 80098 11620 80108
rect 11340 79662 11342 79714
rect 11394 79662 11396 79714
rect 11340 79650 11396 79662
rect 11564 79604 11620 79614
rect 11452 79548 11564 79604
rect 11116 78594 11172 78606
rect 11116 78542 11118 78594
rect 11170 78542 11172 78594
rect 11116 78484 11172 78542
rect 10444 78428 11172 78484
rect 9660 77868 10052 77924
rect 8316 76580 8372 76590
rect 7644 76468 7700 76478
rect 7644 75796 7700 76412
rect 8316 76356 8372 76524
rect 7644 75702 7700 75740
rect 8204 76354 8372 76356
rect 8204 76302 8318 76354
rect 8370 76302 8372 76354
rect 8204 76300 8372 76302
rect 7756 74900 7812 74910
rect 7756 74806 7812 74844
rect 7868 74898 7924 74910
rect 7868 74846 7870 74898
rect 7922 74846 7924 74898
rect 7532 74620 7700 74676
rect 7644 73948 7700 74620
rect 7868 74452 7924 74846
rect 8092 74788 8148 74798
rect 8092 74694 8148 74732
rect 7868 74386 7924 74396
rect 7756 74338 7812 74350
rect 7756 74286 7758 74338
rect 7810 74286 7812 74338
rect 7756 74226 7812 74286
rect 7756 74174 7758 74226
rect 7810 74174 7812 74226
rect 7756 74162 7812 74174
rect 7420 72258 7476 72268
rect 7532 73892 7700 73948
rect 7980 74004 8036 74014
rect 8204 74004 8260 76300
rect 8316 76290 8372 76300
rect 8764 76580 8820 76590
rect 8988 76580 9044 77868
rect 9548 77812 9604 77822
rect 9436 77810 9604 77812
rect 9436 77758 9550 77810
rect 9602 77758 9604 77810
rect 9436 77756 9604 77758
rect 9436 77362 9492 77756
rect 9548 77746 9604 77756
rect 9436 77310 9438 77362
rect 9490 77310 9492 77362
rect 9436 77298 9492 77310
rect 8764 76578 9044 76580
rect 8764 76526 8766 76578
rect 8818 76526 9044 76578
rect 8764 76524 9044 76526
rect 9548 76580 9604 76590
rect 9660 76580 9716 77868
rect 10108 77252 10164 77262
rect 10668 77252 10724 77262
rect 10164 77250 10724 77252
rect 10164 77198 10670 77250
rect 10722 77198 10724 77250
rect 10164 77196 10724 77198
rect 10108 77158 10164 77196
rect 9604 76524 9716 76580
rect 8764 76244 8820 76524
rect 9548 76466 9604 76524
rect 9548 76414 9550 76466
rect 9602 76414 9604 76466
rect 9548 76402 9604 76414
rect 9772 76468 9828 76478
rect 9772 76374 9828 76412
rect 9996 76466 10052 76478
rect 9996 76414 9998 76466
rect 10050 76414 10052 76466
rect 8428 76188 8764 76244
rect 8316 75012 8372 75022
rect 8316 74898 8372 74956
rect 8316 74846 8318 74898
rect 8370 74846 8372 74898
rect 8316 74834 8372 74846
rect 8428 74900 8484 76188
rect 8764 76178 8820 76188
rect 8876 76354 8932 76366
rect 8876 76302 8878 76354
rect 8930 76302 8932 76354
rect 8876 76020 8932 76302
rect 9884 76354 9940 76366
rect 9884 76302 9886 76354
rect 9938 76302 9940 76354
rect 8988 76244 9044 76254
rect 9884 76244 9940 76302
rect 8988 76242 9940 76244
rect 8988 76190 8990 76242
rect 9042 76190 9940 76242
rect 8988 76188 9940 76190
rect 9996 76244 10052 76414
rect 10220 76468 10276 76478
rect 10220 76374 10276 76412
rect 10332 76356 10388 76366
rect 10332 76244 10388 76300
rect 9996 76188 10388 76244
rect 8988 76178 9044 76188
rect 8876 75964 9828 76020
rect 9772 75794 9828 75964
rect 9772 75742 9774 75794
rect 9826 75742 9828 75794
rect 9772 75730 9828 75742
rect 8764 75012 8820 75022
rect 8764 74918 8820 74956
rect 8428 74226 8484 74844
rect 8428 74174 8430 74226
rect 8482 74174 8484 74226
rect 8428 74162 8484 74174
rect 8036 73948 8260 74004
rect 10332 73948 10388 76188
rect 10444 75796 10500 77196
rect 10668 77186 10724 77196
rect 10668 76356 10724 76366
rect 10780 76356 10836 78428
rect 11116 78260 11172 78428
rect 11116 78194 11172 78204
rect 11340 77924 11396 77934
rect 10724 76300 10836 76356
rect 11116 76356 11172 76366
rect 10668 76262 10724 76300
rect 11116 76262 11172 76300
rect 11004 75796 11060 75806
rect 10444 75794 11060 75796
rect 10444 75742 11006 75794
rect 11058 75742 11060 75794
rect 10444 75740 11060 75742
rect 10444 75682 10500 75740
rect 10444 75630 10446 75682
rect 10498 75630 10500 75682
rect 10444 75618 10500 75630
rect 10892 74676 10948 75740
rect 11004 75730 11060 75740
rect 11340 74898 11396 77868
rect 11452 76466 11508 79548
rect 11564 79538 11620 79548
rect 11900 79042 11956 80222
rect 11900 78990 11902 79042
rect 11954 78990 11956 79042
rect 11900 78978 11956 78990
rect 12236 78930 12292 81004
rect 12572 80994 12628 81004
rect 12236 78878 12238 78930
rect 12290 78878 12292 78930
rect 12236 78866 12292 78878
rect 11564 78820 11620 78830
rect 11564 78726 11620 78764
rect 12460 78820 12516 78830
rect 12460 78726 12516 78764
rect 12124 77364 12180 77374
rect 12684 77364 12740 82348
rect 13020 81730 13076 83246
rect 13580 83300 13636 85932
rect 14140 85874 14196 86492
rect 14140 85822 14142 85874
rect 14194 85822 14196 85874
rect 13804 85764 13860 85774
rect 14140 85764 14196 85822
rect 13692 85762 14196 85764
rect 13692 85710 13806 85762
rect 13858 85710 14196 85762
rect 13692 85708 14196 85710
rect 14252 85762 14308 85774
rect 14252 85710 14254 85762
rect 14306 85710 14308 85762
rect 13692 85092 13748 85708
rect 13804 85698 13860 85708
rect 13692 84196 13748 85036
rect 14028 85316 14084 85326
rect 14028 85090 14084 85260
rect 14028 85038 14030 85090
rect 14082 85038 14084 85090
rect 14028 85026 14084 85038
rect 14252 85090 14308 85710
rect 15484 85708 15540 87388
rect 15596 87350 15652 87388
rect 15708 87220 15764 87230
rect 15708 87218 15876 87220
rect 15708 87166 15710 87218
rect 15762 87166 15876 87218
rect 15708 87164 15876 87166
rect 15708 87154 15764 87164
rect 15820 86660 15876 87164
rect 15820 86594 15876 86604
rect 14476 85652 14532 85662
rect 15148 85652 15540 85708
rect 14476 85650 14868 85652
rect 14476 85598 14478 85650
rect 14530 85598 14868 85650
rect 14476 85596 14868 85598
rect 14476 85586 14532 85596
rect 14812 85314 14868 85596
rect 14812 85262 14814 85314
rect 14866 85262 14868 85314
rect 14252 85038 14254 85090
rect 14306 85038 14308 85090
rect 14252 85026 14308 85038
rect 14588 85092 14644 85102
rect 14588 84998 14644 85036
rect 13804 84868 13860 84878
rect 14140 84868 14196 84878
rect 13860 84812 13972 84868
rect 13804 84774 13860 84812
rect 13692 84130 13748 84140
rect 13916 84532 13972 84812
rect 14140 84866 14756 84868
rect 14140 84814 14142 84866
rect 14194 84814 14756 84866
rect 14140 84812 14756 84814
rect 14140 84802 14196 84812
rect 13804 83412 13860 83422
rect 13692 83300 13748 83310
rect 13804 83300 13860 83356
rect 13580 83298 13860 83300
rect 13580 83246 13694 83298
rect 13746 83246 13860 83298
rect 13580 83244 13860 83246
rect 13692 83234 13748 83244
rect 13020 81678 13022 81730
rect 13074 81678 13076 81730
rect 13020 81172 13076 81678
rect 13692 81954 13748 81966
rect 13692 81902 13694 81954
rect 13746 81902 13748 81954
rect 13692 81396 13748 81902
rect 13244 81172 13300 81182
rect 13020 81170 13300 81172
rect 13020 81118 13246 81170
rect 13298 81118 13300 81170
rect 13020 81116 13300 81118
rect 13244 80948 13300 81116
rect 13468 81172 13524 81182
rect 13692 81172 13748 81340
rect 13468 81170 13748 81172
rect 13468 81118 13470 81170
rect 13522 81118 13748 81170
rect 13468 81116 13748 81118
rect 13468 81106 13524 81116
rect 13468 80948 13524 80958
rect 13244 80892 13468 80948
rect 13468 79490 13524 80892
rect 13468 79438 13470 79490
rect 13522 79438 13524 79490
rect 13468 78596 13524 79438
rect 13468 78530 13524 78540
rect 13580 79604 13636 79614
rect 13356 78036 13412 78046
rect 13580 78036 13636 79548
rect 13356 78034 13636 78036
rect 13356 77982 13358 78034
rect 13410 77982 13636 78034
rect 13356 77980 13636 77982
rect 13356 77970 13412 77980
rect 12908 77924 12964 77934
rect 13804 77924 13860 83244
rect 12908 77830 12964 77868
rect 13580 77868 13860 77924
rect 13916 77924 13972 84476
rect 14700 84418 14756 84812
rect 14700 84366 14702 84418
rect 14754 84366 14756 84418
rect 14700 84354 14756 84366
rect 14812 83748 14868 85262
rect 15148 85316 15204 85652
rect 15148 85222 15204 85260
rect 15596 85092 15652 85102
rect 15596 84998 15652 85036
rect 15484 84306 15540 84318
rect 15484 84254 15486 84306
rect 15538 84254 15540 84306
rect 15484 84196 15540 84254
rect 15932 84196 15988 88172
rect 16156 88162 16212 88172
rect 15484 84194 15988 84196
rect 15484 84142 15934 84194
rect 15986 84142 15988 84194
rect 15484 84140 15988 84142
rect 14812 83746 15428 83748
rect 14812 83694 14814 83746
rect 14866 83694 15428 83746
rect 14812 83692 15428 83694
rect 14812 83682 14868 83692
rect 15372 83522 15428 83692
rect 15372 83470 15374 83522
rect 15426 83470 15428 83522
rect 15372 83458 15428 83470
rect 14140 83410 14196 83422
rect 14140 83358 14142 83410
rect 14194 83358 14196 83410
rect 14140 82964 14196 83358
rect 14028 82516 14084 82526
rect 14028 81730 14084 82460
rect 14028 81678 14030 81730
rect 14082 81678 14084 81730
rect 14028 81666 14084 81678
rect 14140 81842 14196 82908
rect 14140 81790 14142 81842
rect 14194 81790 14196 81842
rect 14028 81060 14084 81070
rect 14140 81060 14196 81790
rect 14252 83410 14308 83422
rect 14252 83358 14254 83410
rect 14306 83358 14308 83410
rect 14252 81844 14308 83358
rect 14364 83412 14420 83422
rect 14364 83410 14532 83412
rect 14364 83358 14366 83410
rect 14418 83358 14532 83410
rect 14364 83356 14532 83358
rect 14364 83346 14420 83356
rect 14476 82178 14532 83356
rect 15148 83298 15204 83310
rect 15148 83246 15150 83298
rect 15202 83246 15204 83298
rect 14476 82126 14478 82178
rect 14530 82126 14532 82178
rect 14476 82114 14532 82126
rect 14812 83076 14868 83086
rect 14812 82626 14868 83020
rect 14812 82574 14814 82626
rect 14866 82574 14868 82626
rect 14364 81844 14420 81854
rect 14252 81842 14420 81844
rect 14252 81790 14366 81842
rect 14418 81790 14420 81842
rect 14252 81788 14420 81790
rect 14364 81732 14420 81788
rect 14812 81732 14868 82574
rect 15148 82516 15204 83246
rect 15260 83300 15316 83310
rect 15260 83206 15316 83244
rect 15148 82450 15204 82460
rect 15372 83188 15428 83198
rect 14364 81730 14868 81732
rect 14364 81678 14814 81730
rect 14866 81678 14868 81730
rect 14364 81676 14868 81678
rect 14476 81396 14532 81406
rect 14476 81302 14532 81340
rect 14028 81058 14196 81060
rect 14028 81006 14030 81058
rect 14082 81006 14196 81058
rect 14028 81004 14196 81006
rect 14028 80948 14084 81004
rect 14028 80882 14084 80892
rect 14812 79828 14868 81676
rect 14924 82178 14980 82190
rect 14924 82126 14926 82178
rect 14978 82126 14980 82178
rect 14924 81396 14980 82126
rect 15372 82178 15428 83132
rect 15484 82626 15540 84140
rect 15932 84130 15988 84140
rect 16044 87668 16100 87678
rect 16044 86770 16100 87612
rect 16268 87442 16324 88844
rect 16716 88786 16772 88798
rect 16716 88734 16718 88786
rect 16770 88734 16772 88786
rect 16716 88340 16772 88734
rect 16716 88274 16772 88284
rect 16716 87668 16772 87678
rect 16716 87554 16772 87612
rect 16716 87502 16718 87554
rect 16770 87502 16772 87554
rect 16716 87490 16772 87502
rect 16268 87390 16270 87442
rect 16322 87390 16324 87442
rect 16268 87378 16324 87390
rect 16044 86718 16046 86770
rect 16098 86718 16100 86770
rect 15596 83412 15652 83422
rect 15596 83318 15652 83356
rect 15484 82574 15486 82626
rect 15538 82574 15540 82626
rect 15484 82292 15540 82574
rect 15484 82226 15540 82236
rect 15372 82126 15374 82178
rect 15426 82126 15428 82178
rect 15260 82068 15316 82078
rect 15372 82068 15428 82126
rect 15260 82066 15428 82068
rect 15260 82014 15262 82066
rect 15314 82014 15428 82066
rect 15260 82012 15428 82014
rect 15260 82002 15316 82012
rect 14924 81330 14980 81340
rect 15372 79828 15428 79838
rect 14812 79826 15428 79828
rect 14812 79774 15374 79826
rect 15426 79774 15428 79826
rect 14812 79772 15428 79774
rect 14140 79604 14196 79614
rect 14140 79510 14196 79548
rect 14588 78820 14644 78830
rect 14028 78764 14532 78820
rect 14028 78146 14084 78764
rect 14364 78596 14420 78606
rect 14028 78094 14030 78146
rect 14082 78094 14084 78146
rect 14028 78082 14084 78094
rect 14252 78594 14420 78596
rect 14252 78542 14366 78594
rect 14418 78542 14420 78594
rect 14252 78540 14420 78542
rect 14476 78596 14532 78764
rect 14588 78818 14868 78820
rect 14588 78766 14590 78818
rect 14642 78766 14868 78818
rect 14588 78764 14868 78766
rect 14588 78754 14644 78764
rect 14700 78596 14756 78606
rect 14476 78594 14756 78596
rect 14476 78542 14702 78594
rect 14754 78542 14756 78594
rect 14476 78540 14756 78542
rect 14140 77924 14196 77934
rect 14252 77924 14308 78540
rect 14364 78530 14420 78540
rect 14700 78530 14756 78540
rect 13916 77868 14084 77924
rect 12124 77362 12740 77364
rect 12124 77310 12126 77362
rect 12178 77310 12740 77362
rect 12124 77308 12740 77310
rect 12908 77364 12964 77374
rect 12124 77298 12180 77308
rect 12572 77250 12628 77308
rect 12572 77198 12574 77250
rect 12626 77198 12628 77250
rect 12572 77186 12628 77198
rect 12908 77250 12964 77308
rect 12908 77198 12910 77250
rect 12962 77198 12964 77250
rect 12908 77186 12964 77198
rect 12348 77140 12404 77150
rect 12348 77046 12404 77084
rect 12460 77026 12516 77038
rect 12460 76974 12462 77026
rect 12514 76974 12516 77026
rect 12460 76692 12516 76974
rect 12236 76636 12516 76692
rect 12236 76578 12292 76636
rect 12236 76526 12238 76578
rect 12290 76526 12292 76578
rect 12236 76514 12292 76526
rect 11452 76414 11454 76466
rect 11506 76414 11508 76466
rect 11452 76402 11508 76414
rect 11340 74846 11342 74898
rect 11394 74846 11396 74898
rect 10892 74610 10948 74620
rect 11004 74788 11060 74798
rect 11340 74788 11396 74846
rect 11004 74786 11396 74788
rect 11004 74734 11006 74786
rect 11058 74734 11396 74786
rect 11004 74732 11396 74734
rect 13468 76356 13524 76366
rect 11004 73948 11060 74732
rect 7532 72100 7588 73892
rect 7196 72044 7588 72100
rect 6188 68292 6244 68796
rect 6188 68226 6244 68236
rect 6748 68908 6916 68964
rect 7084 69634 7140 69646
rect 7084 69582 7086 69634
rect 7138 69582 7140 69634
rect 7084 69186 7140 69582
rect 7084 69134 7086 69186
rect 7138 69134 7140 69186
rect 7084 68964 7140 69134
rect 5908 66892 6132 66948
rect 5852 66274 5908 66892
rect 5852 66222 5854 66274
rect 5906 66222 5908 66274
rect 5740 65378 5796 65390
rect 5740 65326 5742 65378
rect 5794 65326 5796 65378
rect 5740 62692 5796 65326
rect 5852 65380 5908 66222
rect 6524 66162 6580 66174
rect 6524 66110 6526 66162
rect 6578 66110 6580 66162
rect 6524 65492 6580 66110
rect 6524 65426 6580 65436
rect 6188 65380 6244 65390
rect 5852 65378 6244 65380
rect 5852 65326 6190 65378
rect 6242 65326 6244 65378
rect 5852 65324 6244 65326
rect 5740 62626 5796 62636
rect 6188 63700 6244 65324
rect 6748 64820 6804 68908
rect 7084 68898 7140 68908
rect 6860 68514 6916 68526
rect 6860 68462 6862 68514
rect 6914 68462 6916 68514
rect 6860 68180 6916 68462
rect 6860 68114 6916 68124
rect 7084 65602 7140 65614
rect 7084 65550 7086 65602
rect 7138 65550 7140 65602
rect 7084 65492 7140 65550
rect 7084 65426 7140 65436
rect 6748 64754 6804 64764
rect 5740 62356 5796 62366
rect 6188 62356 6244 63644
rect 6972 63812 7028 63822
rect 5740 62354 6244 62356
rect 5740 62302 5742 62354
rect 5794 62302 6244 62354
rect 5740 62300 6244 62302
rect 6412 63026 6468 63038
rect 6412 62974 6414 63026
rect 6466 62974 6468 63026
rect 5740 62244 5796 62300
rect 6412 62188 6468 62974
rect 6748 62916 6804 62926
rect 6524 62914 6804 62916
rect 6524 62862 6750 62914
rect 6802 62862 6804 62914
rect 6524 62860 6804 62862
rect 6524 62466 6580 62860
rect 6748 62850 6804 62860
rect 6524 62414 6526 62466
rect 6578 62414 6580 62466
rect 6524 62402 6580 62414
rect 6748 62692 6804 62702
rect 5740 62178 5796 62188
rect 6188 62132 6468 62188
rect 6188 61794 6244 62132
rect 6188 61742 6190 61794
rect 6242 61742 6244 61794
rect 6188 61730 6244 61742
rect 5964 61684 6020 61694
rect 5964 61590 6020 61628
rect 6524 61684 6580 61694
rect 6524 61590 6580 61628
rect 6748 61458 6804 62636
rect 6748 61406 6750 61458
rect 6802 61406 6804 61458
rect 5740 60900 5796 60938
rect 5740 60834 5796 60844
rect 6188 60788 6244 60798
rect 5628 60620 5796 60676
rect 5292 60498 5348 60508
rect 5740 59892 5796 60620
rect 5852 60004 5908 60014
rect 5852 59910 5908 59948
rect 5740 59826 5796 59836
rect 5068 59726 5070 59778
rect 5122 59726 5124 59778
rect 5068 59108 5124 59726
rect 5628 59780 5684 59790
rect 5628 59686 5684 59724
rect 5404 59108 5460 59118
rect 5068 59052 5404 59108
rect 5068 58434 5124 58446
rect 5068 58382 5070 58434
rect 5122 58382 5124 58434
rect 5068 58324 5124 58382
rect 5068 58258 5124 58268
rect 5068 57764 5124 57774
rect 5292 57764 5348 59052
rect 5404 59042 5460 59052
rect 6188 58324 6244 60732
rect 6300 60676 6356 60686
rect 6748 60676 6804 61406
rect 6860 60900 6916 60910
rect 6860 60806 6916 60844
rect 6972 60786 7028 63756
rect 7196 60900 7252 72044
rect 7532 71876 7588 71886
rect 7532 71090 7588 71820
rect 7532 71038 7534 71090
rect 7586 71038 7588 71090
rect 7532 71026 7588 71038
rect 7644 68180 7700 68190
rect 7700 68124 7924 68180
rect 7644 68114 7700 68124
rect 7868 67730 7924 68124
rect 7868 67678 7870 67730
rect 7922 67678 7924 67730
rect 7868 67666 7924 67678
rect 7420 65492 7476 65502
rect 7420 65490 7924 65492
rect 7420 65438 7422 65490
rect 7474 65438 7924 65490
rect 7420 65436 7924 65438
rect 7420 65426 7476 65436
rect 7868 64930 7924 65436
rect 7868 64878 7870 64930
rect 7922 64878 7924 64930
rect 7868 64866 7924 64878
rect 7532 64484 7588 64494
rect 7532 64390 7588 64428
rect 7980 62188 8036 73948
rect 10332 73892 10500 73948
rect 7868 62132 8036 62188
rect 8092 72324 8148 72334
rect 8092 62188 8148 72268
rect 8540 71876 8596 71886
rect 8540 71782 8596 71820
rect 8876 71764 8932 71774
rect 8876 71762 9156 71764
rect 8876 71710 8878 71762
rect 8930 71710 9156 71762
rect 8876 71708 9156 71710
rect 8876 71698 8932 71708
rect 8316 70082 8372 70094
rect 8316 70030 8318 70082
rect 8370 70030 8372 70082
rect 8316 69300 8372 70030
rect 8764 70084 8820 70094
rect 8764 69990 8820 70028
rect 9100 69634 9156 71708
rect 9996 71650 10052 71662
rect 9996 71598 9998 71650
rect 10050 71598 10052 71650
rect 9660 71090 9716 71102
rect 9660 71038 9662 71090
rect 9714 71038 9716 71090
rect 9100 69582 9102 69634
rect 9154 69582 9156 69634
rect 9100 69570 9156 69582
rect 9548 70868 9604 70878
rect 9548 70084 9604 70812
rect 9660 70644 9716 71038
rect 9996 70978 10052 71598
rect 9996 70926 9998 70978
rect 10050 70926 10052 70978
rect 9996 70868 10052 70926
rect 9996 70802 10052 70812
rect 9660 70588 10164 70644
rect 9884 70084 9940 70094
rect 9548 69522 9604 70028
rect 9548 69470 9550 69522
rect 9602 69470 9604 69522
rect 9548 69458 9604 69470
rect 9772 70028 9884 70084
rect 8764 69410 8820 69422
rect 8764 69358 8766 69410
rect 8818 69358 8820 69410
rect 8540 69300 8596 69310
rect 8316 69298 8596 69300
rect 8316 69246 8542 69298
rect 8594 69246 8596 69298
rect 8316 69244 8596 69246
rect 8204 67732 8260 67742
rect 8204 67730 8372 67732
rect 8204 67678 8206 67730
rect 8258 67678 8372 67730
rect 8204 67676 8372 67678
rect 8204 67666 8260 67676
rect 8316 66948 8372 67676
rect 8428 66948 8484 66958
rect 8316 66946 8484 66948
rect 8316 66894 8430 66946
rect 8482 66894 8484 66946
rect 8316 66892 8484 66894
rect 8428 66882 8484 66892
rect 8204 64706 8260 64718
rect 8204 64654 8206 64706
rect 8258 64654 8260 64706
rect 8204 64484 8260 64654
rect 8204 64418 8260 64428
rect 8428 64706 8484 64718
rect 8428 64654 8430 64706
rect 8482 64654 8484 64706
rect 8428 63364 8484 64654
rect 8428 63298 8484 63308
rect 8092 62132 8260 62188
rect 7644 61348 7700 61358
rect 7420 60900 7476 60910
rect 6972 60734 6974 60786
rect 7026 60734 7028 60786
rect 6972 60722 7028 60734
rect 7084 60898 7476 60900
rect 7084 60846 7422 60898
rect 7474 60846 7476 60898
rect 7084 60844 7476 60846
rect 6300 60674 6468 60676
rect 6300 60622 6302 60674
rect 6354 60622 6468 60674
rect 6300 60620 6468 60622
rect 6748 60620 6916 60676
rect 6300 60610 6356 60620
rect 5740 58212 5796 58222
rect 5068 57762 5684 57764
rect 5068 57710 5070 57762
rect 5122 57710 5684 57762
rect 5068 57708 5684 57710
rect 5068 57698 5124 57708
rect 5628 55300 5684 57708
rect 5740 57428 5796 58156
rect 6188 58210 6244 58268
rect 6188 58158 6190 58210
rect 6242 58158 6244 58210
rect 5740 57372 6020 57428
rect 5852 57204 5908 57214
rect 5740 55300 5796 55310
rect 5628 55298 5796 55300
rect 5628 55246 5742 55298
rect 5794 55246 5796 55298
rect 5628 55244 5796 55246
rect 5740 55234 5796 55244
rect 4956 53218 5012 53228
rect 5068 53844 5124 53854
rect 4620 52834 4676 53116
rect 4844 53060 4900 53070
rect 4900 53004 5012 53060
rect 4844 52994 4900 53004
rect 4620 52782 4622 52834
rect 4674 52782 4676 52834
rect 4620 52770 4676 52782
rect 4956 52946 5012 53004
rect 4956 52894 4958 52946
rect 5010 52894 5012 52946
rect 4476 52556 4740 52566
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4476 52490 4740 52500
rect 4844 52276 4900 52286
rect 4956 52276 5012 52894
rect 4844 52274 5012 52276
rect 4844 52222 4846 52274
rect 4898 52222 5012 52274
rect 4844 52220 5012 52222
rect 4844 52210 4900 52220
rect 5068 52164 5124 53788
rect 5852 53506 5908 57148
rect 5852 53454 5854 53506
rect 5906 53454 5908 53506
rect 5404 53172 5460 53182
rect 5404 53078 5460 53116
rect 5180 52948 5236 52958
rect 5180 52854 5236 52892
rect 5628 52948 5684 52958
rect 5852 52948 5908 53454
rect 5628 52946 5908 52948
rect 5628 52894 5630 52946
rect 5682 52894 5908 52946
rect 5628 52892 5908 52894
rect 5964 52948 6020 57372
rect 6188 57204 6244 58158
rect 6188 57138 6244 57148
rect 6188 55076 6244 55086
rect 6188 54514 6244 55020
rect 6188 54462 6190 54514
rect 6242 54462 6244 54514
rect 6188 53844 6244 54462
rect 6188 53778 6244 53788
rect 6300 53620 6356 53630
rect 6300 53170 6356 53564
rect 6300 53118 6302 53170
rect 6354 53118 6356 53170
rect 6300 53106 6356 53118
rect 6076 52948 6132 52958
rect 5964 52892 6076 52948
rect 4956 52052 5012 52062
rect 4844 51996 4956 52052
rect 4172 51380 4228 51390
rect 4172 51286 4228 51324
rect 4476 50988 4740 50998
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4476 50922 4740 50932
rect 4620 49698 4676 49710
rect 4620 49646 4622 49698
rect 4674 49646 4676 49698
rect 4620 49588 4676 49646
rect 4732 49588 4788 49598
rect 4620 49532 4732 49588
rect 4732 49522 4788 49532
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 4060 48244 4116 48254
rect 4732 48244 4788 48254
rect 4060 48242 4788 48244
rect 4060 48190 4062 48242
rect 4114 48190 4734 48242
rect 4786 48190 4788 48242
rect 4060 48188 4788 48190
rect 4060 48178 4116 48188
rect 4732 48178 4788 48188
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 4060 46060 4676 46116
rect 4060 45892 4116 46060
rect 4620 46002 4676 46060
rect 4620 45950 4622 46002
rect 4674 45950 4676 46002
rect 4620 45938 4676 45950
rect 3948 45890 4116 45892
rect 3948 45838 3950 45890
rect 4002 45838 4116 45890
rect 3948 45836 4116 45838
rect 4172 45890 4228 45902
rect 4172 45838 4174 45890
rect 4226 45838 4228 45890
rect 3948 44322 4004 45836
rect 4172 45332 4228 45838
rect 4172 45266 4228 45276
rect 4620 44994 4676 45006
rect 4620 44942 4622 44994
rect 4674 44942 4676 44994
rect 4620 44884 4676 44942
rect 4284 44828 4676 44884
rect 3948 44270 3950 44322
rect 4002 44270 4004 44322
rect 3948 43652 4004 44270
rect 3948 43586 4004 43596
rect 4172 44324 4228 44334
rect 4284 44324 4340 44828
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 4172 44322 4340 44324
rect 4172 44270 4174 44322
rect 4226 44270 4340 44322
rect 4172 44268 4340 44270
rect 3948 40404 4004 40414
rect 3948 40310 4004 40348
rect 4172 39620 4228 44268
rect 4844 44212 4900 51996
rect 4956 51986 5012 51996
rect 5068 51602 5124 52108
rect 5068 51550 5070 51602
rect 5122 51550 5124 51602
rect 5068 50036 5124 51550
rect 5292 52834 5348 52846
rect 5292 52782 5294 52834
rect 5346 52782 5348 52834
rect 5292 50428 5348 52782
rect 5628 52052 5684 52892
rect 6076 52164 6132 52892
rect 6076 52162 6244 52164
rect 6076 52110 6078 52162
rect 6130 52110 6244 52162
rect 6076 52108 6244 52110
rect 6076 52098 6132 52108
rect 5628 51986 5684 51996
rect 5292 50372 5460 50428
rect 5068 49942 5124 49980
rect 4956 49476 5012 49486
rect 4956 45332 5012 49420
rect 5292 48132 5348 48142
rect 5292 48038 5348 48076
rect 5068 48018 5124 48030
rect 5068 47966 5070 48018
rect 5122 47966 5124 48018
rect 5068 47796 5124 47966
rect 5068 47730 5124 47740
rect 5404 47684 5460 50372
rect 5964 50036 6020 50046
rect 5964 48244 6020 49980
rect 5964 48242 6132 48244
rect 5964 48190 5966 48242
rect 6018 48190 6132 48242
rect 5964 48188 6132 48190
rect 5964 48178 6020 48188
rect 5404 47628 6020 47684
rect 5068 47572 5124 47582
rect 5068 47570 5684 47572
rect 5068 47518 5070 47570
rect 5122 47518 5684 47570
rect 5068 47516 5684 47518
rect 5068 47506 5124 47516
rect 4956 45266 5012 45276
rect 5292 47348 5348 47358
rect 5292 47124 5348 47292
rect 5292 46562 5348 47068
rect 5292 46510 5294 46562
rect 5346 46510 5348 46562
rect 5068 44996 5124 45006
rect 5292 44996 5348 46510
rect 5068 44994 5348 44996
rect 5068 44942 5070 44994
rect 5122 44942 5348 44994
rect 5068 44940 5348 44942
rect 5068 44930 5124 44940
rect 4844 44146 4900 44156
rect 4620 44098 4676 44110
rect 4620 44046 4622 44098
rect 4674 44046 4676 44098
rect 4620 43988 4676 44046
rect 4620 43932 4900 43988
rect 4844 43652 4900 43932
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 4844 42756 4900 43596
rect 5180 43540 5236 44940
rect 5516 43540 5572 43550
rect 5180 43484 5516 43540
rect 5516 43446 5572 43484
rect 5068 43428 5124 43438
rect 5068 43426 5460 43428
rect 5068 43374 5070 43426
rect 5122 43374 5460 43426
rect 5068 43372 5460 43374
rect 5068 43362 5124 43372
rect 5404 42868 5460 43372
rect 5628 43092 5684 47516
rect 5740 47236 5796 47246
rect 5740 47142 5796 47180
rect 5628 43036 5796 43092
rect 5628 42868 5684 42878
rect 5404 42866 5684 42868
rect 5404 42814 5630 42866
rect 5682 42814 5684 42866
rect 5404 42812 5684 42814
rect 4844 42690 4900 42700
rect 5068 42756 5124 42766
rect 4956 41636 5012 41646
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 4508 40628 4564 40638
rect 4284 40516 4340 40526
rect 4284 40402 4340 40460
rect 4284 40350 4286 40402
rect 4338 40350 4340 40402
rect 4284 40338 4340 40350
rect 4508 40402 4564 40572
rect 4956 40516 5012 41580
rect 4956 40422 5012 40460
rect 4508 40350 4510 40402
rect 4562 40350 4564 40402
rect 4508 40338 4564 40350
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 5068 39844 5124 42700
rect 5516 42420 5572 42430
rect 5516 41860 5572 42364
rect 5628 42082 5684 42812
rect 5628 42030 5630 42082
rect 5682 42030 5684 42082
rect 5628 42018 5684 42030
rect 5516 41804 5684 41860
rect 4956 39788 5124 39844
rect 5292 41748 5348 41758
rect 4396 39620 4452 39630
rect 4172 39618 4452 39620
rect 4172 39566 4398 39618
rect 4450 39566 4452 39618
rect 4172 39564 4452 39566
rect 4396 39554 4452 39564
rect 4620 39394 4676 39406
rect 4620 39342 4622 39394
rect 4674 39342 4676 39394
rect 4620 39060 4676 39342
rect 4620 38994 4676 39004
rect 4732 39394 4788 39406
rect 4732 39342 4734 39394
rect 4786 39342 4788 39394
rect 4620 38722 4676 38734
rect 4620 38670 4622 38722
rect 4674 38670 4676 38722
rect 4620 38668 4676 38670
rect 4172 38612 4676 38668
rect 4732 38612 4788 39342
rect 4844 39394 4900 39406
rect 4844 39342 4846 39394
rect 4898 39342 4900 39394
rect 4844 38668 4900 39342
rect 4956 39396 5012 39788
rect 5068 39618 5124 39630
rect 5068 39566 5070 39618
rect 5122 39566 5124 39618
rect 5068 39508 5124 39566
rect 5180 39508 5236 39518
rect 5068 39452 5180 39508
rect 4956 39340 5124 39396
rect 5068 38836 5124 39340
rect 5180 39058 5236 39452
rect 5180 39006 5182 39058
rect 5234 39006 5236 39058
rect 5180 38994 5236 39006
rect 5180 38836 5236 38846
rect 5068 38780 5180 38836
rect 5180 38770 5236 38780
rect 4844 38612 5012 38668
rect 3836 37202 3892 37212
rect 3948 37716 4004 37726
rect 3948 35698 4004 37660
rect 4172 36708 4228 38612
rect 4732 38546 4788 38556
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 4844 38164 4900 38174
rect 4844 38070 4900 38108
rect 4620 38050 4676 38062
rect 4620 37998 4622 38050
rect 4674 37998 4676 38050
rect 4284 37828 4340 37838
rect 4284 37734 4340 37772
rect 4620 37828 4676 37998
rect 4620 37762 4676 37772
rect 4620 37156 4676 37166
rect 4172 36642 4228 36652
rect 4284 37154 4676 37156
rect 4284 37102 4622 37154
rect 4674 37102 4676 37154
rect 4284 37100 4676 37102
rect 4284 36372 4340 37100
rect 4620 37090 4676 37100
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4172 35812 4228 35822
rect 4284 35812 4340 36316
rect 4172 35810 4340 35812
rect 4172 35758 4174 35810
rect 4226 35758 4340 35810
rect 4172 35756 4340 35758
rect 4508 36708 4564 36718
rect 4172 35746 4228 35756
rect 3948 35646 3950 35698
rect 4002 35646 4004 35698
rect 3948 35140 4004 35646
rect 4508 35698 4564 36652
rect 4508 35646 4510 35698
rect 4562 35646 4564 35698
rect 4508 35634 4564 35646
rect 4732 35700 4788 35710
rect 4732 35606 4788 35644
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 3948 35084 4452 35140
rect 4396 35026 4452 35084
rect 4396 34974 4398 35026
rect 4450 34974 4452 35026
rect 4396 34962 4452 34974
rect 4956 34468 5012 38612
rect 5068 37828 5124 37838
rect 5068 37490 5124 37772
rect 5068 37438 5070 37490
rect 5122 37438 5124 37490
rect 5068 37426 5124 37438
rect 5180 37268 5236 37278
rect 5180 36594 5236 37212
rect 5180 36542 5182 36594
rect 5234 36542 5236 36594
rect 5180 36530 5236 36542
rect 5068 35476 5124 35486
rect 5068 35474 5236 35476
rect 5068 35422 5070 35474
rect 5122 35422 5236 35474
rect 5068 35420 5236 35422
rect 5068 35410 5124 35420
rect 4844 34412 5012 34468
rect 4620 34020 4676 34030
rect 4620 33926 4676 33964
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4732 33572 4788 33582
rect 4620 33570 4788 33572
rect 4620 33518 4734 33570
rect 4786 33518 4788 33570
rect 4620 33516 4788 33518
rect 3948 33124 4004 33134
rect 3948 32562 4004 33068
rect 4620 32674 4676 33516
rect 4732 33506 4788 33516
rect 4844 33348 4900 34412
rect 4956 34242 5012 34254
rect 4956 34190 4958 34242
rect 5010 34190 5012 34242
rect 4956 33570 5012 34190
rect 5180 34130 5236 35420
rect 5180 34078 5182 34130
rect 5234 34078 5236 34130
rect 5180 34066 5236 34078
rect 4956 33518 4958 33570
rect 5010 33518 5012 33570
rect 4956 33506 5012 33518
rect 4620 32622 4622 32674
rect 4674 32622 4676 32674
rect 4620 32610 4676 32622
rect 4732 33292 4900 33348
rect 3948 32510 3950 32562
rect 4002 32510 4004 32562
rect 3948 32452 4004 32510
rect 3836 30098 3892 30110
rect 3836 30046 3838 30098
rect 3890 30046 3892 30098
rect 3836 29652 3892 30046
rect 3836 29586 3892 29596
rect 3948 29540 4004 32396
rect 4732 32340 4788 33292
rect 4844 33124 4900 33134
rect 4844 33030 4900 33068
rect 4732 32284 4900 32340
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4844 30436 4900 32284
rect 5292 30882 5348 41692
rect 5404 40402 5460 40414
rect 5404 40350 5406 40402
rect 5458 40350 5460 40402
rect 5404 38164 5460 40350
rect 5628 40402 5684 41804
rect 5740 40628 5796 43036
rect 5852 42756 5908 42766
rect 5852 42662 5908 42700
rect 5852 42084 5908 42094
rect 5852 41990 5908 42028
rect 5964 41860 6020 47628
rect 6076 47458 6132 48188
rect 6076 47406 6078 47458
rect 6130 47406 6132 47458
rect 6076 47348 6132 47406
rect 6076 47282 6132 47292
rect 6188 46228 6244 52108
rect 6300 51380 6356 51390
rect 6300 50818 6356 51324
rect 6300 50766 6302 50818
rect 6354 50766 6356 50818
rect 6300 50754 6356 50766
rect 6188 46162 6244 46172
rect 6188 43540 6244 43550
rect 6244 43484 6356 43540
rect 6188 43446 6244 43484
rect 6188 42980 6244 42990
rect 6188 42886 6244 42924
rect 6300 42756 6356 43484
rect 6300 42690 6356 42700
rect 6076 41972 6132 41982
rect 6076 41878 6132 41916
rect 6300 41970 6356 41982
rect 6300 41918 6302 41970
rect 6354 41918 6356 41970
rect 5852 41804 6020 41860
rect 6188 41858 6244 41870
rect 6188 41806 6190 41858
rect 6242 41806 6244 41858
rect 5852 40740 5908 41804
rect 5852 40684 6132 40740
rect 5740 40516 5796 40572
rect 5852 40516 5908 40526
rect 5740 40514 5908 40516
rect 5740 40462 5854 40514
rect 5906 40462 5908 40514
rect 5740 40460 5908 40462
rect 5852 40450 5908 40460
rect 5628 40350 5630 40402
rect 5682 40350 5684 40402
rect 5628 40292 5684 40350
rect 5964 40404 6020 40414
rect 5964 40310 6020 40348
rect 5628 40226 5684 40236
rect 5740 40290 5796 40302
rect 5740 40238 5742 40290
rect 5794 40238 5796 40290
rect 5628 39620 5684 39630
rect 5628 39526 5684 39564
rect 5516 39060 5572 39070
rect 5516 38966 5572 39004
rect 5740 38836 5796 40238
rect 6076 40180 6132 40684
rect 5964 40124 6132 40180
rect 5852 39732 5908 39742
rect 5852 39618 5908 39676
rect 5852 39566 5854 39618
rect 5906 39566 5908 39618
rect 5852 39060 5908 39566
rect 5852 38994 5908 39004
rect 5964 38946 6020 40124
rect 6188 40068 6244 41806
rect 6300 41748 6356 41918
rect 6300 41682 6356 41692
rect 6412 40964 6468 60620
rect 6748 59106 6804 59118
rect 6748 59054 6750 59106
rect 6802 59054 6804 59106
rect 6748 58436 6804 59054
rect 6748 57988 6804 58380
rect 6860 58434 6916 60620
rect 6972 60116 7028 60126
rect 7084 60116 7140 60844
rect 7420 60834 7476 60844
rect 7532 60900 7588 60910
rect 7644 60900 7700 61292
rect 7588 60844 7700 60900
rect 6972 60114 7140 60116
rect 6972 60062 6974 60114
rect 7026 60062 7140 60114
rect 6972 60060 7140 60062
rect 6972 60050 7028 60060
rect 6860 58382 6862 58434
rect 6914 58382 6916 58434
rect 6860 58370 6916 58382
rect 6972 58994 7028 59006
rect 6972 58942 6974 58994
rect 7026 58942 7028 58994
rect 6972 58212 7028 58942
rect 7084 58212 7140 60060
rect 7308 59892 7364 59902
rect 7196 59108 7252 59118
rect 7196 59014 7252 59052
rect 7308 58772 7364 59836
rect 7532 59778 7588 60844
rect 7756 60004 7812 60014
rect 7756 59910 7812 59948
rect 7532 59726 7534 59778
rect 7586 59726 7588 59778
rect 7532 58994 7588 59726
rect 7644 59780 7700 59790
rect 7644 59778 7812 59780
rect 7644 59726 7646 59778
rect 7698 59726 7812 59778
rect 7644 59724 7812 59726
rect 7644 59714 7700 59724
rect 7532 58942 7534 58994
rect 7586 58942 7588 58994
rect 7532 58930 7588 58942
rect 7644 59106 7700 59118
rect 7644 59054 7646 59106
rect 7698 59054 7700 59106
rect 7644 58996 7700 59054
rect 7644 58930 7700 58940
rect 7308 58716 7700 58772
rect 7308 58548 7364 58558
rect 7308 58546 7476 58548
rect 7308 58494 7310 58546
rect 7362 58494 7476 58546
rect 7308 58492 7476 58494
rect 7308 58482 7364 58492
rect 7196 58436 7252 58446
rect 7196 58342 7252 58380
rect 7308 58324 7364 58334
rect 7308 58230 7364 58268
rect 7084 58156 7252 58212
rect 6972 58118 7028 58156
rect 6748 57932 7140 57988
rect 7084 57762 7140 57932
rect 7084 57710 7086 57762
rect 7138 57710 7140 57762
rect 7084 57698 7140 57710
rect 6972 57652 7028 57662
rect 6860 57596 6972 57652
rect 6860 57538 6916 57596
rect 6972 57586 7028 57596
rect 6860 57486 6862 57538
rect 6914 57486 6916 57538
rect 6860 57474 6916 57486
rect 6524 57428 6580 57438
rect 6524 57426 6692 57428
rect 6524 57374 6526 57426
rect 6578 57374 6692 57426
rect 6524 57372 6692 57374
rect 6524 57362 6580 57372
rect 6636 56868 6692 57372
rect 6860 56868 6916 56878
rect 6636 56866 6916 56868
rect 6636 56814 6862 56866
rect 6914 56814 6916 56866
rect 6636 56812 6916 56814
rect 6860 56802 6916 56812
rect 6636 56644 6692 56654
rect 6524 56642 6692 56644
rect 6524 56590 6638 56642
rect 6690 56590 6692 56642
rect 6524 56588 6692 56590
rect 6524 55410 6580 56588
rect 6636 56578 6692 56588
rect 6524 55358 6526 55410
rect 6578 55358 6580 55410
rect 6524 55346 6580 55358
rect 6860 54628 6916 54638
rect 6860 54534 6916 54572
rect 6636 53172 6692 53182
rect 6636 52946 6692 53116
rect 6636 52894 6638 52946
rect 6690 52894 6692 52946
rect 6636 50820 6692 52894
rect 6860 52836 6916 52846
rect 6860 52742 6916 52780
rect 7196 52500 7252 58156
rect 7308 53732 7364 53742
rect 7308 53172 7364 53676
rect 7308 53078 7364 53116
rect 7308 52500 7364 52510
rect 7196 52444 7308 52500
rect 7308 52434 7364 52444
rect 6636 50818 7364 50820
rect 6636 50766 6638 50818
rect 6690 50766 7364 50818
rect 6636 50764 7364 50766
rect 6636 50754 6692 50764
rect 7308 50706 7364 50764
rect 7308 50654 7310 50706
rect 7362 50654 7364 50706
rect 7308 50642 7364 50654
rect 6860 50482 6916 50494
rect 6860 50430 6862 50482
rect 6914 50430 6916 50482
rect 6748 48802 6804 48814
rect 6748 48750 6750 48802
rect 6802 48750 6804 48802
rect 6748 48354 6804 48750
rect 6860 48692 6916 50430
rect 7420 50428 7476 58492
rect 7532 58322 7588 58334
rect 7532 58270 7534 58322
rect 7586 58270 7588 58322
rect 7532 57874 7588 58270
rect 7532 57822 7534 57874
rect 7586 57822 7588 57874
rect 7532 57652 7588 57822
rect 7532 57586 7588 57596
rect 7644 57428 7700 58716
rect 7532 57372 7700 57428
rect 7532 52612 7588 57372
rect 7644 52724 7700 52734
rect 7644 52630 7700 52668
rect 7532 52546 7588 52556
rect 7756 52500 7812 59724
rect 7868 58436 7924 62132
rect 7980 61684 8036 61694
rect 7980 61010 8036 61628
rect 7980 60958 7982 61010
rect 8034 60958 8036 61010
rect 7980 58658 8036 60958
rect 8092 61346 8148 61358
rect 8092 61294 8094 61346
rect 8146 61294 8148 61346
rect 8092 60788 8148 61294
rect 8092 60722 8148 60732
rect 8204 60228 8260 62132
rect 7980 58606 7982 58658
rect 8034 58606 8036 58658
rect 7980 58594 8036 58606
rect 8092 60172 8260 60228
rect 7868 58380 8036 58436
rect 7868 58212 7924 58222
rect 7868 58118 7924 58156
rect 7980 53844 8036 58380
rect 7644 52444 7812 52500
rect 7868 53788 8036 53844
rect 7420 50372 7588 50428
rect 7084 48916 7140 48926
rect 7420 48916 7476 48926
rect 7084 48914 7476 48916
rect 7084 48862 7086 48914
rect 7138 48862 7422 48914
rect 7474 48862 7476 48914
rect 7084 48860 7476 48862
rect 7084 48850 7140 48860
rect 7420 48850 7476 48860
rect 6860 48626 6916 48636
rect 6748 48302 6750 48354
rect 6802 48302 6804 48354
rect 6748 48290 6804 48302
rect 6860 47348 6916 47358
rect 6860 47346 7476 47348
rect 6860 47294 6862 47346
rect 6914 47294 7476 47346
rect 6860 47292 7476 47294
rect 6860 47282 6916 47292
rect 7420 46898 7476 47292
rect 7420 46846 7422 46898
rect 7474 46846 7476 46898
rect 7420 46834 7476 46846
rect 6636 44210 6692 44222
rect 6636 44158 6638 44210
rect 6690 44158 6692 44210
rect 6636 42980 6692 44158
rect 6972 44100 7028 44110
rect 6972 44098 7364 44100
rect 6972 44046 6974 44098
rect 7026 44046 7364 44098
rect 6972 44044 7364 44046
rect 6972 44034 7028 44044
rect 6860 43428 6916 43438
rect 6636 42914 6692 42924
rect 6748 43426 6916 43428
rect 6748 43374 6862 43426
rect 6914 43374 6916 43426
rect 6748 43372 6916 43374
rect 6636 42756 6692 42766
rect 6636 42662 6692 42700
rect 6636 41748 6692 41758
rect 6524 41746 6692 41748
rect 6524 41694 6638 41746
rect 6690 41694 6692 41746
rect 6524 41692 6692 41694
rect 6524 41186 6580 41692
rect 6636 41682 6692 41692
rect 6524 41134 6526 41186
rect 6578 41134 6580 41186
rect 6524 41122 6580 41134
rect 6748 41074 6804 43372
rect 6860 43362 6916 43372
rect 7308 42866 7364 44044
rect 7308 42814 7310 42866
rect 7362 42814 7364 42866
rect 7308 42802 7364 42814
rect 7308 41972 7364 41982
rect 7196 41860 7252 41870
rect 7196 41766 7252 41804
rect 6972 41746 7028 41758
rect 6972 41694 6974 41746
rect 7026 41694 7028 41746
rect 6972 41636 7028 41694
rect 6972 41570 7028 41580
rect 7196 41300 7252 41310
rect 7308 41300 7364 41916
rect 6748 41022 6750 41074
rect 6802 41022 6804 41074
rect 6748 41010 6804 41022
rect 6860 41298 7364 41300
rect 6860 41246 7198 41298
rect 7250 41246 7364 41298
rect 6860 41244 7364 41246
rect 7420 41748 7476 41758
rect 6412 40908 6692 40964
rect 6524 40402 6580 40414
rect 6524 40350 6526 40402
rect 6578 40350 6580 40402
rect 6524 40292 6580 40350
rect 6524 40226 6580 40236
rect 6188 40012 6580 40068
rect 6188 39732 6244 39742
rect 6188 39730 6468 39732
rect 6188 39678 6190 39730
rect 6242 39678 6468 39730
rect 6188 39676 6468 39678
rect 6188 39666 6244 39676
rect 6300 39508 6356 39518
rect 6188 39452 6300 39508
rect 6076 39396 6132 39406
rect 6076 39302 6132 39340
rect 6188 39394 6244 39452
rect 6300 39442 6356 39452
rect 6188 39342 6190 39394
rect 6242 39342 6244 39394
rect 6188 39330 6244 39342
rect 5964 38894 5966 38946
rect 6018 38894 6020 38946
rect 5964 38882 6020 38894
rect 6300 38946 6356 38958
rect 6300 38894 6302 38946
rect 6354 38894 6356 38946
rect 5852 38836 5908 38846
rect 5740 38834 5908 38836
rect 5740 38782 5854 38834
rect 5906 38782 5908 38834
rect 5740 38780 5908 38782
rect 5852 38770 5908 38780
rect 5628 38724 5684 38734
rect 5628 38612 5796 38668
rect 5404 38098 5460 38108
rect 5740 38162 5796 38612
rect 5740 38110 5742 38162
rect 5794 38110 5796 38162
rect 5740 38098 5796 38110
rect 5964 38612 6020 38622
rect 5292 30830 5294 30882
rect 5346 30830 5348 30882
rect 5292 30818 5348 30830
rect 5404 37436 5796 37492
rect 3948 29474 4004 29484
rect 4620 30380 4900 30436
rect 4620 29428 4676 30380
rect 4732 30212 4788 30222
rect 4732 30118 4788 30156
rect 5292 30212 5348 30222
rect 4732 29652 4788 29662
rect 4956 29652 5012 29662
rect 4788 29650 5012 29652
rect 4788 29598 4958 29650
rect 5010 29598 5012 29650
rect 4788 29596 5012 29598
rect 4732 29586 4788 29596
rect 4956 29586 5012 29596
rect 3724 29260 4340 29316
rect 3612 29148 4004 29204
rect 3388 28644 3444 28654
rect 3836 28644 3892 28654
rect 3388 28642 3892 28644
rect 3388 28590 3390 28642
rect 3442 28590 3838 28642
rect 3890 28590 3892 28642
rect 3388 28588 3892 28590
rect 3388 28578 3444 28588
rect 3836 28578 3892 28588
rect 3052 28478 3054 28530
rect 3106 28478 3108 28530
rect 3052 28466 3108 28478
rect 1820 27076 1876 27086
rect 1708 27074 1876 27076
rect 1708 27022 1822 27074
rect 1874 27022 1876 27074
rect 1708 27020 1876 27022
rect 1820 27010 1876 27020
rect 2604 26962 2660 26974
rect 2604 26910 2606 26962
rect 2658 26910 2660 26962
rect 2604 25396 2660 26910
rect 3836 26068 3892 26078
rect 2604 25330 2660 25340
rect 3612 26012 3836 26068
rect 3276 24836 3332 24846
rect 2492 24834 3332 24836
rect 2492 24782 3278 24834
rect 3330 24782 3332 24834
rect 2492 24780 3332 24782
rect 1820 23154 1876 23166
rect 1820 23102 1822 23154
rect 1874 23102 1876 23154
rect 1820 22372 1876 23102
rect 2492 22482 2548 24780
rect 3276 24770 3332 24780
rect 3612 24834 3668 26012
rect 3836 26002 3892 26012
rect 3948 25508 4004 29148
rect 4284 28756 4340 29260
rect 4620 29314 4676 29372
rect 4620 29262 4622 29314
rect 4674 29262 4676 29314
rect 4620 29250 4676 29262
rect 4844 29316 4900 29326
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4396 28756 4452 28766
rect 4284 28754 4452 28756
rect 4284 28702 4398 28754
rect 4450 28702 4452 28754
rect 4284 28700 4452 28702
rect 4172 28644 4228 28654
rect 4172 28550 4228 28588
rect 4284 27300 4340 28700
rect 4396 28690 4452 28700
rect 4844 28754 4900 29260
rect 4844 28702 4846 28754
rect 4898 28702 4900 28754
rect 4620 28644 4676 28654
rect 4620 27746 4676 28588
rect 4844 28644 4900 28702
rect 5292 29202 5348 30156
rect 5292 29150 5294 29202
rect 5346 29150 5348 29202
rect 5292 28756 5348 29150
rect 5292 28690 5348 28700
rect 4844 28578 4900 28588
rect 5404 28532 5460 37436
rect 5516 37266 5572 37278
rect 5516 37214 5518 37266
rect 5570 37214 5572 37266
rect 5516 36708 5572 37214
rect 5628 37268 5684 37278
rect 5628 37174 5684 37212
rect 5740 37266 5796 37436
rect 5740 37214 5742 37266
rect 5794 37214 5796 37266
rect 5740 37202 5796 37214
rect 5964 37266 6020 38556
rect 5964 37214 5966 37266
rect 6018 37214 6020 37266
rect 5964 37202 6020 37214
rect 6076 36708 6132 36718
rect 5516 36652 6020 36708
rect 5964 36594 6020 36652
rect 5964 36542 5966 36594
rect 6018 36542 6020 36594
rect 5964 36530 6020 36542
rect 5852 36484 5908 36494
rect 5628 36372 5684 36382
rect 5628 36278 5684 36316
rect 5852 35924 5908 36428
rect 6076 36482 6132 36652
rect 6076 36430 6078 36482
rect 6130 36430 6132 36482
rect 6076 36418 6132 36430
rect 6188 36258 6244 36270
rect 6188 36206 6190 36258
rect 6242 36206 6244 36258
rect 5852 35868 6020 35924
rect 5516 35700 5572 35710
rect 5516 35364 5572 35644
rect 5516 35298 5572 35308
rect 5852 34914 5908 34926
rect 5852 34862 5854 34914
rect 5906 34862 5908 34914
rect 5852 34020 5908 34862
rect 5964 34916 6020 35868
rect 6188 35700 6244 36206
rect 6188 34916 6244 35644
rect 6300 35252 6356 38894
rect 6412 38834 6468 39676
rect 6412 38782 6414 38834
rect 6466 38782 6468 38834
rect 6412 38770 6468 38782
rect 6412 37042 6468 37054
rect 6412 36990 6414 37042
rect 6466 36990 6468 37042
rect 6412 35812 6468 36990
rect 6412 35746 6468 35756
rect 6524 35588 6580 40012
rect 6636 35924 6692 40908
rect 6748 39732 6804 39742
rect 6860 39732 6916 41244
rect 7196 41234 7252 41244
rect 6804 39676 6916 39732
rect 6972 40852 7028 40862
rect 6972 40626 7028 40796
rect 6972 40574 6974 40626
rect 7026 40574 7028 40626
rect 6972 40404 7028 40574
rect 6748 39638 6804 39676
rect 6860 38948 6916 38958
rect 6860 38854 6916 38892
rect 6972 38668 7028 40348
rect 7196 39732 7252 39742
rect 7420 39732 7476 41692
rect 7196 39730 7476 39732
rect 7196 39678 7198 39730
rect 7250 39678 7476 39730
rect 7196 39676 7476 39678
rect 7196 39508 7252 39676
rect 7196 39442 7252 39452
rect 6972 38612 7252 38668
rect 6748 37156 6804 37194
rect 6748 37090 6804 37100
rect 6748 36932 6804 36942
rect 6748 36594 6804 36876
rect 6748 36542 6750 36594
rect 6802 36542 6804 36594
rect 6748 36484 6804 36542
rect 6748 36418 6804 36428
rect 7196 36258 7252 38612
rect 7420 38164 7476 38174
rect 7420 38070 7476 38108
rect 7532 36596 7588 50372
rect 7644 49476 7700 52444
rect 7868 50428 7924 53788
rect 7980 53620 8036 53630
rect 7980 53526 8036 53564
rect 7980 53172 8036 53182
rect 7980 52946 8036 53116
rect 7980 52894 7982 52946
rect 8034 52894 8036 52946
rect 7980 52882 8036 52894
rect 7644 49410 7700 49420
rect 7756 50372 7924 50428
rect 7756 49252 7812 50372
rect 7980 49588 8036 49598
rect 7644 49196 7812 49252
rect 7868 49586 8036 49588
rect 7868 49534 7982 49586
rect 8034 49534 8036 49586
rect 7868 49532 8036 49534
rect 7644 46452 7700 49196
rect 7756 49028 7812 49038
rect 7868 49028 7924 49532
rect 7980 49522 8036 49532
rect 7980 49252 8036 49262
rect 7980 49138 8036 49196
rect 7980 49086 7982 49138
rect 8034 49086 8036 49138
rect 7980 49074 8036 49086
rect 7756 49026 7924 49028
rect 7756 48974 7758 49026
rect 7810 48974 7924 49026
rect 7756 48972 7924 48974
rect 7756 47236 7812 48972
rect 7756 47170 7812 47180
rect 7756 46676 7812 46686
rect 7756 46674 8036 46676
rect 7756 46622 7758 46674
rect 7810 46622 8036 46674
rect 7756 46620 8036 46622
rect 7756 46610 7812 46620
rect 7644 46396 7924 46452
rect 7644 44994 7700 45006
rect 7644 44942 7646 44994
rect 7698 44942 7700 44994
rect 7644 44884 7700 44942
rect 7644 41858 7700 44828
rect 7644 41806 7646 41858
rect 7698 41806 7700 41858
rect 7644 41636 7700 41806
rect 7644 41570 7700 41580
rect 7532 36530 7588 36540
rect 7196 36206 7198 36258
rect 7250 36206 7252 36258
rect 6636 35868 6804 35924
rect 6300 35186 6356 35196
rect 6412 35532 6580 35588
rect 6636 35700 6692 35710
rect 6636 35586 6692 35644
rect 6636 35534 6638 35586
rect 6690 35534 6692 35586
rect 6300 34916 6356 34926
rect 6188 34914 6356 34916
rect 6188 34862 6302 34914
rect 6354 34862 6356 34914
rect 6188 34860 6356 34862
rect 5964 34822 6020 34860
rect 6300 34850 6356 34860
rect 6076 34690 6132 34702
rect 6076 34638 6078 34690
rect 6130 34638 6132 34690
rect 6076 34130 6132 34638
rect 6188 34690 6244 34702
rect 6188 34638 6190 34690
rect 6242 34638 6244 34690
rect 6188 34356 6244 34638
rect 6412 34692 6468 35532
rect 6636 35522 6692 35534
rect 6524 35252 6580 35262
rect 6748 35252 6804 35868
rect 6972 35700 7028 35710
rect 6580 35196 6692 35252
rect 6524 35186 6580 35196
rect 6412 34636 6580 34692
rect 6188 34300 6468 34356
rect 6076 34078 6078 34130
rect 6130 34078 6132 34130
rect 6076 34066 6132 34078
rect 6188 34132 6244 34142
rect 6188 34038 6244 34076
rect 6300 34130 6356 34142
rect 6300 34078 6302 34130
rect 6354 34078 6356 34130
rect 5852 33460 5908 33964
rect 5964 33460 6020 33470
rect 5852 33458 6020 33460
rect 5852 33406 5966 33458
rect 6018 33406 6020 33458
rect 5852 33404 6020 33406
rect 5964 33394 6020 33404
rect 6188 33348 6244 33358
rect 6188 33254 6244 33292
rect 5740 31780 5796 31790
rect 5740 31218 5796 31724
rect 5740 31166 5742 31218
rect 5794 31166 5796 31218
rect 5740 31154 5796 31166
rect 5516 29428 5572 29438
rect 5516 29334 5572 29372
rect 6300 28868 6356 34078
rect 6412 32452 6468 34300
rect 6524 34130 6580 34636
rect 6524 34078 6526 34130
rect 6578 34078 6580 34130
rect 6524 34066 6580 34078
rect 6524 33908 6580 33918
rect 6524 33570 6580 33852
rect 6524 33518 6526 33570
rect 6578 33518 6580 33570
rect 6524 33506 6580 33518
rect 6412 32386 6468 32396
rect 6188 28812 6356 28868
rect 4620 27694 4622 27746
rect 4674 27694 4676 27746
rect 4620 27636 4676 27694
rect 5292 28476 5460 28532
rect 5740 28532 5796 28542
rect 6076 28532 6132 28542
rect 4620 27580 4900 27636
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 4284 27244 4788 27300
rect 4732 27186 4788 27244
rect 4732 27134 4734 27186
rect 4786 27134 4788 27186
rect 4732 27122 4788 27134
rect 4844 26908 4900 27580
rect 4508 26852 4900 26908
rect 4508 26180 4564 26852
rect 4508 26086 4564 26124
rect 5180 26180 5236 26190
rect 4844 26068 4900 26078
rect 4844 25974 4900 26012
rect 5180 26066 5236 26124
rect 5180 26014 5182 26066
rect 5234 26014 5236 26066
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 3948 25442 4004 25452
rect 3724 25396 3780 25406
rect 3724 25302 3780 25340
rect 4060 25394 4116 25406
rect 4060 25342 4062 25394
rect 4114 25342 4116 25394
rect 3612 24782 3614 24834
rect 3666 24782 3668 24834
rect 3612 24770 3668 24782
rect 3948 24834 4004 24846
rect 3948 24782 3950 24834
rect 4002 24782 4004 24834
rect 2604 23940 2660 23950
rect 2604 23266 2660 23884
rect 3948 23940 4004 24782
rect 4060 24164 4116 25342
rect 4284 25284 4340 25294
rect 4284 24834 4340 25228
rect 4284 24782 4286 24834
rect 4338 24782 4340 24834
rect 4284 24770 4340 24782
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4060 24098 4116 24108
rect 3948 23874 4004 23884
rect 5180 23940 5236 26014
rect 5068 23716 5124 23726
rect 5180 23716 5236 23884
rect 5068 23714 5236 23716
rect 5068 23662 5070 23714
rect 5122 23662 5236 23714
rect 5068 23660 5236 23662
rect 5068 23650 5124 23660
rect 2604 23214 2606 23266
rect 2658 23214 2660 23266
rect 2604 23202 2660 23214
rect 4732 23044 4788 23054
rect 4732 22950 4788 22988
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 5068 22596 5124 22606
rect 2492 22430 2494 22482
rect 2546 22430 2548 22482
rect 2492 22418 2548 22430
rect 4620 22484 4676 22494
rect 1820 22278 1876 22316
rect 4620 21924 4676 22428
rect 5068 22482 5124 22540
rect 5068 22430 5070 22482
rect 5122 22430 5124 22482
rect 5068 22418 5124 22430
rect 4620 21868 4900 21924
rect 4732 21700 4788 21710
rect 4172 21698 4788 21700
rect 4172 21646 4734 21698
rect 4786 21646 4788 21698
rect 4172 21644 4788 21646
rect 4172 20802 4228 21644
rect 4732 21634 4788 21644
rect 4396 21476 4452 21486
rect 4396 21382 4452 21420
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 4172 20750 4174 20802
rect 4226 20750 4228 20802
rect 4172 20738 4228 20750
rect 3836 20580 3892 20590
rect 3500 20578 3892 20580
rect 3500 20526 3838 20578
rect 3890 20526 3892 20578
rect 3500 20524 3892 20526
rect 3500 20188 3556 20524
rect 3836 20514 3892 20524
rect 3276 20132 3556 20188
rect 3276 20130 3332 20132
rect 3276 20078 3278 20130
rect 3330 20078 3332 20130
rect 3276 20066 3332 20078
rect 2604 20018 2660 20030
rect 2604 19966 2606 20018
rect 2658 19966 2660 20018
rect 2268 18452 2324 18462
rect 2604 18452 2660 19966
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4172 19460 4228 19470
rect 3836 19012 3892 19022
rect 2268 18450 2660 18452
rect 2268 18398 2270 18450
rect 2322 18398 2660 18450
rect 2268 18396 2660 18398
rect 2268 18386 2324 18396
rect 2604 18340 2660 18396
rect 3612 19010 3892 19012
rect 3612 18958 3838 19010
rect 3890 18958 3892 19010
rect 3612 18956 3892 18958
rect 2604 18274 2660 18284
rect 2940 18340 2996 18350
rect 2940 18338 3332 18340
rect 2940 18286 2942 18338
rect 2994 18286 3332 18338
rect 2940 18284 3332 18286
rect 2940 18274 2996 18284
rect 3276 17554 3332 18284
rect 3612 17666 3668 18956
rect 3836 18946 3892 18956
rect 3612 17614 3614 17666
rect 3666 17614 3668 17666
rect 3612 17602 3668 17614
rect 3276 17502 3278 17554
rect 3330 17502 3332 17554
rect 3276 17490 3332 17502
rect 4172 15148 4228 19404
rect 4396 19348 4452 19358
rect 4844 19348 4900 21868
rect 5068 21362 5124 21374
rect 5068 21310 5070 21362
rect 5122 21310 5124 21362
rect 5068 20804 5124 21310
rect 5068 20710 5124 20748
rect 4396 19346 4900 19348
rect 4396 19294 4398 19346
rect 4450 19294 4900 19346
rect 4396 19292 4900 19294
rect 4956 19460 5012 19470
rect 5180 19460 5236 23660
rect 5292 23380 5348 28476
rect 5516 27298 5572 27310
rect 5516 27246 5518 27298
rect 5570 27246 5572 27298
rect 5516 26908 5572 27246
rect 5740 27186 5796 28476
rect 5740 27134 5742 27186
rect 5794 27134 5796 27186
rect 5740 27122 5796 27134
rect 5852 28476 6076 28532
rect 5404 26852 5572 26908
rect 5404 26290 5460 26852
rect 5404 26238 5406 26290
rect 5458 26238 5460 26290
rect 5404 26226 5460 26238
rect 5628 25284 5684 25294
rect 5628 25190 5684 25228
rect 5628 24164 5684 24174
rect 5628 24070 5684 24108
rect 5852 23604 5908 28476
rect 6076 28466 6132 28476
rect 6188 27972 6244 28812
rect 6524 28756 6580 28766
rect 6636 28756 6692 35196
rect 6748 35186 6804 35196
rect 6860 35698 7028 35700
rect 6860 35646 6974 35698
rect 7026 35646 7028 35698
rect 6860 35644 7028 35646
rect 6748 34914 6804 34926
rect 6748 34862 6750 34914
rect 6802 34862 6804 34914
rect 6748 34244 6804 34862
rect 6748 34178 6804 34188
rect 6860 33908 6916 35644
rect 6972 35634 7028 35644
rect 7196 35700 7252 36206
rect 7308 35812 7364 35822
rect 7308 35810 7588 35812
rect 7308 35758 7310 35810
rect 7362 35758 7588 35810
rect 7308 35756 7588 35758
rect 7308 35746 7364 35756
rect 7196 35634 7252 35644
rect 7084 35364 7140 35374
rect 6972 34356 7028 34366
rect 6972 34262 7028 34300
rect 6860 33842 6916 33852
rect 6972 33348 7028 33358
rect 6748 32452 6804 32462
rect 6748 32358 6804 32396
rect 6524 28754 6692 28756
rect 6524 28702 6526 28754
rect 6578 28702 6692 28754
rect 6524 28700 6692 28702
rect 6524 28690 6580 28700
rect 6300 28644 6356 28654
rect 6300 28550 6356 28588
rect 6748 28642 6804 28654
rect 6748 28590 6750 28642
rect 6802 28590 6804 28642
rect 6188 27906 6244 27916
rect 6412 28530 6468 28542
rect 6412 28478 6414 28530
rect 6466 28478 6468 28530
rect 6076 27748 6132 27758
rect 6412 27748 6468 28478
rect 6636 28532 6692 28542
rect 6636 28438 6692 28476
rect 6748 28196 6804 28590
rect 6076 27746 6468 27748
rect 6076 27694 6078 27746
rect 6130 27694 6468 27746
rect 6076 27692 6468 27694
rect 6524 28140 6804 28196
rect 6076 27298 6132 27692
rect 6076 27246 6078 27298
rect 6130 27246 6132 27298
rect 6076 27234 6132 27246
rect 6300 27188 6356 27198
rect 6524 27188 6580 28140
rect 6300 27186 6580 27188
rect 6300 27134 6302 27186
rect 6354 27134 6580 27186
rect 6300 27132 6580 27134
rect 6636 27972 6692 27982
rect 6300 26908 6356 27132
rect 6188 26852 6356 26908
rect 6524 26964 6580 26974
rect 6188 25618 6244 26852
rect 6524 25620 6580 26908
rect 6636 25844 6692 27916
rect 6972 27860 7028 33292
rect 7084 32788 7140 35308
rect 7196 35252 7252 35262
rect 7196 34132 7252 35196
rect 7532 35026 7588 35756
rect 7532 34974 7534 35026
rect 7586 34974 7588 35026
rect 7532 34962 7588 34974
rect 7420 34916 7476 34926
rect 7420 34354 7476 34860
rect 7420 34302 7422 34354
rect 7474 34302 7476 34354
rect 7420 34290 7476 34302
rect 7196 34066 7252 34076
rect 7308 34244 7364 34254
rect 7308 34020 7364 34188
rect 7756 34132 7812 34142
rect 7756 34038 7812 34076
rect 7420 34020 7476 34030
rect 7308 33964 7420 34020
rect 7420 33458 7476 33964
rect 7420 33406 7422 33458
rect 7474 33406 7476 33458
rect 7420 33124 7476 33406
rect 7084 32732 7364 32788
rect 7308 32676 7364 32732
rect 7308 32562 7364 32620
rect 7308 32510 7310 32562
rect 7362 32510 7364 32562
rect 7308 32498 7364 32510
rect 7084 32452 7140 32462
rect 7084 32358 7140 32396
rect 7308 31780 7364 31790
rect 7420 31780 7476 33068
rect 7756 32676 7812 32686
rect 7364 31724 7476 31780
rect 7644 32338 7700 32350
rect 7644 32286 7646 32338
rect 7698 32286 7700 32338
rect 7308 31686 7364 31724
rect 7644 31106 7700 32286
rect 7644 31054 7646 31106
rect 7698 31054 7700 31106
rect 7644 31042 7700 31054
rect 7756 31220 7812 32620
rect 7308 30212 7364 30222
rect 6972 26964 7028 27804
rect 6972 26898 7028 26908
rect 7084 29314 7140 29326
rect 7084 29262 7086 29314
rect 7138 29262 7140 29314
rect 7084 28644 7140 29262
rect 6636 25788 6804 25844
rect 6636 25620 6692 25630
rect 6188 25566 6190 25618
rect 6242 25566 6244 25618
rect 6188 25554 6244 25566
rect 6300 25618 6692 25620
rect 6300 25566 6638 25618
rect 6690 25566 6692 25618
rect 6300 25564 6692 25566
rect 5964 25506 6020 25518
rect 5964 25454 5966 25506
rect 6018 25454 6020 25506
rect 5964 25396 6020 25454
rect 6300 25396 6356 25564
rect 6636 25554 6692 25564
rect 6748 25396 6804 25788
rect 5964 25340 6356 25396
rect 6412 25340 6804 25396
rect 5964 23940 6020 23950
rect 5964 23846 6020 23884
rect 6188 23940 6244 23950
rect 6188 23846 6244 23884
rect 5852 23548 6020 23604
rect 5516 23380 5572 23390
rect 5292 23378 5572 23380
rect 5292 23326 5518 23378
rect 5570 23326 5572 23378
rect 5292 23324 5572 23326
rect 5516 23314 5572 23324
rect 5852 23380 5908 23390
rect 5292 23154 5348 23166
rect 5292 23102 5294 23154
rect 5346 23102 5348 23154
rect 5292 23044 5348 23102
rect 5404 23156 5460 23166
rect 5404 23062 5460 23100
rect 5628 23154 5684 23166
rect 5628 23102 5630 23154
rect 5682 23102 5684 23154
rect 5292 21586 5348 22988
rect 5628 22484 5684 23102
rect 5852 23154 5908 23324
rect 5852 23102 5854 23154
rect 5906 23102 5908 23154
rect 5852 23090 5908 23102
rect 5964 23156 6020 23548
rect 6300 23156 6356 23166
rect 5964 23100 6300 23156
rect 5628 22418 5684 22428
rect 5852 22596 5908 22606
rect 5292 21534 5294 21586
rect 5346 21534 5348 21586
rect 5292 21522 5348 21534
rect 5740 22258 5796 22270
rect 5740 22206 5742 22258
rect 5794 22206 5796 22258
rect 5740 20916 5796 22206
rect 5852 21588 5908 22540
rect 5964 22370 6020 23100
rect 6300 23062 6356 23100
rect 6300 22484 6356 22494
rect 6412 22484 6468 25340
rect 6748 23604 6804 23614
rect 7084 23604 7140 28588
rect 7308 28754 7364 30156
rect 7308 28702 7310 28754
rect 7362 28702 7364 28754
rect 7308 28644 7364 28702
rect 7308 28578 7364 28588
rect 7308 23604 7364 23614
rect 7084 23548 7308 23604
rect 6748 23380 6804 23548
rect 6748 23286 6804 23324
rect 6300 22482 6468 22484
rect 6300 22430 6302 22482
rect 6354 22430 6468 22482
rect 6300 22428 6468 22430
rect 6860 23156 6916 23166
rect 6860 22482 6916 23100
rect 6860 22430 6862 22482
rect 6914 22430 6916 22482
rect 6300 22418 6356 22428
rect 6860 22418 6916 22430
rect 7308 22482 7364 23548
rect 7308 22430 7310 22482
rect 7362 22430 7364 22482
rect 5964 22318 5966 22370
rect 6018 22318 6020 22370
rect 5964 22306 6020 22318
rect 6188 22148 6244 22158
rect 6076 22146 6244 22148
rect 6076 22094 6190 22146
rect 6242 22094 6244 22146
rect 6076 22092 6244 22094
rect 5964 21588 6020 21598
rect 5852 21586 6020 21588
rect 5852 21534 5966 21586
rect 6018 21534 6020 21586
rect 5852 21532 6020 21534
rect 5852 21476 5908 21532
rect 5964 21522 6020 21532
rect 5852 21410 5908 21420
rect 5404 20914 5796 20916
rect 5404 20862 5742 20914
rect 5794 20862 5796 20914
rect 5404 20860 5796 20862
rect 5404 19906 5460 20860
rect 5740 20850 5796 20860
rect 5964 20804 6020 20814
rect 5964 20710 6020 20748
rect 5404 19854 5406 19906
rect 5458 19854 5460 19906
rect 5404 19842 5460 19854
rect 5964 19906 6020 19918
rect 5964 19854 5966 19906
rect 6018 19854 6020 19906
rect 5964 19460 6020 19854
rect 5012 19404 5236 19460
rect 5516 19404 6020 19460
rect 4396 19282 4452 19292
rect 4844 19012 4900 19022
rect 4956 19012 5012 19404
rect 4844 19010 5012 19012
rect 4844 18958 4846 19010
rect 4898 18958 5012 19010
rect 4844 18956 5012 18958
rect 4844 18946 4900 18956
rect 4956 18564 5012 18956
rect 5068 18564 5124 18574
rect 4956 18508 5068 18564
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 4956 17780 5012 18508
rect 5068 18498 5124 18508
rect 5068 18340 5124 18350
rect 5516 18340 5572 19404
rect 6076 19348 6132 22092
rect 6188 22082 6244 22092
rect 6300 22148 6356 22158
rect 6300 22054 6356 22092
rect 7308 22148 7364 22430
rect 7308 22082 7364 22092
rect 6748 21476 6804 21486
rect 6748 21474 7028 21476
rect 6748 21422 6750 21474
rect 6802 21422 7028 21474
rect 6748 21420 7028 21422
rect 6748 21410 6804 21420
rect 6300 20692 6356 20702
rect 6636 20692 6692 20702
rect 6300 20690 6692 20692
rect 6300 20638 6302 20690
rect 6354 20638 6638 20690
rect 6690 20638 6692 20690
rect 6300 20636 6692 20638
rect 6300 20626 6356 20636
rect 6636 20626 6692 20636
rect 6972 20690 7028 21420
rect 7420 21140 7476 21150
rect 6972 20638 6974 20690
rect 7026 20638 7028 20690
rect 6972 20626 7028 20638
rect 7308 21084 7420 21140
rect 6300 20244 6356 20254
rect 5068 18338 5348 18340
rect 5068 18286 5070 18338
rect 5122 18286 5348 18338
rect 5068 18284 5348 18286
rect 5068 18274 5124 18284
rect 5292 18226 5348 18284
rect 5292 18174 5294 18226
rect 5346 18174 5348 18226
rect 5292 18162 5348 18174
rect 5068 17780 5124 17790
rect 4956 17778 5124 17780
rect 4956 17726 5070 17778
rect 5122 17726 5124 17778
rect 4956 17724 5124 17726
rect 5068 17714 5124 17724
rect 5516 17108 5572 18284
rect 5628 19292 6132 19348
rect 6188 20188 6300 20244
rect 5628 18226 5684 19292
rect 6188 19236 6244 20188
rect 6300 20178 6356 20188
rect 5628 18174 5630 18226
rect 5682 18174 5684 18226
rect 5628 17778 5684 18174
rect 5852 19180 6244 19236
rect 5852 18564 5908 19180
rect 5852 17890 5908 18508
rect 5852 17838 5854 17890
rect 5906 17838 5908 17890
rect 5852 17826 5908 17838
rect 5628 17726 5630 17778
rect 5682 17726 5684 17778
rect 5628 17714 5684 17726
rect 6188 17668 6244 17678
rect 6748 17668 6804 17678
rect 6188 17666 6804 17668
rect 6188 17614 6190 17666
rect 6242 17614 6750 17666
rect 6802 17614 6804 17666
rect 6188 17612 6804 17614
rect 6188 17602 6244 17612
rect 6748 17602 6804 17612
rect 6524 17444 6580 17454
rect 5404 16884 5460 16894
rect 5516 16884 5572 17052
rect 6076 17442 6580 17444
rect 6076 17390 6526 17442
rect 6578 17390 6580 17442
rect 6076 17388 6580 17390
rect 6076 16994 6132 17388
rect 6524 17378 6580 17388
rect 6076 16942 6078 16994
rect 6130 16942 6132 16994
rect 6076 16930 6132 16942
rect 5404 16882 5572 16884
rect 5404 16830 5406 16882
rect 5458 16830 5572 16882
rect 5404 16828 5572 16830
rect 5404 16818 5460 16828
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 7084 15988 7140 15998
rect 6860 15316 6916 15326
rect 6860 15148 6916 15260
rect 7084 15314 7140 15932
rect 7084 15262 7086 15314
rect 7138 15262 7140 15314
rect 7084 15250 7140 15262
rect 4172 15092 4340 15148
rect 4284 10498 4340 15092
rect 6524 15090 6580 15102
rect 6860 15092 7252 15148
rect 6524 15038 6526 15090
rect 6578 15038 6580 15090
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 6300 14532 6356 14542
rect 6524 14532 6580 15038
rect 6300 14530 6580 14532
rect 6300 14478 6302 14530
rect 6354 14478 6580 14530
rect 6300 14476 6580 14478
rect 6300 14466 6356 14476
rect 5964 14308 6020 14318
rect 5404 14306 6020 14308
rect 5404 14254 5966 14306
rect 6018 14254 6020 14306
rect 5404 14252 6020 14254
rect 5404 13858 5460 14252
rect 5964 14242 6020 14252
rect 5404 13806 5406 13858
rect 5458 13806 5460 13858
rect 5404 13794 5460 13806
rect 4732 13748 4788 13758
rect 4732 13654 4788 13692
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 7196 13076 7252 15092
rect 6972 13074 7252 13076
rect 6972 13022 7198 13074
rect 7250 13022 7252 13074
rect 6972 13020 7252 13022
rect 6076 12460 6468 12516
rect 6076 12178 6132 12460
rect 6412 12404 6468 12460
rect 6636 12404 6692 12414
rect 6412 12402 6692 12404
rect 6412 12350 6638 12402
rect 6690 12350 6692 12402
rect 6412 12348 6692 12350
rect 6636 12338 6692 12348
rect 6972 12404 7028 13020
rect 7196 13010 7252 13020
rect 6300 12292 6356 12302
rect 6300 12290 6468 12292
rect 6300 12238 6302 12290
rect 6354 12238 6468 12290
rect 6300 12236 6468 12238
rect 6300 12226 6356 12236
rect 6076 12126 6078 12178
rect 6130 12126 6132 12178
rect 6076 12114 6132 12126
rect 4844 12068 4900 12078
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4284 10446 4286 10498
rect 4338 10446 4340 10498
rect 4284 9268 4340 10446
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4732 9940 4788 9950
rect 4732 9846 4788 9884
rect 4284 9202 4340 9212
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 4620 2772 4676 2782
rect 4284 2770 4676 2772
rect 4284 2718 4622 2770
rect 4674 2718 4676 2770
rect 4284 2716 4676 2718
rect 3836 1876 3892 1886
rect 3836 1782 3892 1820
rect 4060 1874 4116 1886
rect 4060 1822 4062 1874
rect 4114 1822 4116 1874
rect 3388 1762 3444 1774
rect 3388 1710 3390 1762
rect 3442 1710 3444 1762
rect 3388 1204 3444 1710
rect 4060 1204 4116 1822
rect 4284 1876 4340 2716
rect 4620 2706 4676 2716
rect 4476 2380 4740 2390
rect 4532 2324 4580 2380
rect 4636 2324 4684 2380
rect 4476 2314 4740 2324
rect 4844 2212 4900 12012
rect 5740 11732 5796 11742
rect 5628 11396 5684 11406
rect 5292 11394 5684 11396
rect 5292 11342 5630 11394
rect 5682 11342 5684 11394
rect 5292 11340 5684 11342
rect 5292 10722 5348 11340
rect 5292 10670 5294 10722
rect 5346 10670 5348 10722
rect 5292 10658 5348 10670
rect 5516 9940 5572 11340
rect 5628 11330 5684 11340
rect 5740 10610 5796 11676
rect 6412 10722 6468 12236
rect 6972 12178 7028 12348
rect 7308 12292 7364 21084
rect 7420 21074 7476 21084
rect 7420 20804 7476 20814
rect 7420 20710 7476 20748
rect 7532 16772 7588 16782
rect 7532 15538 7588 16716
rect 7532 15486 7534 15538
rect 7586 15486 7588 15538
rect 7532 15316 7588 15486
rect 7532 15250 7588 15260
rect 7644 13748 7700 13758
rect 7532 13636 7588 13646
rect 6972 12126 6974 12178
rect 7026 12126 7028 12178
rect 6972 11506 7028 12126
rect 6972 11454 6974 11506
rect 7026 11454 7028 11506
rect 6972 11442 7028 11454
rect 7084 12236 7364 12292
rect 7420 13634 7588 13636
rect 7420 13582 7534 13634
rect 7586 13582 7588 13634
rect 7420 13580 7588 13582
rect 6412 10670 6414 10722
rect 6466 10670 6468 10722
rect 6412 10658 6468 10670
rect 5740 10558 5742 10610
rect 5794 10558 5796 10610
rect 5740 10546 5796 10558
rect 5516 9828 5572 9884
rect 5628 9828 5684 9838
rect 5516 9826 5684 9828
rect 5516 9774 5630 9826
rect 5682 9774 5684 9826
rect 5516 9772 5684 9774
rect 5628 9762 5684 9772
rect 5068 9716 5124 9726
rect 5068 8932 5124 9660
rect 7084 9716 7140 12236
rect 7196 12068 7252 12078
rect 7420 12068 7476 13580
rect 7532 13570 7588 13580
rect 7644 12964 7700 13692
rect 7196 12066 7476 12068
rect 7196 12014 7198 12066
rect 7250 12014 7476 12066
rect 7196 12012 7476 12014
rect 7532 12962 7700 12964
rect 7532 12910 7646 12962
rect 7698 12910 7700 12962
rect 7532 12908 7700 12910
rect 7196 10612 7252 12012
rect 7532 11732 7588 12908
rect 7644 12898 7700 12908
rect 7644 12068 7700 12078
rect 7644 11974 7700 12012
rect 7532 11666 7588 11676
rect 7196 10546 7252 10556
rect 7084 9650 7140 9660
rect 7420 9716 7476 9726
rect 7756 9716 7812 31164
rect 7420 9714 7812 9716
rect 7420 9662 7422 9714
rect 7474 9662 7812 9714
rect 7420 9660 7812 9662
rect 5292 8932 5348 8942
rect 5068 8930 5348 8932
rect 5068 8878 5294 8930
rect 5346 8878 5348 8930
rect 5068 8876 5348 8878
rect 5292 5236 5348 8876
rect 5964 7474 6020 7486
rect 5964 7422 5966 7474
rect 6018 7422 6020 7474
rect 5964 7252 6020 7422
rect 6636 7364 6692 7374
rect 6636 7270 6692 7308
rect 7420 7362 7476 9660
rect 7420 7310 7422 7362
rect 7474 7310 7476 7362
rect 5964 7186 6020 7196
rect 7420 7252 7476 7310
rect 7420 7186 7476 7196
rect 7308 6690 7364 6702
rect 7308 6638 7310 6690
rect 7362 6638 7364 6690
rect 7308 6580 7364 6638
rect 7308 6514 7364 6524
rect 7868 6468 7924 46396
rect 7980 45330 8036 46620
rect 7980 45278 7982 45330
rect 8034 45278 8036 45330
rect 7980 45266 8036 45278
rect 8092 44436 8148 60172
rect 8428 60002 8484 60014
rect 8428 59950 8430 60002
rect 8482 59950 8484 60002
rect 8428 59668 8484 59950
rect 8540 59890 8596 69244
rect 8764 68068 8820 69358
rect 9660 69188 9716 69198
rect 9772 69188 9828 70028
rect 9884 69990 9940 70028
rect 10108 70082 10164 70588
rect 10108 70030 10110 70082
rect 10162 70030 10164 70082
rect 9996 69188 10052 69198
rect 9716 69132 9828 69188
rect 9884 69186 10052 69188
rect 9884 69134 9998 69186
rect 10050 69134 10052 69186
rect 9884 69132 10052 69134
rect 9660 69122 9716 69132
rect 8988 68514 9044 68526
rect 8988 68462 8990 68514
rect 9042 68462 9044 68514
rect 8988 68404 9044 68462
rect 9548 68516 9604 68526
rect 9548 68422 9604 68460
rect 8988 68338 9044 68348
rect 9884 68402 9940 69132
rect 9996 69122 10052 69132
rect 10108 68740 10164 70030
rect 10332 70084 10388 70094
rect 10332 69990 10388 70028
rect 10108 68684 10388 68740
rect 10108 68516 10164 68526
rect 10108 68422 10164 68460
rect 9884 68350 9886 68402
rect 9938 68350 9940 68402
rect 9100 68292 9156 68302
rect 9324 68292 9380 68302
rect 8876 68068 8932 68078
rect 8764 68066 8932 68068
rect 8764 68014 8878 68066
rect 8930 68014 8932 68066
rect 8764 68012 8932 68014
rect 8764 67058 8820 68012
rect 8876 68002 8932 68012
rect 8764 67006 8766 67058
rect 8818 67006 8820 67058
rect 8764 66994 8820 67006
rect 8988 66946 9044 66958
rect 8988 66894 8990 66946
rect 9042 66894 9044 66946
rect 8764 66500 8820 66510
rect 8988 66500 9044 66894
rect 8652 66444 8764 66500
rect 8820 66444 9044 66500
rect 8652 66386 8708 66444
rect 8764 66434 8820 66444
rect 8652 66334 8654 66386
rect 8706 66334 8708 66386
rect 8652 66322 8708 66334
rect 8764 66276 8820 66286
rect 8652 62242 8708 62254
rect 8652 62190 8654 62242
rect 8706 62190 8708 62242
rect 8652 60004 8708 62190
rect 8652 59938 8708 59948
rect 8540 59838 8542 59890
rect 8594 59838 8596 59890
rect 8540 59826 8596 59838
rect 8764 59668 8820 66220
rect 9100 66274 9156 68236
rect 9212 68236 9324 68292
rect 9212 68066 9268 68236
rect 9324 68226 9380 68236
rect 9884 68292 9940 68350
rect 9884 68226 9940 68236
rect 9212 68014 9214 68066
rect 9266 68014 9268 68066
rect 9212 67954 9268 68014
rect 9212 67902 9214 67954
rect 9266 67902 9268 67954
rect 9212 67890 9268 67902
rect 9996 66500 10052 66510
rect 9996 66386 10052 66444
rect 9996 66334 9998 66386
rect 10050 66334 10052 66386
rect 9996 66322 10052 66334
rect 9100 66222 9102 66274
rect 9154 66222 9156 66274
rect 9100 66210 9156 66222
rect 9324 66276 9380 66286
rect 10220 66276 10276 66286
rect 9324 66182 9380 66220
rect 10108 66220 10220 66276
rect 9660 66052 9716 66062
rect 9660 65958 9716 65996
rect 10108 65828 10164 66220
rect 10220 66182 10276 66220
rect 9884 65772 10164 65828
rect 9884 65714 9940 65772
rect 9884 65662 9886 65714
rect 9938 65662 9940 65714
rect 9884 65650 9940 65662
rect 10332 65716 10388 68684
rect 10444 65828 10500 73892
rect 10556 73892 11060 73948
rect 11452 74676 11508 74686
rect 10556 68740 10612 73892
rect 11004 72324 11060 72334
rect 10780 72268 11004 72324
rect 10780 71090 10836 72268
rect 11004 72258 11060 72268
rect 11116 71764 11172 71774
rect 11116 71670 11172 71708
rect 10780 71038 10782 71090
rect 10834 71038 10836 71090
rect 10780 71026 10836 71038
rect 10668 70308 10724 70318
rect 10668 70306 11172 70308
rect 10668 70254 10670 70306
rect 10722 70254 11172 70306
rect 10668 70252 11172 70254
rect 10668 70242 10724 70252
rect 11004 70082 11060 70094
rect 11004 70030 11006 70082
rect 11058 70030 11060 70082
rect 10556 68674 10612 68684
rect 10668 69748 10724 69758
rect 10668 69522 10724 69692
rect 10668 69470 10670 69522
rect 10722 69470 10724 69522
rect 10556 68514 10612 68526
rect 10556 68462 10558 68514
rect 10610 68462 10612 68514
rect 10556 68292 10612 68462
rect 10556 67508 10612 68236
rect 10556 67442 10612 67452
rect 10668 66388 10724 69470
rect 10668 66322 10724 66332
rect 10892 68516 10948 68526
rect 10892 66386 10948 68460
rect 11004 66500 11060 70030
rect 11116 69748 11172 70252
rect 11228 69972 11284 69982
rect 11228 69878 11284 69916
rect 11116 69692 11284 69748
rect 11228 69410 11284 69692
rect 11228 69358 11230 69410
rect 11282 69358 11284 69410
rect 11228 69346 11284 69358
rect 11452 67956 11508 74620
rect 11788 72546 11844 72558
rect 13468 72548 13524 76300
rect 13580 74788 13636 77868
rect 13804 77364 13860 77374
rect 13804 77270 13860 77308
rect 13692 77140 13748 77150
rect 13692 77046 13748 77084
rect 13916 77026 13972 77038
rect 13916 76974 13918 77026
rect 13970 76974 13972 77026
rect 13916 75572 13972 76974
rect 13916 75506 13972 75516
rect 13692 74788 13748 74798
rect 13580 74732 13692 74788
rect 13692 74694 13748 74732
rect 14028 73948 14084 77868
rect 14196 77868 14308 77924
rect 14140 77252 14196 77868
rect 14476 77252 14532 77262
rect 14140 77250 14532 77252
rect 14140 77198 14478 77250
rect 14530 77198 14532 77250
rect 14140 77196 14532 77198
rect 14140 77138 14196 77196
rect 14140 77086 14142 77138
rect 14194 77086 14196 77138
rect 14140 77074 14196 77086
rect 14364 76354 14420 76366
rect 14364 76302 14366 76354
rect 14418 76302 14420 76354
rect 14364 74114 14420 76302
rect 14476 75684 14532 77196
rect 14812 77140 14868 78764
rect 14924 78818 14980 79772
rect 15372 79762 15428 79772
rect 14924 78766 14926 78818
rect 14978 78766 14980 78818
rect 14924 78754 14980 78766
rect 15036 78818 15092 78830
rect 15036 78766 15038 78818
rect 15090 78766 15092 78818
rect 15036 77362 15092 78766
rect 15820 78596 15876 78606
rect 15820 78148 15876 78540
rect 15820 78082 15876 78092
rect 15036 77310 15038 77362
rect 15090 77310 15092 77362
rect 15036 77298 15092 77310
rect 15260 77924 15316 77934
rect 14812 77074 14868 77084
rect 15148 77140 15204 77150
rect 15148 77046 15204 77084
rect 14924 77028 14980 77038
rect 14924 77026 15092 77028
rect 14924 76974 14926 77026
rect 14978 76974 15092 77026
rect 14924 76972 15092 76974
rect 14924 76962 14980 76972
rect 15036 76690 15092 76972
rect 15036 76638 15038 76690
rect 15090 76638 15092 76690
rect 15036 76020 15092 76638
rect 15036 75954 15092 75964
rect 14476 75618 14532 75628
rect 14588 75684 14644 75694
rect 15260 75684 15316 77868
rect 15484 77028 15540 77038
rect 15484 76690 15540 76972
rect 16044 77028 16100 86718
rect 16828 86770 16884 88958
rect 17500 89010 17556 89516
rect 19516 89572 19572 89582
rect 19516 89478 19572 89516
rect 19628 89124 19684 89740
rect 19964 89702 20020 89740
rect 19836 89404 20100 89414
rect 19892 89348 19940 89404
rect 19996 89348 20044 89404
rect 19836 89338 20100 89348
rect 19684 89068 19908 89124
rect 19628 89030 19684 89068
rect 17500 88958 17502 89010
rect 17554 88958 17556 89010
rect 17500 88946 17556 88958
rect 18284 88900 18340 88910
rect 18284 88806 18340 88844
rect 19516 88900 19572 88910
rect 19180 88788 19236 88798
rect 19068 88676 19124 88686
rect 16940 88340 16996 88350
rect 16940 88246 16996 88284
rect 17500 87668 17556 87678
rect 17500 87574 17556 87612
rect 18732 87668 18788 87678
rect 18172 87556 18228 87566
rect 18172 87554 18340 87556
rect 18172 87502 18174 87554
rect 18226 87502 18340 87554
rect 18172 87500 18340 87502
rect 18172 87490 18228 87500
rect 17836 87444 17892 87454
rect 17836 87350 17892 87388
rect 16828 86718 16830 86770
rect 16882 86718 16884 86770
rect 16828 86706 16884 86718
rect 18284 86772 18340 87500
rect 18732 87554 18788 87612
rect 18732 87502 18734 87554
rect 18786 87502 18788 87554
rect 18732 87490 18788 87502
rect 19068 87554 19124 88620
rect 19068 87502 19070 87554
rect 19122 87502 19124 87554
rect 19068 87490 19124 87502
rect 19180 88002 19236 88732
rect 19516 88226 19572 88844
rect 19516 88174 19518 88226
rect 19570 88174 19572 88226
rect 19516 88162 19572 88174
rect 19852 88226 19908 89068
rect 20636 89068 20804 89124
rect 20636 89012 20692 89068
rect 20412 88956 20692 89012
rect 20748 89010 20804 89068
rect 20748 88958 20750 89010
rect 20802 88958 20804 89010
rect 20412 88898 20468 88956
rect 20748 88946 20804 88958
rect 20412 88846 20414 88898
rect 20466 88846 20468 88898
rect 20412 88834 20468 88846
rect 19852 88174 19854 88226
rect 19906 88174 19908 88226
rect 19852 88162 19908 88174
rect 20636 88452 20692 88462
rect 20636 88226 20692 88396
rect 20636 88174 20638 88226
rect 20690 88174 20692 88226
rect 20636 88162 20692 88174
rect 19180 87950 19182 88002
rect 19234 87950 19236 88002
rect 19180 86772 19236 87950
rect 19740 88004 19796 88042
rect 19740 87938 19796 87948
rect 20188 88004 20244 88014
rect 20300 88004 20356 88014
rect 20244 88002 20356 88004
rect 20244 87950 20302 88002
rect 20354 87950 20356 88002
rect 20244 87948 20356 87950
rect 19836 87836 20100 87846
rect 19892 87780 19940 87836
rect 19996 87780 20044 87836
rect 19836 87770 20100 87780
rect 20076 87668 20132 87678
rect 20076 87574 20132 87612
rect 18284 86770 19236 86772
rect 18284 86718 18286 86770
rect 18338 86718 19182 86770
rect 19234 86718 19236 86770
rect 18284 86716 19236 86718
rect 16940 86660 16996 86670
rect 16940 86566 16996 86604
rect 17500 86660 17556 86670
rect 18284 86660 18340 86716
rect 19180 86706 19236 86716
rect 19628 87444 19684 87454
rect 19684 87388 19908 87444
rect 17500 86658 18340 86660
rect 17500 86606 17502 86658
rect 17554 86606 18340 86658
rect 17500 86604 18340 86606
rect 17500 85708 17556 86604
rect 19628 86100 19684 87388
rect 19852 86770 19908 87388
rect 19852 86718 19854 86770
rect 19906 86718 19908 86770
rect 19852 86706 19908 86718
rect 19836 86268 20100 86278
rect 19892 86212 19940 86268
rect 19996 86212 20044 86268
rect 19836 86202 20100 86212
rect 19628 86044 19908 86100
rect 19628 85762 19684 85774
rect 19628 85710 19630 85762
rect 19682 85710 19684 85762
rect 17500 85652 18004 85708
rect 17612 84532 17668 84542
rect 17612 84438 17668 84476
rect 16156 84084 16212 84094
rect 16156 83634 16212 84028
rect 16156 83582 16158 83634
rect 16210 83582 16212 83634
rect 16156 83076 16212 83582
rect 17724 83748 17780 83758
rect 17724 83634 17780 83692
rect 17724 83582 17726 83634
rect 17778 83582 17780 83634
rect 17724 83570 17780 83582
rect 17836 83522 17892 83534
rect 17836 83470 17838 83522
rect 17890 83470 17892 83522
rect 17836 83412 17892 83470
rect 16604 83300 16660 83310
rect 16604 83206 16660 83244
rect 17164 83300 17220 83310
rect 17164 83206 17220 83244
rect 17836 83076 17892 83356
rect 16156 83010 16212 83020
rect 17612 83020 17892 83076
rect 17612 82962 17668 83020
rect 17612 82910 17614 82962
rect 17666 82910 17668 82962
rect 17612 82898 17668 82910
rect 16940 82516 16996 82526
rect 16380 82292 16436 82302
rect 16380 81060 16436 82236
rect 16940 81394 16996 82460
rect 17388 81954 17444 81966
rect 17388 81902 17390 81954
rect 17442 81902 17444 81954
rect 16940 81342 16942 81394
rect 16994 81342 16996 81394
rect 16940 81330 16996 81342
rect 17052 81730 17108 81742
rect 17052 81678 17054 81730
rect 17106 81678 17108 81730
rect 16268 79828 16324 79838
rect 16268 79492 16324 79772
rect 16380 79492 16436 81004
rect 16492 81284 16548 81294
rect 16492 80386 16548 81228
rect 17052 81060 17108 81678
rect 17052 80994 17108 81004
rect 17388 81170 17444 81902
rect 17388 81118 17390 81170
rect 17442 81118 17444 81170
rect 17388 81060 17444 81118
rect 17388 80994 17444 81004
rect 17388 80612 17444 80622
rect 17388 80518 17444 80556
rect 17052 80500 17108 80510
rect 17052 80406 17108 80444
rect 17836 80388 17892 80398
rect 16492 80334 16494 80386
rect 16546 80334 16548 80386
rect 16492 80322 16548 80334
rect 17724 80332 17836 80388
rect 17612 80276 17668 80286
rect 17500 80274 17668 80276
rect 17500 80222 17614 80274
rect 17666 80222 17668 80274
rect 17500 80220 17668 80222
rect 16268 79490 16436 79492
rect 16268 79438 16382 79490
rect 16434 79438 16436 79490
rect 16268 79436 16436 79438
rect 16268 78818 16324 79436
rect 16380 79426 16436 79436
rect 16716 80162 16772 80174
rect 16716 80110 16718 80162
rect 16770 80110 16772 80162
rect 16268 78766 16270 78818
rect 16322 78766 16324 78818
rect 16044 76962 16100 76972
rect 16156 77922 16212 77934
rect 16156 77870 16158 77922
rect 16210 77870 16212 77922
rect 16156 76804 16212 77870
rect 16268 77924 16324 78766
rect 16716 78372 16772 80110
rect 16828 79492 16884 79502
rect 16828 79398 16884 79436
rect 17500 78932 17556 80220
rect 17612 80210 17668 80220
rect 17612 79828 17668 79838
rect 17724 79828 17780 80332
rect 17836 80322 17892 80332
rect 17948 80052 18004 85652
rect 19068 85314 19124 85326
rect 19068 85262 19070 85314
rect 19122 85262 19124 85314
rect 18844 85204 18900 85214
rect 18732 84868 18788 84878
rect 18732 84774 18788 84812
rect 18844 84532 18900 85148
rect 18844 84438 18900 84476
rect 19068 84530 19124 85262
rect 19628 85314 19684 85710
rect 19852 85708 19908 86044
rect 19852 85652 20132 85708
rect 19628 85262 19630 85314
rect 19682 85262 19684 85314
rect 19628 85250 19684 85262
rect 19068 84478 19070 84530
rect 19122 84478 19124 84530
rect 19068 84466 19124 84478
rect 19180 85092 19236 85102
rect 18508 84308 18564 84318
rect 18844 84308 18900 84318
rect 18508 84306 18844 84308
rect 18508 84254 18510 84306
rect 18562 84254 18844 84306
rect 18508 84252 18844 84254
rect 18508 84242 18564 84252
rect 18060 84194 18116 84206
rect 18060 84142 18062 84194
rect 18114 84142 18116 84194
rect 18060 83412 18116 84142
rect 18732 84082 18788 84094
rect 18732 84030 18734 84082
rect 18786 84030 18788 84082
rect 18396 83524 18452 83534
rect 18060 83346 18116 83356
rect 18172 83522 18452 83524
rect 18172 83470 18398 83522
rect 18450 83470 18452 83522
rect 18172 83468 18452 83470
rect 18172 82852 18228 83468
rect 18396 83458 18452 83468
rect 18508 83524 18564 83534
rect 18508 83430 18564 83468
rect 18284 83300 18340 83310
rect 18284 83206 18340 83244
rect 18732 83076 18788 84030
rect 18060 82796 18228 82852
rect 18284 83020 18788 83076
rect 18060 82068 18116 82796
rect 18172 82626 18228 82638
rect 18172 82574 18174 82626
rect 18226 82574 18228 82626
rect 18172 82516 18228 82574
rect 18172 82450 18228 82460
rect 18172 82068 18228 82078
rect 18060 82066 18228 82068
rect 18060 82014 18174 82066
rect 18226 82014 18228 82066
rect 18060 82012 18228 82014
rect 18172 82002 18228 82012
rect 18172 81284 18228 81294
rect 18284 81284 18340 83020
rect 18844 82964 18900 84252
rect 19180 83748 19236 85036
rect 19740 84868 19796 84878
rect 19628 84866 19796 84868
rect 19628 84814 19742 84866
rect 19794 84814 19796 84866
rect 19628 84812 19796 84814
rect 19180 83522 19236 83692
rect 19404 84306 19460 84318
rect 19404 84254 19406 84306
rect 19458 84254 19460 84306
rect 19292 83636 19348 83646
rect 19292 83542 19348 83580
rect 19180 83470 19182 83522
rect 19234 83470 19236 83522
rect 19180 83458 19236 83470
rect 18732 82908 18900 82964
rect 19292 83412 19348 83422
rect 18620 82850 18676 82862
rect 18620 82798 18622 82850
rect 18674 82798 18676 82850
rect 18172 81282 18340 81284
rect 18172 81230 18174 81282
rect 18226 81230 18340 81282
rect 18172 81228 18340 81230
rect 18396 82516 18452 82526
rect 18172 81218 18228 81228
rect 18396 81060 18452 82460
rect 18508 82514 18564 82526
rect 18508 82462 18510 82514
rect 18562 82462 18564 82514
rect 18508 81284 18564 82462
rect 18508 81218 18564 81228
rect 18060 81004 18452 81060
rect 18620 81060 18676 82798
rect 18060 80274 18116 81004
rect 18620 80994 18676 81004
rect 18060 80222 18062 80274
rect 18114 80222 18116 80274
rect 18060 80210 18116 80222
rect 17948 79996 18228 80052
rect 18060 79828 18116 79838
rect 17612 79826 17780 79828
rect 17612 79774 17614 79826
rect 17666 79774 17780 79826
rect 17612 79772 17780 79774
rect 17948 79772 18060 79828
rect 17612 79762 17668 79772
rect 17948 79714 18004 79772
rect 18060 79762 18116 79772
rect 17948 79662 17950 79714
rect 18002 79662 18004 79714
rect 17948 79650 18004 79662
rect 17500 78866 17556 78876
rect 18060 79492 18116 79502
rect 16940 78708 16996 78718
rect 16940 78706 17780 78708
rect 16940 78654 16942 78706
rect 16994 78654 17780 78706
rect 16940 78652 17780 78654
rect 16940 78642 16996 78652
rect 16716 78306 16772 78316
rect 17724 78258 17780 78652
rect 17724 78206 17726 78258
rect 17778 78206 17780 78258
rect 17724 78194 17780 78206
rect 17612 78148 17668 78158
rect 17612 78054 17668 78092
rect 16268 77858 16324 77868
rect 16716 78036 16772 78046
rect 16156 76748 16324 76804
rect 15484 76638 15486 76690
rect 15538 76638 15540 76690
rect 15484 76626 15540 76638
rect 15932 76692 15988 76702
rect 15932 76598 15988 76636
rect 16156 76466 16212 76478
rect 16156 76414 16158 76466
rect 16210 76414 16212 76466
rect 14588 75682 15316 75684
rect 14588 75630 14590 75682
rect 14642 75630 15316 75682
rect 14588 75628 15316 75630
rect 15932 75684 15988 75694
rect 16156 75684 16212 76414
rect 15988 75628 16212 75684
rect 16268 75682 16324 76748
rect 16604 76692 16660 76702
rect 16604 76598 16660 76636
rect 16716 76690 16772 77980
rect 17388 78036 17444 78046
rect 17388 77942 17444 77980
rect 17948 78034 18004 78046
rect 17948 77982 17950 78034
rect 18002 77982 18004 78034
rect 16828 77924 16884 77934
rect 16828 77830 16884 77868
rect 16716 76638 16718 76690
rect 16770 76638 16772 76690
rect 16716 76626 16772 76638
rect 16828 77140 16884 77150
rect 16828 76692 16884 77084
rect 17948 77140 18004 77982
rect 17948 77074 18004 77084
rect 17724 77028 17780 77038
rect 16828 76690 17332 76692
rect 16828 76638 16830 76690
rect 16882 76638 17332 76690
rect 16828 76636 17332 76638
rect 16828 76626 16884 76636
rect 17276 76466 17332 76636
rect 17724 76578 17780 76972
rect 17724 76526 17726 76578
rect 17778 76526 17780 76578
rect 17724 76514 17780 76526
rect 17276 76414 17278 76466
rect 17330 76414 17332 76466
rect 17276 76402 17332 76414
rect 17836 76466 17892 76478
rect 17836 76414 17838 76466
rect 17890 76414 17892 76466
rect 16268 75630 16270 75682
rect 16322 75630 16324 75682
rect 14588 75618 14644 75628
rect 14364 74062 14366 74114
rect 14418 74062 14420 74114
rect 14364 74050 14420 74062
rect 15036 75460 15092 75470
rect 13804 73892 14084 73948
rect 15036 74004 15092 75404
rect 15036 73938 15092 73948
rect 13692 72548 13748 72558
rect 11788 72494 11790 72546
rect 11842 72494 11844 72546
rect 11564 72324 11620 72334
rect 11564 72230 11620 72268
rect 11788 71876 11844 72494
rect 11564 71820 11844 71876
rect 13356 72492 13524 72548
rect 13580 72546 13748 72548
rect 13580 72494 13694 72546
rect 13746 72494 13748 72546
rect 13580 72492 13748 72494
rect 11564 70418 11620 71820
rect 11788 71652 11844 71662
rect 11564 70366 11566 70418
rect 11618 70366 11620 70418
rect 11564 70354 11620 70366
rect 11676 71650 11844 71652
rect 11676 71598 11790 71650
rect 11842 71598 11844 71650
rect 11676 71596 11844 71598
rect 11564 69300 11620 69310
rect 11676 69300 11732 71596
rect 11788 71586 11844 71596
rect 12684 71428 12740 71438
rect 11900 70868 11956 70878
rect 11900 70194 11956 70812
rect 12684 70306 12740 71372
rect 12908 71090 12964 71102
rect 12908 71038 12910 71090
rect 12962 71038 12964 71090
rect 12908 70644 12964 71038
rect 13356 70980 13412 72492
rect 13468 72322 13524 72334
rect 13468 72270 13470 72322
rect 13522 72270 13524 72322
rect 13468 71428 13524 72270
rect 13468 71362 13524 71372
rect 13468 71204 13524 71214
rect 13580 71204 13636 72492
rect 13692 72482 13748 72492
rect 13804 71204 13860 73892
rect 13916 73218 13972 73230
rect 13916 73166 13918 73218
rect 13970 73166 13972 73218
rect 13916 72212 13972 73166
rect 15148 72658 15204 75628
rect 15148 72606 15150 72658
rect 15202 72606 15204 72658
rect 15148 72594 15204 72606
rect 15260 74788 15316 74798
rect 13916 72146 13972 72156
rect 14476 71764 14532 71774
rect 14476 71670 14532 71708
rect 15036 71764 15092 71774
rect 13916 71652 13972 71662
rect 13916 71650 14420 71652
rect 13916 71598 13918 71650
rect 13970 71598 14420 71650
rect 13916 71596 14420 71598
rect 13916 71586 13972 71596
rect 13468 71202 13636 71204
rect 13468 71150 13470 71202
rect 13522 71150 13636 71202
rect 13468 71148 13636 71150
rect 13692 71202 13860 71204
rect 13692 71150 13806 71202
rect 13858 71150 13860 71202
rect 13692 71148 13860 71150
rect 13468 71138 13524 71148
rect 13356 70924 13524 70980
rect 12908 70578 12964 70588
rect 12684 70254 12686 70306
rect 12738 70254 12740 70306
rect 12684 70242 12740 70254
rect 11900 70142 11902 70194
rect 11954 70142 11956 70194
rect 11900 69524 11956 70142
rect 11900 69458 11956 69468
rect 11564 69298 11732 69300
rect 11564 69246 11566 69298
rect 11618 69246 11732 69298
rect 11564 69244 11732 69246
rect 11564 69234 11620 69244
rect 11116 67900 11508 67956
rect 13468 68404 13524 70924
rect 13692 69972 13748 71148
rect 13804 71138 13860 71148
rect 14364 71092 14420 71596
rect 14476 71092 14532 71102
rect 14364 71090 14532 71092
rect 14364 71038 14478 71090
rect 14530 71038 14532 71090
rect 14364 71036 14532 71038
rect 14476 71026 14532 71036
rect 14028 70978 14084 70990
rect 14028 70926 14030 70978
rect 14082 70926 14084 70978
rect 14028 70644 14084 70926
rect 15036 70978 15092 71708
rect 15036 70926 15038 70978
rect 15090 70926 15092 70978
rect 14028 70578 14084 70588
rect 14588 70754 14644 70766
rect 14588 70702 14590 70754
rect 14642 70702 14644 70754
rect 14588 70308 14644 70702
rect 14588 70242 14644 70252
rect 14812 70084 14868 70094
rect 13580 69524 13636 69534
rect 13692 69524 13748 69916
rect 14700 70082 14868 70084
rect 14700 70030 14814 70082
rect 14866 70030 14868 70082
rect 14700 70028 14868 70030
rect 14028 69524 14084 69534
rect 13580 69522 13972 69524
rect 13580 69470 13582 69522
rect 13634 69470 13972 69522
rect 13580 69468 13972 69470
rect 13580 69458 13636 69468
rect 11116 67172 11172 67900
rect 11676 67508 11732 67518
rect 11116 67170 11396 67172
rect 11116 67118 11118 67170
rect 11170 67118 11396 67170
rect 11116 67116 11396 67118
rect 11116 67106 11172 67116
rect 11004 66444 11284 66500
rect 10892 66334 10894 66386
rect 10946 66334 10948 66386
rect 10892 66322 10948 66334
rect 11116 66276 11172 66286
rect 11004 66220 11116 66276
rect 10556 66052 10612 66062
rect 10556 65958 10612 65996
rect 11004 65828 11060 66220
rect 11116 66182 11172 66220
rect 10444 65772 10612 65828
rect 10332 65660 10500 65716
rect 8876 65378 8932 65390
rect 8876 65326 8878 65378
rect 8930 65326 8932 65378
rect 8876 63700 8932 65326
rect 8932 63644 9044 63700
rect 8876 63634 8932 63644
rect 8988 63140 9044 63644
rect 8988 63046 9044 63084
rect 9212 63364 9268 63374
rect 8428 59612 8820 59668
rect 8988 61684 9044 61694
rect 8316 59108 8372 59118
rect 8428 59108 8484 59612
rect 8988 59442 9044 61628
rect 9100 61348 9156 61358
rect 9100 61254 9156 61292
rect 9100 60116 9156 60126
rect 9212 60116 9268 63308
rect 9660 63140 9716 63150
rect 9660 62580 9716 63084
rect 9772 63028 9828 63038
rect 9772 63026 10052 63028
rect 9772 62974 9774 63026
rect 9826 62974 10052 63026
rect 9772 62972 10052 62974
rect 9772 62962 9828 62972
rect 9660 62486 9716 62524
rect 9996 62578 10052 62972
rect 9996 62526 9998 62578
rect 10050 62526 10052 62578
rect 9996 62514 10052 62526
rect 10332 62354 10388 62366
rect 10332 62302 10334 62354
rect 10386 62302 10388 62354
rect 9996 61684 10052 61694
rect 9772 61628 9996 61684
rect 9548 60900 9604 60910
rect 9100 60114 9268 60116
rect 9100 60062 9102 60114
rect 9154 60062 9268 60114
rect 9100 60060 9268 60062
rect 9324 60898 9604 60900
rect 9324 60846 9550 60898
rect 9602 60846 9604 60898
rect 9324 60844 9604 60846
rect 9100 60050 9156 60060
rect 8988 59390 8990 59442
rect 9042 59390 9044 59442
rect 8988 59378 9044 59390
rect 8540 59108 8596 59118
rect 8428 59106 8596 59108
rect 8428 59054 8542 59106
rect 8594 59054 8596 59106
rect 8428 59052 8596 59054
rect 8316 58884 8372 59052
rect 8316 58828 8484 58884
rect 8428 58434 8484 58828
rect 8428 58382 8430 58434
rect 8482 58382 8484 58434
rect 8428 58212 8484 58382
rect 8428 58146 8484 58156
rect 8204 57652 8260 57662
rect 8204 56532 8260 57596
rect 8204 53954 8260 56476
rect 8540 55412 8596 59052
rect 9100 58548 9156 58558
rect 9324 58548 9380 60844
rect 9548 60834 9604 60844
rect 9548 60004 9604 60014
rect 9548 59330 9604 59948
rect 9548 59278 9550 59330
rect 9602 59278 9604 59330
rect 9548 59266 9604 59278
rect 9772 59218 9828 61628
rect 9996 61590 10052 61628
rect 10332 61010 10388 62302
rect 10332 60958 10334 61010
rect 10386 60958 10388 61010
rect 10332 60946 10388 60958
rect 9884 60788 9940 60798
rect 9884 60786 10052 60788
rect 9884 60734 9886 60786
rect 9938 60734 10052 60786
rect 9884 60732 10052 60734
rect 9884 60722 9940 60732
rect 9996 59444 10052 60732
rect 10108 59444 10164 59454
rect 9996 59442 10164 59444
rect 9996 59390 10110 59442
rect 10162 59390 10164 59442
rect 9996 59388 10164 59390
rect 10108 59378 10164 59388
rect 9772 59166 9774 59218
rect 9826 59166 9828 59218
rect 9772 59154 9828 59166
rect 9100 58546 9380 58548
rect 9100 58494 9102 58546
rect 9154 58494 9380 58546
rect 9100 58492 9380 58494
rect 9100 58482 9156 58492
rect 9772 58212 9828 58222
rect 8540 55346 8596 55356
rect 8652 55410 8708 55422
rect 8652 55358 8654 55410
rect 8706 55358 8708 55410
rect 8428 54516 8484 54526
rect 8204 53902 8206 53954
rect 8258 53902 8260 53954
rect 8204 53732 8260 53902
rect 8204 53666 8260 53676
rect 8316 54460 8428 54516
rect 8204 53060 8260 53070
rect 8316 53060 8372 54460
rect 8428 54450 8484 54460
rect 8652 54180 8708 55358
rect 9772 55410 9828 58156
rect 9772 55358 9774 55410
rect 9826 55358 9828 55410
rect 9772 55346 9828 55358
rect 9324 55076 9380 55086
rect 9324 54982 9380 55020
rect 9548 54628 9604 54638
rect 9548 54534 9604 54572
rect 10444 54626 10500 65660
rect 10444 54574 10446 54626
rect 10498 54574 10500 54626
rect 10444 54562 10500 54574
rect 8988 54516 9044 54526
rect 9772 54516 9828 54526
rect 8988 54402 9044 54460
rect 8988 54350 8990 54402
rect 9042 54350 9044 54402
rect 8988 54338 9044 54350
rect 9660 54514 9828 54516
rect 9660 54462 9774 54514
rect 9826 54462 9828 54514
rect 9660 54460 9828 54462
rect 8428 54124 8708 54180
rect 8428 53620 8484 54124
rect 9660 54068 9716 54460
rect 9772 54450 9828 54460
rect 8540 54012 9716 54068
rect 10444 54402 10500 54414
rect 10444 54350 10446 54402
rect 10498 54350 10500 54402
rect 8540 53954 8596 54012
rect 8540 53902 8542 53954
rect 8594 53902 8596 53954
rect 8540 53890 8596 53902
rect 8428 53554 8484 53564
rect 8652 53732 8708 53742
rect 8652 53172 8708 53676
rect 8988 53732 9044 53742
rect 8988 53638 9044 53676
rect 10108 53730 10164 53742
rect 10108 53678 10110 53730
rect 10162 53678 10164 53730
rect 9660 53620 9716 53630
rect 8652 53170 8820 53172
rect 8652 53118 8654 53170
rect 8706 53118 8820 53170
rect 8652 53116 8820 53118
rect 8652 53106 8708 53116
rect 8204 53058 8372 53060
rect 8204 53006 8206 53058
rect 8258 53006 8372 53058
rect 8204 53004 8372 53006
rect 8204 52994 8260 53004
rect 8204 52612 8260 52622
rect 8204 49698 8260 52556
rect 8204 49646 8206 49698
rect 8258 49646 8260 49698
rect 8204 49586 8260 49646
rect 8204 49534 8206 49586
rect 8258 49534 8260 49586
rect 8204 49522 8260 49534
rect 8316 52500 8372 52510
rect 8316 49364 8372 52444
rect 8204 49308 8372 49364
rect 8204 44548 8260 49308
rect 8316 49138 8372 49150
rect 8316 49086 8318 49138
rect 8370 49086 8372 49138
rect 8316 48692 8372 49086
rect 8316 48626 8372 48636
rect 8764 48020 8820 53116
rect 9324 51268 9380 51278
rect 9324 50594 9380 51212
rect 9436 50708 9492 50718
rect 9436 50614 9492 50652
rect 9324 50542 9326 50594
rect 9378 50542 9380 50594
rect 8876 50482 8932 50494
rect 8876 50430 8878 50482
rect 8930 50430 8932 50482
rect 8876 49252 8932 50430
rect 9324 50428 9380 50542
rect 9660 50594 9716 53564
rect 10108 53508 10164 53678
rect 10108 53442 10164 53452
rect 9660 50542 9662 50594
rect 9714 50542 9716 50594
rect 9660 50530 9716 50542
rect 10220 52052 10276 52062
rect 10220 50428 10276 51996
rect 9324 50372 9716 50428
rect 8932 49196 9044 49252
rect 8876 49186 8932 49196
rect 8876 48132 8932 48142
rect 8876 48038 8932 48076
rect 8764 47954 8820 47964
rect 8988 47570 9044 49196
rect 9660 48580 9716 50372
rect 10108 50372 10276 50428
rect 10108 50370 10164 50372
rect 10108 50318 10110 50370
rect 10162 50318 10164 50370
rect 10108 50036 10164 50318
rect 10444 50036 10500 54350
rect 10556 51044 10612 65772
rect 10780 65772 11060 65828
rect 10780 65714 10836 65772
rect 10780 65662 10782 65714
rect 10834 65662 10836 65714
rect 10780 65650 10836 65662
rect 11228 63812 11284 66444
rect 11228 63746 11284 63756
rect 10668 61684 10724 61694
rect 10668 60786 10724 61628
rect 10668 60734 10670 60786
rect 10722 60734 10724 60786
rect 10668 60722 10724 60734
rect 10892 60674 10948 60686
rect 10892 60622 10894 60674
rect 10946 60622 10948 60674
rect 10892 60564 10948 60622
rect 11116 60564 11172 60574
rect 10892 60562 11172 60564
rect 10892 60510 11118 60562
rect 11170 60510 11172 60562
rect 10892 60508 11172 60510
rect 11116 60498 11172 60508
rect 11228 59892 11284 59902
rect 11004 59890 11284 59892
rect 11004 59838 11230 59890
rect 11282 59838 11284 59890
rect 11004 59836 11284 59838
rect 10892 59220 10948 59230
rect 10892 59126 10948 59164
rect 10892 57876 10948 57886
rect 11004 57876 11060 59836
rect 11228 59826 11284 59836
rect 11340 58772 11396 67116
rect 11452 66050 11508 66062
rect 11452 65998 11454 66050
rect 11506 65998 11508 66050
rect 11452 65716 11508 65998
rect 11452 65650 11508 65660
rect 11452 64260 11508 64270
rect 11452 63922 11508 64204
rect 11452 63870 11454 63922
rect 11506 63870 11508 63922
rect 11452 63858 11508 63870
rect 11676 62188 11732 67452
rect 11900 66276 11956 66286
rect 11900 66050 11956 66220
rect 11900 65998 11902 66050
rect 11954 65998 11956 66050
rect 11788 65490 11844 65502
rect 11788 65438 11790 65490
rect 11842 65438 11844 65490
rect 11788 64260 11844 65438
rect 11900 64372 11956 65998
rect 12460 65380 12516 65390
rect 12460 65286 12516 65324
rect 12460 64932 12516 64942
rect 12460 64818 12516 64876
rect 13468 64932 13524 68348
rect 13468 64838 13524 64876
rect 13580 65380 13636 65390
rect 12460 64766 12462 64818
rect 12514 64766 12516 64818
rect 12460 64754 12516 64766
rect 13020 64820 13076 64830
rect 13020 64726 13076 64764
rect 13580 64818 13636 65324
rect 13580 64766 13582 64818
rect 13634 64766 13636 64818
rect 13580 64754 13636 64766
rect 13692 64820 13748 64830
rect 13692 64596 13748 64764
rect 13804 64708 13860 64718
rect 13804 64614 13860 64652
rect 13580 64540 13748 64596
rect 11900 64306 11956 64316
rect 12124 64484 12180 64494
rect 11788 64194 11844 64204
rect 12124 64034 12180 64428
rect 12124 63982 12126 64034
rect 12178 63982 12180 64034
rect 12124 63970 12180 63982
rect 11900 63812 11956 63822
rect 11900 63252 11956 63756
rect 11900 63158 11956 63196
rect 13468 63364 13524 63374
rect 13468 63250 13524 63308
rect 13468 63198 13470 63250
rect 13522 63198 13524 63250
rect 13468 63186 13524 63198
rect 12348 62914 12404 62926
rect 12348 62862 12350 62914
rect 12402 62862 12404 62914
rect 11564 62132 11732 62188
rect 12012 62580 12068 62590
rect 12348 62580 12404 62862
rect 12068 62524 12404 62580
rect 10892 57874 11060 57876
rect 10892 57822 10894 57874
rect 10946 57822 11060 57874
rect 10892 57820 11060 57822
rect 11116 58716 11396 58772
rect 11452 60674 11508 60686
rect 11452 60622 11454 60674
rect 11506 60622 11508 60674
rect 11452 60562 11508 60622
rect 11452 60510 11454 60562
rect 11506 60510 11508 60562
rect 10892 57810 10948 57820
rect 10668 57652 10724 57662
rect 10668 57650 10836 57652
rect 10668 57598 10670 57650
rect 10722 57598 10836 57650
rect 10668 57596 10836 57598
rect 10668 57586 10724 57596
rect 10780 56756 10836 57596
rect 11116 56868 11172 58716
rect 11228 58548 11284 58558
rect 11452 58548 11508 60510
rect 11228 58546 11508 58548
rect 11228 58494 11230 58546
rect 11282 58494 11508 58546
rect 11228 58492 11508 58494
rect 11228 58482 11284 58492
rect 11116 56812 11396 56868
rect 10780 56700 11284 56756
rect 11228 56306 11284 56700
rect 11228 56254 11230 56306
rect 11282 56254 11284 56306
rect 11228 56242 11284 56254
rect 10892 55412 10948 55422
rect 10892 54514 10948 55356
rect 10892 54462 10894 54514
rect 10946 54462 10948 54514
rect 10892 53956 10948 54462
rect 11228 54516 11284 54526
rect 11228 54422 11284 54460
rect 10892 53890 10948 53900
rect 10780 53844 10836 53854
rect 10780 53750 10836 53788
rect 10780 51268 10836 51278
rect 10780 51174 10836 51212
rect 10556 50988 10836 51044
rect 10780 50428 10836 50988
rect 11340 50708 11396 56812
rect 11452 54852 11508 58492
rect 11564 56084 11620 62132
rect 12012 60116 12068 62524
rect 13580 61460 13636 64540
rect 13692 64372 13748 64382
rect 13692 63138 13748 64316
rect 13692 63086 13694 63138
rect 13746 63086 13748 63138
rect 13692 62580 13748 63086
rect 13916 62804 13972 69468
rect 14028 69430 14084 69468
rect 14476 69524 14532 69534
rect 14476 69430 14532 69468
rect 14364 68740 14420 68750
rect 14252 66162 14308 66174
rect 14252 66110 14254 66162
rect 14306 66110 14308 66162
rect 14140 66052 14196 66062
rect 14028 66050 14196 66052
rect 14028 65998 14142 66050
rect 14194 65998 14196 66050
rect 14028 65996 14196 65998
rect 14028 65492 14084 65996
rect 14140 65986 14196 65996
rect 14028 64708 14084 65436
rect 14252 64708 14308 66110
rect 14028 64642 14084 64652
rect 14140 64652 14308 64708
rect 14364 64820 14420 68684
rect 14364 64706 14420 64764
rect 14364 64654 14366 64706
rect 14418 64654 14420 64706
rect 14028 64484 14084 64494
rect 14028 64390 14084 64428
rect 14028 64036 14084 64046
rect 14028 63362 14084 63980
rect 14140 63812 14196 64652
rect 14364 64642 14420 64654
rect 14588 65378 14644 65390
rect 14588 65326 14590 65378
rect 14642 65326 14644 65378
rect 14252 64484 14308 64494
rect 14252 64482 14420 64484
rect 14252 64430 14254 64482
rect 14306 64430 14420 64482
rect 14252 64428 14420 64430
rect 14252 64418 14308 64428
rect 14364 63924 14420 64428
rect 14588 64034 14644 65326
rect 14588 63982 14590 64034
rect 14642 63982 14644 64034
rect 14588 63970 14644 63982
rect 14700 63924 14756 70028
rect 14812 70018 14868 70028
rect 14812 69524 14868 69534
rect 14812 69410 14868 69468
rect 14812 69358 14814 69410
rect 14866 69358 14868 69410
rect 14812 69346 14868 69358
rect 15036 68964 15092 70926
rect 15260 70418 15316 74732
rect 15260 70366 15262 70418
rect 15314 70366 15316 70418
rect 15260 70196 15316 70366
rect 15036 68908 15204 68964
rect 14924 68852 14980 68862
rect 14812 68796 14924 68852
rect 14812 66386 14868 68796
rect 14924 68786 14980 68796
rect 15148 68852 15204 68908
rect 15148 68786 15204 68796
rect 15260 68740 15316 70140
rect 15372 74004 15428 74014
rect 15820 74002 15876 74014
rect 15820 73950 15822 74002
rect 15874 73950 15876 74002
rect 15820 73948 15876 73950
rect 15372 73892 15876 73948
rect 15932 74004 15988 75628
rect 16268 75618 16324 75630
rect 17500 76354 17556 76366
rect 17500 76302 17502 76354
rect 17554 76302 17556 76354
rect 15932 73938 15988 73948
rect 16044 75124 16100 75134
rect 15372 68740 15428 73892
rect 16044 73442 16100 75068
rect 17500 75124 17556 76302
rect 17500 75058 17556 75068
rect 17724 75124 17780 75134
rect 17724 75030 17780 75068
rect 17500 73892 17556 73902
rect 17500 73554 17556 73836
rect 17500 73502 17502 73554
rect 17554 73502 17556 73554
rect 17500 73490 17556 73502
rect 17836 73554 17892 76414
rect 18060 75572 18116 79436
rect 18060 75506 18116 75516
rect 18172 75124 18228 79996
rect 18284 79604 18340 79614
rect 18284 79510 18340 79548
rect 18620 79604 18676 79614
rect 18620 79510 18676 79548
rect 18396 79490 18452 79502
rect 18396 79438 18398 79490
rect 18450 79438 18452 79490
rect 18396 78820 18452 79438
rect 18732 79380 18788 82908
rect 18844 82514 18900 82526
rect 18844 82462 18846 82514
rect 18898 82462 18900 82514
rect 18844 80724 18900 82462
rect 18844 80658 18900 80668
rect 19292 80610 19348 83356
rect 19404 82628 19460 84254
rect 19628 84084 19684 84812
rect 19740 84802 19796 84812
rect 20076 84868 20132 85652
rect 20188 85092 20244 87948
rect 20300 87938 20356 87948
rect 20748 88002 20804 88014
rect 20748 87950 20750 88002
rect 20802 87950 20804 88002
rect 20412 87780 20468 87790
rect 20300 86658 20356 86670
rect 20300 86606 20302 86658
rect 20354 86606 20356 86658
rect 20300 85092 20356 86606
rect 20412 86546 20468 87724
rect 20636 87442 20692 87454
rect 20636 87390 20638 87442
rect 20690 87390 20692 87442
rect 20636 86772 20692 87390
rect 20748 86884 20804 87950
rect 20748 86818 20804 86828
rect 20636 86706 20692 86716
rect 20748 86660 20804 86670
rect 20748 86566 20804 86604
rect 20412 86494 20414 86546
rect 20466 86494 20468 86546
rect 20412 85314 20468 86494
rect 20412 85262 20414 85314
rect 20466 85262 20468 85314
rect 20412 85250 20468 85262
rect 20636 86436 20692 86446
rect 20860 86436 20916 97412
rect 23436 96292 23492 96302
rect 23324 96290 23492 96292
rect 23324 96238 23438 96290
rect 23490 96238 23492 96290
rect 23324 96236 23492 96238
rect 21420 96066 21476 96078
rect 21420 96014 21422 96066
rect 21474 96014 21476 96066
rect 21420 95844 21476 96014
rect 22316 96066 22372 96078
rect 22316 96014 22318 96066
rect 22370 96014 22372 96066
rect 21420 95778 21476 95788
rect 22092 95844 22148 95854
rect 22148 95788 22260 95844
rect 22092 95778 22148 95788
rect 21196 95284 21252 95294
rect 21196 95190 21252 95228
rect 22204 95282 22260 95788
rect 22204 95230 22206 95282
rect 22258 95230 22260 95282
rect 22204 94610 22260 95230
rect 22316 95284 22372 96014
rect 22316 95218 22372 95228
rect 23324 95284 23380 96236
rect 23436 96226 23492 96236
rect 23548 95508 23604 99600
rect 26012 97468 26068 99600
rect 26012 97412 26404 97468
rect 25340 96180 25396 96190
rect 24220 95956 24276 95966
rect 25004 95956 25060 95966
rect 24220 95862 24276 95900
rect 24444 95954 25060 95956
rect 24444 95902 25006 95954
rect 25058 95902 25060 95954
rect 24444 95900 25060 95902
rect 23548 95442 23604 95452
rect 23884 95842 23940 95854
rect 23884 95790 23886 95842
rect 23938 95790 23940 95842
rect 22204 94558 22206 94610
rect 22258 94558 22260 94610
rect 22204 94546 22260 94558
rect 21532 94498 21588 94510
rect 21532 94446 21534 94498
rect 21586 94446 21588 94498
rect 21308 94274 21364 94286
rect 21308 94222 21310 94274
rect 21362 94222 21364 94274
rect 20972 93716 21028 93726
rect 21308 93716 21364 94222
rect 21532 93940 21588 94446
rect 22316 94500 22372 94510
rect 22652 94500 22708 94510
rect 22316 94498 22708 94500
rect 22316 94446 22318 94498
rect 22370 94446 22654 94498
rect 22706 94446 22708 94498
rect 22316 94444 22708 94446
rect 22316 94434 22372 94444
rect 22652 94434 22708 94444
rect 21980 94388 22036 94398
rect 21980 94294 22036 94332
rect 22764 94386 22820 94398
rect 22764 94334 22766 94386
rect 22818 94334 22820 94386
rect 22764 94276 22820 94334
rect 23212 94276 23268 94286
rect 22764 94274 23268 94276
rect 22764 94222 23214 94274
rect 23266 94222 23268 94274
rect 22764 94220 23268 94222
rect 21532 93874 21588 93884
rect 20972 93714 21364 93716
rect 20972 93662 20974 93714
rect 21026 93662 21364 93714
rect 20972 93660 21364 93662
rect 20972 93650 21028 93660
rect 20972 93044 21028 93054
rect 20972 92146 21028 92988
rect 21308 92930 21364 93660
rect 21308 92878 21310 92930
rect 21362 92878 21364 92930
rect 21308 92866 21364 92878
rect 21980 93714 22036 93726
rect 21980 93662 21982 93714
rect 22034 93662 22036 93714
rect 21980 92932 22036 93662
rect 23212 93380 23268 94220
rect 23212 93314 23268 93324
rect 23324 93938 23380 95228
rect 23548 95172 23604 95182
rect 23884 95172 23940 95790
rect 23548 95170 23940 95172
rect 23548 95118 23550 95170
rect 23602 95118 23940 95170
rect 23548 95116 23940 95118
rect 23548 95106 23604 95116
rect 23324 93886 23326 93938
rect 23378 93886 23380 93938
rect 23324 93156 23380 93886
rect 23436 93156 23492 93166
rect 23324 93154 23492 93156
rect 23324 93102 23438 93154
rect 23490 93102 23492 93154
rect 23324 93100 23492 93102
rect 22316 92932 22372 92942
rect 21980 92930 22372 92932
rect 21980 92878 22318 92930
rect 22370 92878 22372 92930
rect 21980 92876 22372 92878
rect 22204 92708 22260 92718
rect 20972 92094 20974 92146
rect 21026 92094 21028 92146
rect 20972 91924 21028 92094
rect 21644 92146 21700 92158
rect 21644 92094 21646 92146
rect 21698 92094 21700 92146
rect 21644 92036 21700 92094
rect 21644 91970 21700 91980
rect 20972 91858 21028 91868
rect 22204 91812 22260 92652
rect 22316 92372 22372 92876
rect 23212 92372 23268 92382
rect 22316 92370 23268 92372
rect 22316 92318 23214 92370
rect 23266 92318 23268 92370
rect 22316 92316 23268 92318
rect 23212 92306 23268 92316
rect 22316 92034 22372 92046
rect 23324 92036 23380 92046
rect 22316 91982 22318 92034
rect 22370 91982 22372 92034
rect 22316 91924 22372 91982
rect 23100 91980 23324 92036
rect 22428 91924 22484 91934
rect 22316 91868 22428 91924
rect 22428 91858 22484 91868
rect 22204 91756 22372 91812
rect 21756 90468 21812 90478
rect 21868 90468 21924 90478
rect 21756 90466 21868 90468
rect 21756 90414 21758 90466
rect 21810 90414 21868 90466
rect 21756 90412 21868 90414
rect 21756 90402 21812 90412
rect 21644 89908 21700 89918
rect 21644 89814 21700 89852
rect 21756 89572 21812 89582
rect 21196 89012 21252 89022
rect 21196 88898 21252 88956
rect 21196 88846 21198 88898
rect 21250 88846 21252 88898
rect 21196 88004 21252 88846
rect 21756 88450 21812 89516
rect 21868 89460 21924 90412
rect 22204 90466 22260 90478
rect 22204 90414 22206 90466
rect 22258 90414 22260 90466
rect 21868 89394 21924 89404
rect 21980 89908 22036 89918
rect 21980 89010 22036 89852
rect 22092 89684 22148 89694
rect 22092 89590 22148 89628
rect 21980 88958 21982 89010
rect 22034 88958 22036 89010
rect 21980 88946 22036 88958
rect 22092 89124 22148 89134
rect 21756 88398 21758 88450
rect 21810 88398 21812 88450
rect 21756 88386 21812 88398
rect 22092 88450 22148 89068
rect 22204 89012 22260 90414
rect 22204 88946 22260 88956
rect 22316 89796 22372 91756
rect 22988 90580 23044 90590
rect 22988 90486 23044 90524
rect 22652 90468 22708 90478
rect 22652 90466 22932 90468
rect 22652 90414 22654 90466
rect 22706 90414 22932 90466
rect 22652 90412 22932 90414
rect 22652 90402 22708 90412
rect 22764 89796 22820 89806
rect 22316 89794 22820 89796
rect 22316 89742 22766 89794
rect 22818 89742 22820 89794
rect 22316 89740 22820 89742
rect 22092 88398 22094 88450
rect 22146 88398 22148 88450
rect 22092 88386 22148 88398
rect 21532 88228 21588 88238
rect 21532 88134 21588 88172
rect 22204 88228 22260 88238
rect 21196 87938 21252 87948
rect 21196 87668 21252 87678
rect 21084 87556 21140 87566
rect 21084 87462 21140 87500
rect 20972 87444 21028 87454
rect 20972 87350 21028 87388
rect 21196 87442 21252 87612
rect 21196 87390 21198 87442
rect 21250 87390 21252 87442
rect 21196 87378 21252 87390
rect 22204 87442 22260 88172
rect 22204 87390 22206 87442
rect 22258 87390 22260 87442
rect 21980 86772 22036 86782
rect 21980 86658 22036 86716
rect 21980 86606 21982 86658
rect 22034 86606 22036 86658
rect 20636 86434 20916 86436
rect 20636 86382 20638 86434
rect 20690 86382 20916 86434
rect 20636 86380 20916 86382
rect 21084 86436 21140 86446
rect 20524 85092 20580 85102
rect 20300 85090 20580 85092
rect 20300 85038 20526 85090
rect 20578 85038 20580 85090
rect 20300 85036 20580 85038
rect 20188 85026 20244 85036
rect 20524 85026 20580 85036
rect 20132 84812 20244 84868
rect 20076 84802 20132 84812
rect 19836 84700 20100 84710
rect 19892 84644 19940 84700
rect 19996 84644 20044 84700
rect 19836 84634 20100 84644
rect 20188 84532 20244 84812
rect 20076 84476 20244 84532
rect 20412 84644 20468 84654
rect 19964 84420 20020 84430
rect 19964 84326 20020 84364
rect 19740 84084 19796 84094
rect 19628 84028 19740 84084
rect 19740 84018 19796 84028
rect 19852 84082 19908 84094
rect 19852 84030 19854 84082
rect 19906 84030 19908 84082
rect 19516 83524 19572 83534
rect 19516 83298 19572 83468
rect 19852 83412 19908 84030
rect 20076 83748 20132 84476
rect 20412 84418 20468 84588
rect 20636 84532 20692 86380
rect 20748 85876 20804 85886
rect 20748 85090 20804 85820
rect 20748 85038 20750 85090
rect 20802 85038 20804 85090
rect 20748 85026 20804 85038
rect 20412 84366 20414 84418
rect 20466 84366 20468 84418
rect 20412 84354 20468 84366
rect 20524 84476 20692 84532
rect 21084 84530 21140 86380
rect 21756 86212 21812 86222
rect 21756 85316 21812 86156
rect 21980 85764 22036 86606
rect 21980 85698 22036 85708
rect 22092 86770 22148 86782
rect 22092 86718 22094 86770
rect 22146 86718 22148 86770
rect 21084 84478 21086 84530
rect 21138 84478 21140 84530
rect 20188 84308 20244 84318
rect 20188 84306 20356 84308
rect 20188 84254 20190 84306
rect 20242 84254 20356 84306
rect 20188 84252 20356 84254
rect 20188 84242 20244 84252
rect 20076 83682 20132 83692
rect 19964 83636 20020 83646
rect 19964 83524 20020 83580
rect 19964 83522 20244 83524
rect 19964 83470 19966 83522
rect 20018 83470 20244 83522
rect 19964 83468 20244 83470
rect 19964 83458 20020 83468
rect 19516 83246 19518 83298
rect 19570 83246 19572 83298
rect 19516 83234 19572 83246
rect 19628 83356 19908 83412
rect 19628 82738 19684 83356
rect 19836 83132 20100 83142
rect 19892 83076 19940 83132
rect 19996 83076 20044 83132
rect 19836 83066 20100 83076
rect 19628 82686 19630 82738
rect 19682 82686 19684 82738
rect 19628 82674 19684 82686
rect 19404 82562 19460 82572
rect 20188 82068 20244 83468
rect 20300 83412 20356 84252
rect 20300 83346 20356 83356
rect 20412 83748 20468 83758
rect 20412 83634 20468 83692
rect 20412 83582 20414 83634
rect 20466 83582 20468 83634
rect 20412 83300 20468 83582
rect 20412 82516 20468 83244
rect 20524 82852 20580 84476
rect 21084 84466 21140 84478
rect 21308 85314 21812 85316
rect 21308 85262 21758 85314
rect 21810 85262 21812 85314
rect 21308 85260 21812 85262
rect 21308 84530 21364 85260
rect 21756 85250 21812 85260
rect 21420 85092 21476 85102
rect 21868 85092 21924 85102
rect 21476 85090 22036 85092
rect 21476 85038 21870 85090
rect 21922 85038 22036 85090
rect 21476 85036 22036 85038
rect 21420 84998 21476 85036
rect 21868 85026 21924 85036
rect 21308 84478 21310 84530
rect 21362 84478 21364 84530
rect 21308 84466 21364 84478
rect 20636 84308 20692 84318
rect 20636 84214 20692 84252
rect 20524 82786 20580 82796
rect 21196 84194 21252 84206
rect 21196 84142 21198 84194
rect 21250 84142 21252 84194
rect 20412 82450 20468 82460
rect 20972 82628 21028 82638
rect 20300 82068 20356 82078
rect 20188 82066 20356 82068
rect 20188 82014 20302 82066
rect 20354 82014 20356 82066
rect 20188 82012 20356 82014
rect 19836 81564 20100 81574
rect 19892 81508 19940 81564
rect 19996 81508 20044 81564
rect 19836 81498 20100 81508
rect 20188 81284 20244 82012
rect 20300 82002 20356 82012
rect 20188 80836 20244 81228
rect 20972 81282 21028 82572
rect 20972 81230 20974 81282
rect 21026 81230 21028 81282
rect 20972 81218 21028 81230
rect 21084 82516 21140 82526
rect 20860 81170 20916 81182
rect 20860 81118 20862 81170
rect 20914 81118 20916 81170
rect 20300 81060 20356 81070
rect 20636 81060 20692 81070
rect 20356 81058 20692 81060
rect 20356 81006 20638 81058
rect 20690 81006 20692 81058
rect 20356 81004 20692 81006
rect 20300 80966 20356 81004
rect 20636 80994 20692 81004
rect 20188 80780 20356 80836
rect 20076 80724 20132 80734
rect 20132 80668 20244 80724
rect 20076 80658 20132 80668
rect 19292 80558 19294 80610
rect 19346 80558 19348 80610
rect 19292 80546 19348 80558
rect 19404 80386 19460 80398
rect 19404 80334 19406 80386
rect 19458 80334 19460 80386
rect 19404 80164 19460 80334
rect 19404 80098 19460 80108
rect 20076 80386 20132 80398
rect 20076 80334 20078 80386
rect 20130 80334 20132 80386
rect 20076 80164 20132 80334
rect 20076 80098 20132 80108
rect 19836 79996 20100 80006
rect 19892 79940 19940 79996
rect 19996 79940 20044 79996
rect 19836 79930 20100 79940
rect 18396 78754 18452 78764
rect 18620 79324 18788 79380
rect 19068 79602 19124 79614
rect 19068 79550 19070 79602
rect 19122 79550 19124 79602
rect 18620 78260 18676 79324
rect 19068 78930 19124 79550
rect 19068 78878 19070 78930
rect 19122 78878 19124 78930
rect 19068 78866 19124 78878
rect 20076 78818 20132 78830
rect 20076 78766 20078 78818
rect 20130 78766 20132 78818
rect 19852 78596 19908 78606
rect 20076 78596 20132 78766
rect 19628 78594 20076 78596
rect 19628 78542 19854 78594
rect 19906 78542 20076 78594
rect 19628 78540 20076 78542
rect 18620 78166 18676 78204
rect 18732 78372 18788 78382
rect 18732 76466 18788 78316
rect 19628 78260 19684 78540
rect 19852 78530 19908 78540
rect 20076 78530 20132 78540
rect 19836 78428 20100 78438
rect 19892 78372 19940 78428
rect 19996 78372 20044 78428
rect 19836 78362 20100 78372
rect 19628 78194 19684 78204
rect 20188 78146 20244 80668
rect 20300 80610 20356 80780
rect 20300 80558 20302 80610
rect 20354 80558 20356 80610
rect 20300 80546 20356 80558
rect 20860 80500 20916 81118
rect 21084 81172 21140 82460
rect 21196 81956 21252 84142
rect 21868 83524 21924 83534
rect 21868 83430 21924 83468
rect 21980 83300 22036 85036
rect 21868 83244 22036 83300
rect 22092 85090 22148 86718
rect 22204 86772 22260 87390
rect 22204 86706 22260 86716
rect 22316 86770 22372 89740
rect 22764 89730 22820 89740
rect 22876 89684 22932 90412
rect 22540 89570 22596 89582
rect 22540 89518 22542 89570
rect 22594 89518 22596 89570
rect 22540 89460 22596 89518
rect 22540 89394 22596 89404
rect 22652 89570 22708 89582
rect 22652 89518 22654 89570
rect 22706 89518 22708 89570
rect 22428 88228 22484 88238
rect 22428 88134 22484 88172
rect 22652 87668 22708 89518
rect 22876 89236 22932 89628
rect 22876 89170 22932 89180
rect 22988 89570 23044 89582
rect 22988 89518 22990 89570
rect 23042 89518 23044 89570
rect 22764 88898 22820 88910
rect 22764 88846 22766 88898
rect 22818 88846 22820 88898
rect 22764 88452 22820 88846
rect 22764 88386 22820 88396
rect 22988 88900 23044 89518
rect 22988 87892 23044 88844
rect 22876 87836 23044 87892
rect 22316 86718 22318 86770
rect 22370 86718 22372 86770
rect 22316 86706 22372 86718
rect 22428 87612 22708 87668
rect 22764 87780 22820 87790
rect 22876 87780 22932 87836
rect 22820 87724 22932 87780
rect 22764 87666 22820 87724
rect 22764 87614 22766 87666
rect 22818 87614 22820 87666
rect 22428 85708 22484 87612
rect 22764 87602 22820 87614
rect 22988 87668 23044 87678
rect 23100 87668 23156 91980
rect 23324 91942 23380 91980
rect 23436 89908 23492 93100
rect 23548 90468 23604 90478
rect 23548 90374 23604 90412
rect 23436 89842 23492 89852
rect 23660 89796 23716 95116
rect 24332 94388 24388 94398
rect 24220 94386 24388 94388
rect 24220 94334 24334 94386
rect 24386 94334 24388 94386
rect 24220 94332 24388 94334
rect 24108 94274 24164 94286
rect 24108 94222 24110 94274
rect 24162 94222 24164 94274
rect 23884 93714 23940 93726
rect 23884 93662 23886 93714
rect 23938 93662 23940 93714
rect 23884 92484 23940 93662
rect 23884 92418 23940 92428
rect 23996 93604 24052 93614
rect 24108 93604 24164 94222
rect 23996 93602 24164 93604
rect 23996 93550 23998 93602
rect 24050 93550 24164 93602
rect 23996 93548 24164 93550
rect 23996 91924 24052 93548
rect 24108 93156 24164 93166
rect 24220 93156 24276 94332
rect 24332 94322 24388 94332
rect 24444 93492 24500 95900
rect 25004 95890 25060 95900
rect 25340 95954 25396 96124
rect 25340 95902 25342 95954
rect 25394 95902 25396 95954
rect 25340 95890 25396 95902
rect 25676 95844 25732 95854
rect 25452 95842 25732 95844
rect 25452 95790 25678 95842
rect 25730 95790 25732 95842
rect 25452 95788 25732 95790
rect 25452 95508 25508 95788
rect 25676 95778 25732 95788
rect 26012 95842 26068 95854
rect 26012 95790 26014 95842
rect 26066 95790 26068 95842
rect 26012 95732 26068 95790
rect 26012 95666 26068 95676
rect 25228 95452 25508 95508
rect 24668 95284 24724 95294
rect 24668 95190 24724 95228
rect 25004 94500 25060 94510
rect 24444 93426 24500 93436
rect 24556 94498 25060 94500
rect 24556 94446 25006 94498
rect 25058 94446 25060 94498
rect 24556 94444 25060 94446
rect 24556 93602 24612 94444
rect 25004 94434 25060 94444
rect 24668 94274 24724 94286
rect 24668 94222 24670 94274
rect 24722 94222 24724 94274
rect 24668 93716 24724 94222
rect 25228 93940 25284 95452
rect 25340 95282 25396 95294
rect 25340 95230 25342 95282
rect 25394 95230 25396 95282
rect 25340 94722 25396 95230
rect 26012 95284 26068 95294
rect 26068 95228 26292 95284
rect 26012 95190 26068 95228
rect 25340 94670 25342 94722
rect 25394 94670 25396 94722
rect 25340 94658 25396 94670
rect 26236 94612 26292 95228
rect 26236 94518 26292 94556
rect 25340 94500 25396 94510
rect 25676 94500 25732 94510
rect 25340 94498 25732 94500
rect 25340 94446 25342 94498
rect 25394 94446 25678 94498
rect 25730 94446 25732 94498
rect 25340 94444 25732 94446
rect 25340 94434 25396 94444
rect 25676 94434 25732 94444
rect 25788 94386 25844 94398
rect 25788 94334 25790 94386
rect 25842 94334 25844 94386
rect 25788 93940 25844 94334
rect 25228 93884 25508 93940
rect 25788 93884 26180 93940
rect 25228 93716 25284 93726
rect 24668 93714 25284 93716
rect 24668 93662 25230 93714
rect 25282 93662 25284 93714
rect 24668 93660 25284 93662
rect 25228 93650 25284 93660
rect 24556 93550 24558 93602
rect 24610 93550 24612 93602
rect 24108 93154 24276 93156
rect 24108 93102 24110 93154
rect 24162 93102 24276 93154
rect 24108 93100 24276 93102
rect 24444 93156 24500 93166
rect 24556 93156 24612 93550
rect 24444 93154 24612 93156
rect 24444 93102 24446 93154
rect 24498 93102 24612 93154
rect 24444 93100 24612 93102
rect 24668 93380 24724 93390
rect 24108 93090 24164 93100
rect 24444 93090 24500 93100
rect 24668 92930 24724 93324
rect 24668 92878 24670 92930
rect 24722 92878 24724 92930
rect 24668 92708 24724 92878
rect 25116 92708 25172 92718
rect 25228 92708 25284 92718
rect 24668 92706 25228 92708
rect 24668 92654 25118 92706
rect 25170 92654 25228 92706
rect 24668 92652 25228 92654
rect 25116 92642 25172 92652
rect 23996 91858 24052 91868
rect 24220 92034 24276 92046
rect 24220 91982 24222 92034
rect 24274 91982 24276 92034
rect 23548 89740 23716 89796
rect 23772 91250 23828 91262
rect 23772 91198 23774 91250
rect 23826 91198 23828 91250
rect 23324 89572 23380 89582
rect 23324 89478 23380 89516
rect 23436 89570 23492 89582
rect 23436 89518 23438 89570
rect 23490 89518 23492 89570
rect 22988 87666 23156 87668
rect 22988 87614 22990 87666
rect 23042 87614 23156 87666
rect 22988 87612 23156 87614
rect 23212 89460 23268 89470
rect 23212 87668 23268 89404
rect 23436 89012 23492 89518
rect 23548 89348 23604 89740
rect 23548 89282 23604 89292
rect 23660 89570 23716 89582
rect 23660 89518 23662 89570
rect 23714 89518 23716 89570
rect 23660 89236 23716 89518
rect 23660 89170 23716 89180
rect 23436 88946 23492 88956
rect 23548 89012 23604 89022
rect 23772 89012 23828 91198
rect 24108 90692 24164 90702
rect 24108 90598 24164 90636
rect 24220 89796 24276 91982
rect 24668 92034 24724 92046
rect 24668 91982 24670 92034
rect 24722 91982 24724 92034
rect 24668 91924 24724 91982
rect 24668 91858 24724 91868
rect 25116 90580 25172 90590
rect 25228 90580 25284 92652
rect 25340 92148 25396 92158
rect 25340 92054 25396 92092
rect 25452 90692 25508 93884
rect 26012 93716 26068 93726
rect 25676 93714 26068 93716
rect 25676 93662 26014 93714
rect 26066 93662 26068 93714
rect 25676 93660 26068 93662
rect 25676 93154 25732 93660
rect 26012 93650 26068 93660
rect 25676 93102 25678 93154
rect 25730 93102 25732 93154
rect 25676 93090 25732 93102
rect 25564 92818 25620 92830
rect 25564 92766 25566 92818
rect 25618 92766 25620 92818
rect 25564 92484 25620 92766
rect 26124 92708 26180 93884
rect 26124 92614 26180 92652
rect 26236 92820 26292 92830
rect 25564 92418 25620 92428
rect 26124 92260 26180 92298
rect 25900 92204 26124 92260
rect 25172 90524 25284 90580
rect 25340 90636 25508 90692
rect 25676 92148 25732 92158
rect 25116 90514 25172 90524
rect 24780 90468 24836 90478
rect 24780 90466 24948 90468
rect 24780 90414 24782 90466
rect 24834 90414 24948 90466
rect 24780 90412 24948 90414
rect 24780 90402 24836 90412
rect 23996 89740 24276 89796
rect 23548 89010 23828 89012
rect 23548 88958 23550 89010
rect 23602 88958 23828 89010
rect 23548 88956 23828 88958
rect 23884 89684 23940 89694
rect 23996 89684 24052 89740
rect 23884 89682 24052 89684
rect 23884 89630 23886 89682
rect 23938 89630 24052 89682
rect 23884 89628 24052 89630
rect 23548 88946 23604 88956
rect 23884 88564 23940 89628
rect 24220 89570 24276 89582
rect 24220 89518 24222 89570
rect 24274 89518 24276 89570
rect 24108 89348 24164 89358
rect 23996 89010 24052 89022
rect 23996 88958 23998 89010
rect 24050 88958 24052 89010
rect 23996 88900 24052 88958
rect 23996 88834 24052 88844
rect 23884 88498 23940 88508
rect 23884 88340 23940 88350
rect 24108 88340 24164 89292
rect 24220 89124 24276 89518
rect 24556 89572 24612 89582
rect 24556 89570 24836 89572
rect 24556 89518 24558 89570
rect 24610 89518 24836 89570
rect 24556 89516 24836 89518
rect 24556 89506 24612 89516
rect 24444 89460 24500 89470
rect 24444 89236 24500 89404
rect 24668 89236 24724 89246
rect 24444 89234 24724 89236
rect 24444 89182 24670 89234
rect 24722 89182 24724 89234
rect 24444 89180 24724 89182
rect 24668 89170 24724 89180
rect 24220 89058 24276 89068
rect 24780 89124 24836 89516
rect 24780 89058 24836 89068
rect 24892 89236 24948 90412
rect 24444 89012 24500 89022
rect 24444 88918 24500 88956
rect 23548 87668 23604 87678
rect 23212 87666 23604 87668
rect 23212 87614 23214 87666
rect 23266 87614 23550 87666
rect 23602 87614 23604 87666
rect 23212 87612 23604 87614
rect 22092 85038 22094 85090
rect 22146 85038 22148 85090
rect 22092 84194 22148 85038
rect 22092 84142 22094 84194
rect 22146 84142 22148 84194
rect 22092 83300 22148 84142
rect 21196 81890 21252 81900
rect 21420 83076 21476 83086
rect 21196 81172 21252 81182
rect 21084 81170 21252 81172
rect 21084 81118 21198 81170
rect 21250 81118 21252 81170
rect 21084 81116 21252 81118
rect 21196 81106 21252 81116
rect 21420 81170 21476 83020
rect 21420 81118 21422 81170
rect 21474 81118 21476 81170
rect 21420 81106 21476 81118
rect 21868 81172 21924 83244
rect 22092 83234 22148 83244
rect 22204 85652 22484 85708
rect 22652 86884 22708 86894
rect 21980 81284 22036 81294
rect 21980 81190 22036 81228
rect 21868 80612 21924 81116
rect 22092 81170 22148 81182
rect 22092 81118 22094 81170
rect 22146 81118 22148 81170
rect 22092 81060 22148 81118
rect 22092 80994 22148 81004
rect 21980 80948 22036 80958
rect 21980 80854 22036 80892
rect 21532 80556 21924 80612
rect 20860 80444 21028 80500
rect 20524 80388 20580 80398
rect 20188 78094 20190 78146
rect 20242 78094 20244 78146
rect 20188 78082 20244 78094
rect 20412 80332 20524 80388
rect 18732 76414 18734 76466
rect 18786 76414 18788 76466
rect 18732 76402 18788 76414
rect 19516 77252 19572 77262
rect 19292 76020 19348 76030
rect 19292 75908 19348 75964
rect 19516 75908 19572 77196
rect 19836 76860 20100 76870
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 19836 76794 20100 76804
rect 19292 75906 19572 75908
rect 19292 75854 19518 75906
rect 19570 75854 19572 75906
rect 19292 75852 19572 75854
rect 17836 73502 17838 73554
rect 17890 73502 17892 73554
rect 17836 73490 17892 73502
rect 17948 74898 18004 74910
rect 17948 74846 17950 74898
rect 18002 74846 18004 74898
rect 17948 74116 18004 74846
rect 18172 74898 18228 75068
rect 19068 75572 19124 75582
rect 18172 74846 18174 74898
rect 18226 74846 18228 74898
rect 18172 74834 18228 74846
rect 18508 74900 18564 74910
rect 19068 74900 19124 75516
rect 18508 74898 18900 74900
rect 18508 74846 18510 74898
rect 18562 74846 18900 74898
rect 18508 74844 18900 74846
rect 18508 74834 18564 74844
rect 18060 74788 18116 74798
rect 18060 74694 18116 74732
rect 18844 74338 18900 74844
rect 19068 74898 19236 74900
rect 19068 74846 19070 74898
rect 19122 74846 19236 74898
rect 19068 74844 19236 74846
rect 19068 74834 19124 74844
rect 18844 74286 18846 74338
rect 18898 74286 18900 74338
rect 18844 74274 18900 74286
rect 19068 74228 19124 74238
rect 19068 74134 19124 74172
rect 17948 73554 18004 74060
rect 17948 73502 17950 73554
rect 18002 73502 18004 73554
rect 17948 73490 18004 73502
rect 18844 73892 18900 73902
rect 18844 73554 18900 73836
rect 18844 73502 18846 73554
rect 18898 73502 18900 73554
rect 18844 73490 18900 73502
rect 16044 73390 16046 73442
rect 16098 73390 16100 73442
rect 16044 73378 16100 73390
rect 16828 73330 16884 73342
rect 16828 73278 16830 73330
rect 16882 73278 16884 73330
rect 16828 71764 16884 73278
rect 17724 73330 17780 73342
rect 17724 73278 17726 73330
rect 17778 73278 17780 73330
rect 17724 73220 17780 73278
rect 17724 73154 17780 73164
rect 18396 73220 18452 73230
rect 18396 73126 18452 73164
rect 18844 72212 18900 72222
rect 16828 71698 16884 71708
rect 17500 71764 17556 71774
rect 17500 71670 17556 71708
rect 18844 71762 18900 72156
rect 18844 71710 18846 71762
rect 18898 71710 18900 71762
rect 18844 71698 18900 71710
rect 19180 71764 19236 74844
rect 19180 71698 19236 71708
rect 17836 71092 17892 71102
rect 18284 71092 18340 71102
rect 17836 71090 18340 71092
rect 17836 71038 17838 71090
rect 17890 71038 18286 71090
rect 18338 71038 18340 71090
rect 17836 71036 18340 71038
rect 17836 71026 17892 71036
rect 18284 71026 18340 71036
rect 15708 70868 15764 70878
rect 15708 70866 15988 70868
rect 15708 70814 15710 70866
rect 15762 70814 15988 70866
rect 15708 70812 15988 70814
rect 15708 70802 15764 70812
rect 15484 70644 15540 70654
rect 15484 69076 15540 70588
rect 15932 70418 15988 70812
rect 15932 70366 15934 70418
rect 15986 70366 15988 70418
rect 15932 70354 15988 70366
rect 18396 70754 18452 70766
rect 18396 70702 18398 70754
rect 18450 70702 18452 70754
rect 15708 70308 15764 70318
rect 15708 70214 15764 70252
rect 16604 70308 16660 70318
rect 15596 70196 15652 70206
rect 15596 70102 15652 70140
rect 16268 70082 16324 70094
rect 16268 70030 16270 70082
rect 16322 70030 16324 70082
rect 16268 69524 16324 70030
rect 16268 69458 16324 69468
rect 15596 69300 15652 69310
rect 15596 69298 16324 69300
rect 15596 69246 15598 69298
rect 15650 69246 16324 69298
rect 15596 69244 16324 69246
rect 15596 69234 15652 69244
rect 15484 69020 15764 69076
rect 15372 68684 15652 68740
rect 15260 68674 15316 68684
rect 15372 68514 15428 68526
rect 15372 68462 15374 68514
rect 15426 68462 15428 68514
rect 15372 68404 15428 68462
rect 15372 68338 15428 68348
rect 15036 67060 15092 67070
rect 15036 66966 15092 67004
rect 15484 67060 15540 67070
rect 15484 66946 15540 67004
rect 15484 66894 15486 66946
rect 15538 66894 15540 66946
rect 14812 66334 14814 66386
rect 14866 66334 14868 66386
rect 14812 66322 14868 66334
rect 15260 66834 15316 66846
rect 15260 66782 15262 66834
rect 15314 66782 15316 66834
rect 15036 65490 15092 65502
rect 15036 65438 15038 65490
rect 15090 65438 15092 65490
rect 15036 64930 15092 65438
rect 15036 64878 15038 64930
rect 15090 64878 15092 64930
rect 15036 64866 15092 64878
rect 15036 64708 15092 64718
rect 15260 64708 15316 66782
rect 15484 66612 15540 66894
rect 15484 66546 15540 66556
rect 15596 66388 15652 68684
rect 15036 64706 15316 64708
rect 15036 64654 15038 64706
rect 15090 64654 15316 64706
rect 15036 64652 15316 64654
rect 15036 64642 15092 64652
rect 14924 64260 14980 64270
rect 14700 63868 14868 63924
rect 14252 63812 14308 63822
rect 14140 63810 14308 63812
rect 14140 63758 14254 63810
rect 14306 63758 14308 63810
rect 14140 63756 14308 63758
rect 14252 63746 14308 63756
rect 14028 63310 14030 63362
rect 14082 63310 14084 63362
rect 14028 63298 14084 63310
rect 13916 62738 13972 62748
rect 14252 62580 14308 62590
rect 13692 62578 14308 62580
rect 13692 62526 14254 62578
rect 14306 62526 14308 62578
rect 13692 62524 14308 62526
rect 14252 62514 14308 62524
rect 14364 62188 14420 63868
rect 14700 63700 14756 63710
rect 14588 63698 14756 63700
rect 14588 63646 14702 63698
rect 14754 63646 14756 63698
rect 14588 63644 14756 63646
rect 14476 63028 14532 63038
rect 14476 62934 14532 62972
rect 14028 62132 14420 62188
rect 14476 62692 14532 62702
rect 14028 61794 14084 62132
rect 14028 61742 14030 61794
rect 14082 61742 14084 61794
rect 14028 61730 14084 61742
rect 13916 61460 13972 61470
rect 13580 61394 13636 61404
rect 13804 61458 13972 61460
rect 13804 61406 13918 61458
rect 13970 61406 13972 61458
rect 13804 61404 13972 61406
rect 12460 60116 12516 60126
rect 12012 60114 12516 60116
rect 12012 60062 12462 60114
rect 12514 60062 12516 60114
rect 12012 60060 12516 60062
rect 12012 60002 12068 60060
rect 12460 60050 12516 60060
rect 12012 59950 12014 60002
rect 12066 59950 12068 60002
rect 12012 59938 12068 59950
rect 13468 60002 13524 60014
rect 13468 59950 13470 60002
rect 13522 59950 13524 60002
rect 13468 59220 13524 59950
rect 13524 59164 13636 59220
rect 13468 59154 13524 59164
rect 11676 59106 11732 59118
rect 11676 59054 11678 59106
rect 11730 59054 11732 59106
rect 11676 58436 11732 59054
rect 13468 58548 13524 58558
rect 11676 58380 12180 58436
rect 11676 58212 11732 58222
rect 11676 58118 11732 58156
rect 12124 57874 12180 58380
rect 12124 57822 12126 57874
rect 12178 57822 12180 57874
rect 12124 57810 12180 57822
rect 12460 57652 12516 57662
rect 12460 57558 12516 57596
rect 13020 56644 13076 56654
rect 12236 56084 12292 56094
rect 11564 55990 11620 56028
rect 12012 56028 12236 56084
rect 11452 54786 11508 54796
rect 11788 55970 11844 55982
rect 11788 55918 11790 55970
rect 11842 55918 11844 55970
rect 11676 54740 11732 54750
rect 11564 53508 11620 53518
rect 11452 53172 11508 53182
rect 11452 53078 11508 53116
rect 10892 50706 11396 50708
rect 10892 50654 11342 50706
rect 11394 50654 11396 50706
rect 10892 50652 11396 50654
rect 10892 50594 10948 50652
rect 11340 50642 11396 50652
rect 10892 50542 10894 50594
rect 10946 50542 10948 50594
rect 10892 50530 10948 50542
rect 10556 50372 10612 50382
rect 10780 50372 10948 50428
rect 10556 50370 10724 50372
rect 10556 50318 10558 50370
rect 10610 50318 10724 50370
rect 10556 50316 10724 50318
rect 10556 50306 10612 50316
rect 10444 49980 10612 50036
rect 10108 49970 10164 49980
rect 10220 49922 10276 49934
rect 10220 49870 10222 49922
rect 10274 49870 10276 49922
rect 10220 49588 10276 49870
rect 10444 49812 10500 49822
rect 10444 49718 10500 49756
rect 10220 49532 10500 49588
rect 10332 49364 10388 49374
rect 9660 48466 9716 48524
rect 9660 48414 9662 48466
rect 9714 48414 9716 48466
rect 9660 48402 9716 48414
rect 10108 49028 10164 49038
rect 9996 48242 10052 48254
rect 9996 48190 9998 48242
rect 10050 48190 10052 48242
rect 9996 48132 10052 48190
rect 9996 48066 10052 48076
rect 8988 47518 8990 47570
rect 9042 47518 9044 47570
rect 8988 47506 9044 47518
rect 9436 47460 9492 47470
rect 8316 47236 8372 47246
rect 8316 44884 8372 47180
rect 9436 46564 9492 47404
rect 10108 47460 10164 48972
rect 10108 47366 10164 47404
rect 10220 48580 10276 48590
rect 10220 48466 10276 48524
rect 10220 48414 10222 48466
rect 10274 48414 10276 48466
rect 9660 46564 9716 46574
rect 9436 46562 9716 46564
rect 9436 46510 9662 46562
rect 9714 46510 9716 46562
rect 9436 46508 9716 46510
rect 8540 44996 8596 45006
rect 8540 44994 9044 44996
rect 8540 44942 8542 44994
rect 8594 44942 9044 44994
rect 8540 44940 9044 44942
rect 8540 44930 8596 44940
rect 8316 44790 8372 44828
rect 8204 44492 8372 44548
rect 8092 44380 8260 44436
rect 8092 41972 8148 41982
rect 8092 41878 8148 41916
rect 7980 39396 8036 39406
rect 7980 31892 8036 39340
rect 8092 32676 8148 32686
rect 8092 32582 8148 32620
rect 7980 31836 8148 31892
rect 7980 31666 8036 31678
rect 7980 31614 7982 31666
rect 8034 31614 8036 31666
rect 7980 31218 8036 31614
rect 7980 31166 7982 31218
rect 8034 31166 8036 31218
rect 7980 31154 8036 31166
rect 8092 30212 8148 31836
rect 8092 30146 8148 30156
rect 8204 29988 8260 44380
rect 7980 29932 8260 29988
rect 7980 28756 8036 29932
rect 7980 28690 8036 28700
rect 8204 28756 8260 28766
rect 8204 28642 8260 28700
rect 8204 28590 8206 28642
rect 8258 28590 8260 28642
rect 8204 28578 8260 28590
rect 8316 28644 8372 44492
rect 8988 43428 9044 44940
rect 8988 43334 9044 43372
rect 9660 43426 9716 46508
rect 10220 44548 10276 48414
rect 10332 48466 10388 49308
rect 10444 49138 10500 49532
rect 10444 49086 10446 49138
rect 10498 49086 10500 49138
rect 10444 49074 10500 49086
rect 10332 48414 10334 48466
rect 10386 48414 10388 48466
rect 10332 48402 10388 48414
rect 10444 48692 10500 48702
rect 10444 48466 10500 48636
rect 10444 48414 10446 48466
rect 10498 48414 10500 48466
rect 10444 48402 10500 48414
rect 10220 44492 10388 44548
rect 9660 43374 9662 43426
rect 9714 43374 9716 43426
rect 9660 43316 9716 43374
rect 10108 43426 10164 43438
rect 10108 43374 10110 43426
rect 10162 43374 10164 43426
rect 10108 43316 10164 43374
rect 9660 43260 10164 43316
rect 10220 43428 10276 43438
rect 9436 42866 9492 42878
rect 9436 42814 9438 42866
rect 9490 42814 9492 42866
rect 9324 42532 9380 42542
rect 9324 38668 9380 42476
rect 9436 42084 9492 42814
rect 9884 42756 9940 43260
rect 9772 42642 9828 42654
rect 9772 42590 9774 42642
rect 9826 42590 9828 42642
rect 9548 42084 9604 42094
rect 9772 42084 9828 42590
rect 9436 42082 9828 42084
rect 9436 42030 9550 42082
rect 9602 42030 9828 42082
rect 9436 42028 9828 42030
rect 9548 42018 9604 42028
rect 9772 41860 9828 41870
rect 9772 41766 9828 41804
rect 9884 41188 9940 42700
rect 10220 42754 10276 43372
rect 10220 42702 10222 42754
rect 10274 42702 10276 42754
rect 10220 42690 10276 42702
rect 10332 42756 10388 44492
rect 10556 44324 10612 49980
rect 10668 49924 10724 50316
rect 10668 49868 10836 49924
rect 10668 48242 10724 48254
rect 10668 48190 10670 48242
rect 10722 48190 10724 48242
rect 10668 48132 10724 48190
rect 10668 48066 10724 48076
rect 10780 47572 10836 49868
rect 10556 44258 10612 44268
rect 10668 47516 10836 47572
rect 9996 42644 10052 42654
rect 9996 42084 10052 42588
rect 10108 42532 10164 42542
rect 10108 42438 10164 42476
rect 9996 42018 10052 42028
rect 10332 42084 10388 42700
rect 10332 42018 10388 42028
rect 10556 41970 10612 41982
rect 10556 41918 10558 41970
rect 10610 41918 10612 41970
rect 10108 41860 10164 41870
rect 10556 41860 10612 41918
rect 10108 41858 10612 41860
rect 10108 41806 10110 41858
rect 10162 41806 10612 41858
rect 10108 41804 10612 41806
rect 10108 41794 10164 41804
rect 10668 41748 10724 47516
rect 10780 47346 10836 47358
rect 10780 47294 10782 47346
rect 10834 47294 10836 47346
rect 10780 46898 10836 47294
rect 10780 46846 10782 46898
rect 10834 46846 10836 46898
rect 10780 46834 10836 46846
rect 10892 42308 10948 50372
rect 11116 50036 11172 50046
rect 11116 49942 11172 49980
rect 11004 49812 11060 49822
rect 11060 49756 11172 49812
rect 11004 49746 11060 49756
rect 11116 48804 11172 49756
rect 11564 49140 11620 53452
rect 11676 50036 11732 54684
rect 11788 53732 11844 55918
rect 11788 53666 11844 53676
rect 11900 55412 11956 55422
rect 11900 54404 11956 55356
rect 11788 52834 11844 52846
rect 11788 52782 11790 52834
rect 11842 52782 11844 52834
rect 11788 52276 11844 52782
rect 11788 52210 11844 52220
rect 11900 50428 11956 54348
rect 12012 53172 12068 56028
rect 12236 55990 12292 56028
rect 12236 55074 12292 55086
rect 12236 55022 12238 55074
rect 12290 55022 12292 55074
rect 12236 53956 12292 55022
rect 12684 55074 12740 55086
rect 12684 55022 12686 55074
rect 12738 55022 12740 55074
rect 12684 54740 12740 55022
rect 12684 54674 12740 54684
rect 13020 54626 13076 56588
rect 13020 54574 13022 54626
rect 13074 54574 13076 54626
rect 13020 54562 13076 54574
rect 12348 54514 12404 54526
rect 12348 54462 12350 54514
rect 12402 54462 12404 54514
rect 12348 54068 12404 54462
rect 13468 54068 13524 58492
rect 13580 58548 13636 59164
rect 13804 59106 13860 61404
rect 13916 61394 13972 61404
rect 14364 61348 14420 61358
rect 14252 61346 14420 61348
rect 14252 61294 14366 61346
rect 14418 61294 14420 61346
rect 14252 61292 14420 61294
rect 14252 60114 14308 61292
rect 14364 61282 14420 61292
rect 14252 60062 14254 60114
rect 14306 60062 14308 60114
rect 14252 60050 14308 60062
rect 14476 59668 14532 62636
rect 14588 62356 14644 63644
rect 14700 63634 14756 63644
rect 14812 62916 14868 63868
rect 14812 62850 14868 62860
rect 14700 62580 14756 62590
rect 14924 62580 14980 64204
rect 15148 63922 15204 63934
rect 15148 63870 15150 63922
rect 15202 63870 15204 63922
rect 15148 63362 15204 63870
rect 15148 63310 15150 63362
rect 15202 63310 15204 63362
rect 15148 63298 15204 63310
rect 15036 63140 15092 63150
rect 15260 63140 15316 64652
rect 15036 63138 15316 63140
rect 15036 63086 15038 63138
rect 15090 63086 15316 63138
rect 15036 63084 15316 63086
rect 15036 63074 15092 63084
rect 14700 62578 14980 62580
rect 14700 62526 14702 62578
rect 14754 62526 14980 62578
rect 14700 62524 14980 62526
rect 15036 62916 15092 62926
rect 14700 62514 14756 62524
rect 14588 61458 14644 62300
rect 14588 61406 14590 61458
rect 14642 61406 14644 61458
rect 14588 61394 14644 61406
rect 14700 61460 14756 61470
rect 13804 59054 13806 59106
rect 13858 59054 13860 59106
rect 13804 59042 13860 59054
rect 14252 59612 14532 59668
rect 14252 59442 14308 59612
rect 14700 59556 14756 61404
rect 14252 59390 14254 59442
rect 14306 59390 14308 59442
rect 14252 59108 14308 59390
rect 14252 59042 14308 59052
rect 14364 59500 14756 59556
rect 14364 58884 14420 59500
rect 14252 58828 14420 58884
rect 14476 59332 14532 59342
rect 13804 58660 13860 58670
rect 13804 58548 13860 58604
rect 13580 58546 13860 58548
rect 13580 58494 13582 58546
rect 13634 58494 13860 58546
rect 13580 58492 13860 58494
rect 13580 58482 13636 58492
rect 13804 58212 13860 58492
rect 14028 58436 14084 58446
rect 14028 58342 14084 58380
rect 13804 58156 14196 58212
rect 14140 57762 14196 58156
rect 14140 57710 14142 57762
rect 14194 57710 14196 57762
rect 14140 57698 14196 57710
rect 13692 57652 13748 57662
rect 13468 54012 13636 54068
rect 12348 54002 12404 54012
rect 12236 53890 12292 53900
rect 12908 53842 12964 53854
rect 12908 53790 12910 53842
rect 12962 53790 12964 53842
rect 12908 53732 12964 53790
rect 12012 52946 12068 53116
rect 12348 53620 12404 53630
rect 12348 53170 12404 53564
rect 12348 53118 12350 53170
rect 12402 53118 12404 53170
rect 12348 53106 12404 53118
rect 12012 52894 12014 52946
rect 12066 52894 12068 52946
rect 12012 51268 12068 52894
rect 12908 52612 12964 53676
rect 13468 53844 13524 53854
rect 13468 53618 13524 53788
rect 13468 53566 13470 53618
rect 13522 53566 13524 53618
rect 13468 53554 13524 53566
rect 13020 52836 13076 52846
rect 13020 52742 13076 52780
rect 12908 52556 13076 52612
rect 12908 52276 12964 52286
rect 12908 52182 12964 52220
rect 13020 52164 13076 52556
rect 13020 52098 13076 52108
rect 12012 51202 12068 51212
rect 13580 50428 13636 54012
rect 11676 49970 11732 49980
rect 11788 50372 11956 50428
rect 13468 50372 13636 50428
rect 11676 49812 11732 49822
rect 11676 49718 11732 49756
rect 11676 49140 11732 49150
rect 11228 49138 11732 49140
rect 11228 49086 11678 49138
rect 11730 49086 11732 49138
rect 11228 49084 11732 49086
rect 11228 49028 11284 49084
rect 11676 49074 11732 49084
rect 11228 48934 11284 48972
rect 11116 48748 11396 48804
rect 11340 48466 11396 48748
rect 11340 48414 11342 48466
rect 11394 48414 11396 48466
rect 11340 48402 11396 48414
rect 11452 48692 11508 48702
rect 11004 46900 11060 46910
rect 11228 46900 11284 46910
rect 11004 46898 11284 46900
rect 11004 46846 11006 46898
rect 11058 46846 11230 46898
rect 11282 46846 11284 46898
rect 11004 46844 11284 46846
rect 11452 46900 11508 48636
rect 11676 48020 11732 48030
rect 11564 46900 11620 46910
rect 11452 46844 11564 46900
rect 11004 46834 11060 46844
rect 11228 46834 11284 46844
rect 11564 46834 11620 46844
rect 11452 46674 11508 46686
rect 11452 46622 11454 46674
rect 11506 46622 11508 46674
rect 11340 45332 11396 45342
rect 11452 45332 11508 46622
rect 11340 45330 11508 45332
rect 11340 45278 11342 45330
rect 11394 45278 11508 45330
rect 11340 45276 11508 45278
rect 11340 45266 11396 45276
rect 11004 44996 11060 45006
rect 11676 44996 11732 47964
rect 11004 44994 11732 44996
rect 11004 44942 11006 44994
rect 11058 44942 11678 44994
rect 11730 44942 11732 44994
rect 11004 44940 11732 44942
rect 11004 44930 11060 44940
rect 11004 42532 11060 42542
rect 11004 42438 11060 42476
rect 10892 42252 11060 42308
rect 10332 41692 10724 41748
rect 10892 42082 10948 42094
rect 10892 42030 10894 42082
rect 10946 42030 10948 42082
rect 9996 41188 10052 41198
rect 9884 41186 10052 41188
rect 9884 41134 9998 41186
rect 10050 41134 10052 41186
rect 9884 41132 10052 41134
rect 9996 40628 10052 41132
rect 9996 40402 10052 40572
rect 9996 40350 9998 40402
rect 10050 40350 10052 40402
rect 9996 40338 10052 40350
rect 10108 38834 10164 38846
rect 10108 38782 10110 38834
rect 10162 38782 10164 38834
rect 9324 38612 9492 38668
rect 8540 36596 8596 36606
rect 8540 36502 8596 36540
rect 9100 36596 9156 36606
rect 8988 36482 9044 36494
rect 8988 36430 8990 36482
rect 9042 36430 9044 36482
rect 8988 35924 9044 36430
rect 9100 36482 9156 36540
rect 9100 36430 9102 36482
rect 9154 36430 9156 36482
rect 9100 36418 9156 36430
rect 9436 36482 9492 38612
rect 9548 37940 9604 37950
rect 9548 37846 9604 37884
rect 9772 37828 9828 37838
rect 9772 37266 9828 37772
rect 10108 37490 10164 38782
rect 10108 37438 10110 37490
rect 10162 37438 10164 37490
rect 10108 37426 10164 37438
rect 10220 38052 10276 38062
rect 9772 37214 9774 37266
rect 9826 37214 9828 37266
rect 9772 37202 9828 37214
rect 9436 36430 9438 36482
rect 9490 36430 9492 36482
rect 9436 36418 9492 36430
rect 9548 37154 9604 37166
rect 9548 37102 9550 37154
rect 9602 37102 9604 37154
rect 9212 36370 9268 36382
rect 9212 36318 9214 36370
rect 9266 36318 9268 36370
rect 9100 35924 9156 35934
rect 8988 35868 9100 35924
rect 9100 35858 9156 35868
rect 9212 31668 9268 36318
rect 9548 35812 9604 37102
rect 10220 37156 10276 37996
rect 9772 36484 9828 36494
rect 9772 35922 9828 36428
rect 9884 36260 9940 36270
rect 9884 36166 9940 36204
rect 9772 35870 9774 35922
rect 9826 35870 9828 35922
rect 9772 35858 9828 35870
rect 9884 35924 9940 35934
rect 9884 35830 9940 35868
rect 9548 35810 9716 35812
rect 9548 35758 9550 35810
rect 9602 35758 9716 35810
rect 9548 35756 9716 35758
rect 9548 35746 9604 35756
rect 9660 35026 9716 35756
rect 9996 35698 10052 35710
rect 9996 35646 9998 35698
rect 10050 35646 10052 35698
rect 9996 35140 10052 35646
rect 10108 35700 10164 35710
rect 10108 35606 10164 35644
rect 9660 34974 9662 35026
rect 9714 34974 9716 35026
rect 9660 34962 9716 34974
rect 9884 35084 10052 35140
rect 9884 34244 9940 35084
rect 10108 34916 10164 34926
rect 10220 34916 10276 37100
rect 10108 34914 10276 34916
rect 10108 34862 10110 34914
rect 10162 34862 10276 34914
rect 10108 34860 10276 34862
rect 9884 34188 10052 34244
rect 9884 34020 9940 34030
rect 9884 33926 9940 33964
rect 8652 31612 9268 31668
rect 9324 31892 9380 31902
rect 9996 31892 10052 34188
rect 10108 34020 10164 34860
rect 10108 33954 10164 33964
rect 10108 31892 10164 31902
rect 8316 28588 8484 28644
rect 7980 28532 8036 28542
rect 7980 28530 8148 28532
rect 7980 28478 7982 28530
rect 8034 28478 8148 28530
rect 7980 28476 8148 28478
rect 7980 28466 8036 28476
rect 7980 28308 8036 28318
rect 7980 18004 8036 28252
rect 8092 27972 8148 28476
rect 8428 28308 8484 28588
rect 8316 28252 8484 28308
rect 8204 27972 8260 27982
rect 8092 27970 8260 27972
rect 8092 27918 8206 27970
rect 8258 27918 8260 27970
rect 8092 27916 8260 27918
rect 8204 27906 8260 27916
rect 8316 27748 8372 28252
rect 8204 27692 8372 27748
rect 8092 27636 8148 27646
rect 8092 26290 8148 27580
rect 8092 26238 8094 26290
rect 8146 26238 8148 26290
rect 8092 26226 8148 26238
rect 8204 21140 8260 27692
rect 8428 26962 8484 26974
rect 8428 26910 8430 26962
rect 8482 26910 8484 26962
rect 8428 26908 8484 26910
rect 8316 26852 8484 26908
rect 8316 26514 8372 26852
rect 8316 26462 8318 26514
rect 8370 26462 8372 26514
rect 8316 26450 8372 26462
rect 8428 23604 8484 23614
rect 8316 23548 8428 23604
rect 8316 23154 8372 23548
rect 8428 23538 8484 23548
rect 8652 23378 8708 31612
rect 8988 31220 9044 31230
rect 8988 31126 9044 31164
rect 9212 28756 9268 28766
rect 9324 28756 9380 31836
rect 9884 31890 10164 31892
rect 9884 31838 10110 31890
rect 10162 31838 10164 31890
rect 9884 31836 10164 31838
rect 9884 30994 9940 31836
rect 10108 31826 10164 31836
rect 9884 30942 9886 30994
rect 9938 30942 9940 30994
rect 9884 30930 9940 30942
rect 10108 31220 10164 31230
rect 10108 30994 10164 31164
rect 10108 30942 10110 30994
rect 10162 30942 10164 30994
rect 10108 30772 10164 30942
rect 10108 30706 10164 30716
rect 9884 29652 9940 29662
rect 9884 29558 9940 29596
rect 8988 28754 9380 28756
rect 8988 28702 9214 28754
rect 9266 28702 9380 28754
rect 8988 28700 9380 28702
rect 10220 29202 10276 29214
rect 10220 29150 10222 29202
rect 10274 29150 10276 29202
rect 8988 27858 9044 28700
rect 9212 28690 9268 28700
rect 10108 28644 10164 28654
rect 10108 28550 10164 28588
rect 8988 27806 8990 27858
rect 9042 27806 9044 27858
rect 8988 27076 9044 27806
rect 9884 27860 9940 27870
rect 9884 27766 9940 27804
rect 10108 27748 10164 27758
rect 10108 27654 10164 27692
rect 9548 27636 9604 27646
rect 9548 27542 9604 27580
rect 9100 27076 9156 27086
rect 9660 27076 9716 27086
rect 8988 27074 9716 27076
rect 8988 27022 9102 27074
rect 9154 27022 9662 27074
rect 9714 27022 9716 27074
rect 8988 27020 9716 27022
rect 9100 27010 9156 27020
rect 9660 24722 9716 27020
rect 9660 24670 9662 24722
rect 9714 24670 9716 24722
rect 9660 24658 9716 24670
rect 9996 24612 10052 24622
rect 9772 23940 9828 23950
rect 9772 23938 9940 23940
rect 9772 23886 9774 23938
rect 9826 23886 9940 23938
rect 9772 23884 9940 23886
rect 9772 23874 9828 23884
rect 9212 23714 9268 23726
rect 9212 23662 9214 23714
rect 9266 23662 9268 23714
rect 9212 23604 9268 23662
rect 9212 23538 9268 23548
rect 9884 23492 9940 23884
rect 9996 23826 10052 24556
rect 9996 23774 9998 23826
rect 10050 23774 10052 23826
rect 9996 23762 10052 23774
rect 9884 23436 10164 23492
rect 8652 23326 8654 23378
rect 8706 23326 8708 23378
rect 8652 23314 8708 23326
rect 9772 23380 9828 23390
rect 8316 23102 8318 23154
rect 8370 23102 8372 23154
rect 8316 23090 8372 23102
rect 8540 23154 8596 23166
rect 8540 23102 8542 23154
rect 8594 23102 8596 23154
rect 8540 22596 8596 23102
rect 8764 23156 8820 23166
rect 8764 23062 8820 23100
rect 8876 23154 8932 23166
rect 8876 23102 8878 23154
rect 8930 23102 8932 23154
rect 8876 23044 8932 23102
rect 9772 23154 9828 23324
rect 10108 23378 10164 23436
rect 10108 23326 10110 23378
rect 10162 23326 10164 23378
rect 10108 23314 10164 23326
rect 9772 23102 9774 23154
rect 9826 23102 9828 23154
rect 9772 23090 9828 23102
rect 9548 23044 9604 23054
rect 8876 23042 9604 23044
rect 8876 22990 9550 23042
rect 9602 22990 9604 23042
rect 8876 22988 9604 22990
rect 8204 21074 8260 21084
rect 8428 22540 8596 22596
rect 8652 22596 8708 22606
rect 8428 20802 8484 22540
rect 8652 22370 8708 22540
rect 8652 22318 8654 22370
rect 8706 22318 8708 22370
rect 8652 22306 8708 22318
rect 8876 21474 8932 22988
rect 9548 22978 9604 22988
rect 10220 22708 10276 29150
rect 10332 26908 10388 41692
rect 10780 41300 10836 41310
rect 10892 41300 10948 42030
rect 10780 41298 10948 41300
rect 10780 41246 10782 41298
rect 10834 41246 10948 41298
rect 10780 41244 10948 41246
rect 10780 41234 10836 41244
rect 10668 40292 10724 40302
rect 10444 40290 10724 40292
rect 10444 40238 10670 40290
rect 10722 40238 10724 40290
rect 10444 40236 10724 40238
rect 10444 39058 10500 40236
rect 10668 40226 10724 40236
rect 10444 39006 10446 39058
rect 10498 39006 10500 39058
rect 10444 38994 10500 39006
rect 11004 38668 11060 42252
rect 10892 38612 11060 38668
rect 10668 37940 10724 37950
rect 10668 37846 10724 37884
rect 10556 37828 10612 37838
rect 10556 37490 10612 37772
rect 10556 37438 10558 37490
rect 10610 37438 10612 37490
rect 10556 37426 10612 37438
rect 10668 36484 10724 36494
rect 10668 35922 10724 36428
rect 10668 35870 10670 35922
rect 10722 35870 10724 35922
rect 10668 35858 10724 35870
rect 10780 35474 10836 35486
rect 10780 35422 10782 35474
rect 10834 35422 10836 35474
rect 10780 35026 10836 35422
rect 10780 34974 10782 35026
rect 10834 34974 10836 35026
rect 10780 34962 10836 34974
rect 10556 34020 10612 34030
rect 10556 31892 10612 33964
rect 10556 31798 10612 31836
rect 10444 30772 10500 30782
rect 10444 30770 10724 30772
rect 10444 30718 10446 30770
rect 10498 30718 10724 30770
rect 10444 30716 10724 30718
rect 10444 30706 10500 30716
rect 10556 30212 10612 30222
rect 10556 29652 10612 30156
rect 10668 30210 10724 30716
rect 10668 30158 10670 30210
rect 10722 30158 10724 30210
rect 10668 30146 10724 30158
rect 10892 30100 10948 38612
rect 11004 37940 11060 37950
rect 11004 37846 11060 37884
rect 11116 35924 11172 44940
rect 11676 44930 11732 44940
rect 11452 43540 11508 43550
rect 11452 43538 11620 43540
rect 11452 43486 11454 43538
rect 11506 43486 11620 43538
rect 11452 43484 11620 43486
rect 11452 43474 11508 43484
rect 11228 42756 11284 42766
rect 11284 42700 11396 42756
rect 11228 42690 11284 42700
rect 11340 42642 11396 42700
rect 11340 42590 11342 42642
rect 11394 42590 11396 42642
rect 11340 42578 11396 42590
rect 11452 42532 11508 42542
rect 11340 41860 11396 41870
rect 11340 41766 11396 41804
rect 11452 39620 11508 42476
rect 11564 41972 11620 43484
rect 11676 41972 11732 41982
rect 11564 41916 11676 41972
rect 11676 41906 11732 41916
rect 11452 39554 11508 39564
rect 11788 38668 11844 50372
rect 12348 49700 12404 49710
rect 12348 49606 12404 49644
rect 12460 49252 12516 49262
rect 12460 49138 12516 49196
rect 13468 49252 13524 50372
rect 13468 49158 13524 49196
rect 13580 49700 13636 49710
rect 12460 49086 12462 49138
rect 12514 49086 12516 49138
rect 12460 49074 12516 49086
rect 13580 49138 13636 49644
rect 13580 49086 13582 49138
rect 13634 49086 13636 49138
rect 13580 49074 13636 49086
rect 13020 48916 13076 48926
rect 13692 48916 13748 57596
rect 14140 56642 14196 56654
rect 14140 56590 14142 56642
rect 14194 56590 14196 56642
rect 14140 56420 14196 56590
rect 14252 56420 14308 58828
rect 14476 58772 14532 59276
rect 14588 59220 14644 59230
rect 15036 59220 15092 62860
rect 15260 62692 15316 63084
rect 15484 66386 15652 66388
rect 15484 66334 15598 66386
rect 15650 66334 15652 66386
rect 15484 66332 15652 66334
rect 15484 64706 15540 66332
rect 15596 66322 15652 66332
rect 15596 65492 15652 65502
rect 15596 65398 15652 65436
rect 15708 65156 15764 69020
rect 15820 68852 15876 68862
rect 15820 68758 15876 68796
rect 16268 68850 16324 69244
rect 16268 68798 16270 68850
rect 16322 68798 16324 68850
rect 16268 68786 16324 68798
rect 16380 68738 16436 68750
rect 16380 68686 16382 68738
rect 16434 68686 16436 68738
rect 16156 68404 16212 68414
rect 16156 67732 16212 68348
rect 16156 67666 16212 67676
rect 16044 66946 16100 66958
rect 16044 66894 16046 66946
rect 16098 66894 16100 66946
rect 16044 65380 16100 66894
rect 16380 66164 16436 68686
rect 16492 66946 16548 66958
rect 16492 66894 16494 66946
rect 16546 66894 16548 66946
rect 16492 66834 16548 66894
rect 16492 66782 16494 66834
rect 16546 66782 16548 66834
rect 16492 66770 16548 66782
rect 16604 66386 16660 70252
rect 18396 70308 18452 70702
rect 18844 70754 18900 70766
rect 18844 70702 18846 70754
rect 18898 70702 18900 70754
rect 18396 70306 18788 70308
rect 18396 70254 18398 70306
rect 18450 70254 18788 70306
rect 18396 70252 18788 70254
rect 18396 70242 18452 70252
rect 17836 70084 17892 70094
rect 18172 70084 18228 70094
rect 17612 70082 18228 70084
rect 17612 70030 17838 70082
rect 17890 70030 18174 70082
rect 18226 70030 18228 70082
rect 17612 70028 18228 70030
rect 16940 68852 16996 68862
rect 16828 67732 16884 67742
rect 16828 67638 16884 67676
rect 16940 67172 16996 68796
rect 17500 68852 17556 68862
rect 17500 68626 17556 68796
rect 17500 68574 17502 68626
rect 17554 68574 17556 68626
rect 17500 68562 17556 68574
rect 17612 67732 17668 70028
rect 17836 70018 17892 70028
rect 18172 70018 18228 70028
rect 18508 70084 18564 70094
rect 18508 69990 18564 70028
rect 17724 69524 17780 69534
rect 18172 69524 18228 69534
rect 17724 69522 18228 69524
rect 17724 69470 17726 69522
rect 17778 69470 18174 69522
rect 18226 69470 18228 69522
rect 17724 69468 18228 69470
rect 17724 69458 17780 69468
rect 18172 69458 18228 69468
rect 18060 69188 18116 69198
rect 17836 69186 18116 69188
rect 17836 69134 18062 69186
rect 18114 69134 18116 69186
rect 17836 69132 18116 69134
rect 17836 67732 17892 69132
rect 18060 69122 18116 69132
rect 18172 68516 18228 68526
rect 17948 68514 18228 68516
rect 17948 68462 18174 68514
rect 18226 68462 18228 68514
rect 17948 68460 18228 68462
rect 17948 68066 18004 68460
rect 18172 68450 18228 68460
rect 17948 68014 17950 68066
rect 18002 68014 18004 68066
rect 17948 68002 18004 68014
rect 17612 67638 17668 67676
rect 17724 67730 17892 67732
rect 17724 67678 17838 67730
rect 17890 67678 17892 67730
rect 17724 67676 17892 67678
rect 16604 66334 16606 66386
rect 16658 66334 16660 66386
rect 16604 66322 16660 66334
rect 16828 67116 16996 67172
rect 17388 67618 17444 67630
rect 17388 67566 17390 67618
rect 17442 67566 17444 67618
rect 16492 66276 16548 66286
rect 16492 66182 16548 66220
rect 16380 66098 16436 66108
rect 16268 65604 16324 65614
rect 16268 65510 16324 65548
rect 16716 65380 16772 65390
rect 16044 65378 16772 65380
rect 16044 65326 16046 65378
rect 16098 65326 16718 65378
rect 16770 65326 16772 65378
rect 16044 65324 16772 65326
rect 16044 65314 16100 65324
rect 15708 65100 16212 65156
rect 15484 64654 15486 64706
rect 15538 64654 15540 64706
rect 15484 63138 15540 64654
rect 16044 64706 16100 64718
rect 16044 64654 16046 64706
rect 16098 64654 16100 64706
rect 16044 64148 16100 64654
rect 16156 64594 16212 65100
rect 16156 64542 16158 64594
rect 16210 64542 16212 64594
rect 16156 64530 16212 64542
rect 15484 63086 15486 63138
rect 15538 63086 15540 63138
rect 15484 62804 15540 63086
rect 15596 64092 16100 64148
rect 15596 63140 15652 64092
rect 15708 63924 15764 63934
rect 16268 63924 16324 65324
rect 16716 65314 16772 65324
rect 16828 64260 16884 67116
rect 16940 66948 16996 66958
rect 17388 66948 17444 67566
rect 17612 67060 17668 67070
rect 17724 67060 17780 67676
rect 17836 67666 17892 67676
rect 18620 67956 18676 67966
rect 17948 67060 18004 67070
rect 17612 67058 17780 67060
rect 17612 67006 17614 67058
rect 17666 67006 17780 67058
rect 17612 67004 17780 67006
rect 17836 67004 17948 67060
rect 17612 66994 17668 67004
rect 16940 66946 17108 66948
rect 16940 66894 16942 66946
rect 16994 66894 17108 66946
rect 16940 66892 17108 66894
rect 16940 66882 16996 66892
rect 16828 64146 16884 64204
rect 16828 64094 16830 64146
rect 16882 64094 16884 64146
rect 16828 64082 16884 64094
rect 16940 64594 16996 64606
rect 16940 64542 16942 64594
rect 16994 64542 16996 64594
rect 15708 63830 15764 63868
rect 15820 63922 16324 63924
rect 15820 63870 16270 63922
rect 16322 63870 16324 63922
rect 15820 63868 16324 63870
rect 15708 63140 15764 63150
rect 15596 63084 15708 63140
rect 15708 63074 15764 63084
rect 15484 62738 15540 62748
rect 15260 62626 15316 62636
rect 15372 62356 15428 62366
rect 15372 62262 15428 62300
rect 15820 62242 15876 63868
rect 16268 63858 16324 63868
rect 16380 64034 16436 64046
rect 16380 63982 16382 64034
rect 16434 63982 16436 64034
rect 16380 63924 16436 63982
rect 16380 63858 16436 63868
rect 16940 63364 16996 64542
rect 16268 63308 16996 63364
rect 16044 63140 16100 63150
rect 16044 63046 16100 63084
rect 16156 63028 16212 63038
rect 16156 62934 16212 62972
rect 15820 62190 15822 62242
rect 15874 62190 15876 62242
rect 15148 61572 15204 61582
rect 15148 61478 15204 61516
rect 15820 61124 15876 62190
rect 16268 62130 16324 63308
rect 16604 63140 16660 63150
rect 17052 63140 17108 66892
rect 17388 66882 17444 66892
rect 17388 66498 17444 66510
rect 17388 66446 17390 66498
rect 17442 66446 17444 66498
rect 17388 63922 17444 66446
rect 17724 66276 17780 66286
rect 17836 66276 17892 67004
rect 17948 66966 18004 67004
rect 18620 67060 18676 67900
rect 18620 66994 18676 67004
rect 18732 67058 18788 70252
rect 18844 68852 18900 70702
rect 18956 70196 19012 70206
rect 18956 70102 19012 70140
rect 18844 68786 18900 68796
rect 19292 67284 19348 75852
rect 19516 75842 19572 75852
rect 19628 76580 19684 76590
rect 19628 75684 19684 76524
rect 19404 75628 19684 75684
rect 20412 76356 20468 80332
rect 20524 80294 20580 80332
rect 20636 80388 20692 80398
rect 20636 80386 20916 80388
rect 20636 80334 20638 80386
rect 20690 80334 20916 80386
rect 20636 80332 20916 80334
rect 20636 80322 20692 80332
rect 20860 80276 20916 80332
rect 20860 80210 20916 80220
rect 20636 80164 20692 80174
rect 20636 80070 20692 80108
rect 20972 80052 21028 80444
rect 21532 80386 21588 80556
rect 21532 80334 21534 80386
rect 21586 80334 21588 80386
rect 21532 80322 21588 80334
rect 22092 80386 22148 80398
rect 22092 80334 22094 80386
rect 22146 80334 22148 80386
rect 20972 79986 21028 79996
rect 21532 80162 21588 80174
rect 21532 80110 21534 80162
rect 21586 80110 21588 80162
rect 21532 80052 21588 80110
rect 22092 80164 22148 80334
rect 22092 80098 22148 80108
rect 21532 79986 21588 79996
rect 22204 79828 22260 85652
rect 22316 85090 22372 85102
rect 22316 85038 22318 85090
rect 22370 85038 22372 85090
rect 22316 84532 22372 85038
rect 22652 85090 22708 86828
rect 22876 86772 22932 86782
rect 22652 85038 22654 85090
rect 22706 85038 22708 85090
rect 22652 85026 22708 85038
rect 22764 86716 22876 86772
rect 22764 86658 22820 86716
rect 22876 86706 22932 86716
rect 22764 86606 22766 86658
rect 22818 86606 22820 86658
rect 22372 84476 22484 84532
rect 22316 84466 22372 84476
rect 22316 84306 22372 84318
rect 22316 84254 22318 84306
rect 22370 84254 22372 84306
rect 22316 84084 22372 84254
rect 22316 84018 22372 84028
rect 22316 83298 22372 83310
rect 22316 83246 22318 83298
rect 22370 83246 22372 83298
rect 22316 82740 22372 83246
rect 22316 82674 22372 82684
rect 22428 81170 22484 84476
rect 22764 83972 22820 86606
rect 22988 85708 23044 87612
rect 23212 87602 23268 87612
rect 23548 87602 23604 87612
rect 23772 87668 23828 87678
rect 23772 87574 23828 87612
rect 23100 87330 23156 87342
rect 23100 87278 23102 87330
rect 23154 87278 23156 87330
rect 23100 86660 23156 87278
rect 23660 87330 23716 87342
rect 23660 87278 23662 87330
rect 23714 87278 23716 87330
rect 23212 86660 23268 86670
rect 23100 86658 23268 86660
rect 23100 86606 23214 86658
rect 23266 86606 23268 86658
rect 23100 86604 23268 86606
rect 23212 86594 23268 86604
rect 23548 86658 23604 86670
rect 23548 86606 23550 86658
rect 23602 86606 23604 86658
rect 23548 86100 23604 86606
rect 23660 86660 23716 87278
rect 23660 86594 23716 86604
rect 23772 86546 23828 86558
rect 23772 86494 23774 86546
rect 23826 86494 23828 86546
rect 23660 86436 23716 86446
rect 23660 86342 23716 86380
rect 23772 86100 23828 86494
rect 23548 86034 23604 86044
rect 23660 86044 23828 86100
rect 22876 85652 23044 85708
rect 23548 85874 23604 85886
rect 23548 85822 23550 85874
rect 23602 85822 23604 85874
rect 22876 84194 22932 85652
rect 23324 84420 23380 84430
rect 23324 84326 23380 84364
rect 22876 84142 22878 84194
rect 22930 84142 22932 84194
rect 22876 84130 22932 84142
rect 22988 84306 23044 84318
rect 22988 84254 22990 84306
rect 23042 84254 23044 84306
rect 22988 83972 23044 84254
rect 22764 83916 23044 83972
rect 22876 83410 22932 83422
rect 22876 83358 22878 83410
rect 22930 83358 22932 83410
rect 22876 83076 22932 83358
rect 22876 83010 22932 83020
rect 22988 82740 23044 83916
rect 22988 82674 23044 82684
rect 23436 84306 23492 84318
rect 23436 84254 23438 84306
rect 23490 84254 23492 84306
rect 23436 82066 23492 84254
rect 23436 82014 23438 82066
rect 23490 82014 23492 82066
rect 23436 82002 23492 82014
rect 23548 82626 23604 85822
rect 23548 82574 23550 82626
rect 23602 82574 23604 82626
rect 23100 81732 23156 81742
rect 22428 81118 22430 81170
rect 22482 81118 22484 81170
rect 22428 80276 22484 81118
rect 22204 79762 22260 79772
rect 22316 80052 22372 80062
rect 22316 79602 22372 79996
rect 22316 79550 22318 79602
rect 22370 79550 22372 79602
rect 22316 79538 22372 79550
rect 22428 79490 22484 80220
rect 22652 81284 22708 81294
rect 22652 81170 22708 81228
rect 22652 81118 22654 81170
rect 22706 81118 22708 81170
rect 22652 79602 22708 81118
rect 23100 81172 23156 81676
rect 23100 81078 23156 81116
rect 23324 81060 23380 81070
rect 22652 79550 22654 79602
rect 22706 79550 22708 79602
rect 22652 79538 22708 79550
rect 22764 80836 22820 80846
rect 22428 79438 22430 79490
rect 22482 79438 22484 79490
rect 22428 79426 22484 79438
rect 21196 79380 21252 79390
rect 21196 79378 21588 79380
rect 21196 79326 21198 79378
rect 21250 79326 21588 79378
rect 21196 79324 21588 79326
rect 21196 79314 21252 79324
rect 20524 78820 20580 78830
rect 20524 78726 20580 78764
rect 20636 78708 20692 78718
rect 20636 78614 20692 78652
rect 20748 78594 20804 78606
rect 20748 78542 20750 78594
rect 20802 78542 20804 78594
rect 20748 77364 20804 78542
rect 21532 77588 21588 79324
rect 21868 79378 21924 79390
rect 21868 79326 21870 79378
rect 21922 79326 21924 79378
rect 21644 78596 21700 78606
rect 21644 78502 21700 78540
rect 21868 78594 21924 79326
rect 22764 78820 22820 80780
rect 23324 79714 23380 81004
rect 23324 79662 23326 79714
rect 23378 79662 23380 79714
rect 23324 79650 23380 79662
rect 23436 79604 23492 79614
rect 23436 79510 23492 79548
rect 22652 78764 22820 78820
rect 21868 78542 21870 78594
rect 21922 78542 21924 78594
rect 21868 77700 21924 78542
rect 21868 77634 21924 77644
rect 21980 78594 22036 78606
rect 21980 78542 21982 78594
rect 22034 78542 22036 78594
rect 21532 77532 21700 77588
rect 21532 77364 21588 77374
rect 20748 77362 21588 77364
rect 20748 77310 21534 77362
rect 21586 77310 21588 77362
rect 20748 77308 21588 77310
rect 21532 77298 21588 77308
rect 20636 77250 20692 77262
rect 20636 77198 20638 77250
rect 20690 77198 20692 77250
rect 20636 76580 20692 77198
rect 20636 76486 20692 76524
rect 21644 76692 21700 77532
rect 20412 76300 20804 76356
rect 19404 73330 19460 75628
rect 20412 75572 20468 76300
rect 20748 75794 20804 76300
rect 20748 75742 20750 75794
rect 20802 75742 20804 75794
rect 20748 75730 20804 75742
rect 20412 75506 20468 75516
rect 21644 75682 21700 76636
rect 21980 75908 22036 78542
rect 22092 78594 22148 78606
rect 22092 78542 22094 78594
rect 22146 78542 22148 78594
rect 22092 77812 22148 78542
rect 22540 78596 22596 78606
rect 22540 78502 22596 78540
rect 22092 77746 22148 77756
rect 22540 78036 22596 78046
rect 21980 75842 22036 75852
rect 21644 75630 21646 75682
rect 21698 75630 21700 75682
rect 19836 75292 20100 75302
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 19836 75226 20100 75236
rect 19740 74788 19796 74798
rect 19740 74694 19796 74732
rect 19628 74340 19684 74350
rect 20076 74340 20132 74350
rect 19628 74338 20020 74340
rect 19628 74286 19630 74338
rect 19682 74286 20020 74338
rect 19628 74284 20020 74286
rect 19628 74274 19684 74284
rect 19964 74226 20020 74284
rect 19964 74174 19966 74226
rect 20018 74174 20020 74226
rect 19964 74162 20020 74174
rect 19852 74116 19908 74126
rect 19852 74022 19908 74060
rect 20076 74114 20132 74284
rect 21420 74340 21476 74350
rect 21420 74226 21476 74284
rect 21420 74174 21422 74226
rect 21474 74174 21476 74226
rect 21420 74162 21476 74174
rect 21644 74228 21700 75630
rect 22428 74900 22484 74910
rect 22204 74898 22484 74900
rect 22204 74846 22430 74898
rect 22482 74846 22484 74898
rect 22204 74844 22484 74846
rect 21868 74788 21924 74798
rect 21868 74786 22036 74788
rect 21868 74734 21870 74786
rect 21922 74734 22036 74786
rect 21868 74732 22036 74734
rect 21868 74722 21924 74732
rect 20076 74062 20078 74114
rect 20130 74062 20132 74114
rect 20076 74050 20132 74062
rect 20524 74114 20580 74126
rect 20524 74062 20526 74114
rect 20578 74062 20580 74114
rect 19740 74004 19796 74014
rect 19516 73892 19796 73948
rect 20524 74004 20580 74062
rect 20524 73938 20580 73948
rect 21644 73948 21700 74172
rect 21644 73892 21812 73948
rect 19516 73798 19572 73836
rect 19836 73724 20100 73734
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 19836 73658 20100 73668
rect 19404 73278 19406 73330
rect 19458 73278 19460 73330
rect 19404 73266 19460 73278
rect 21084 73220 21140 73230
rect 19964 72548 20020 72558
rect 19964 72454 20020 72492
rect 20412 72548 20468 72558
rect 20412 72454 20468 72492
rect 19836 72156 20100 72166
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 19836 72090 20100 72100
rect 21084 71650 21140 73164
rect 21084 71598 21086 71650
rect 21138 71598 21140 71650
rect 19836 70588 20100 70598
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 19836 70522 20100 70532
rect 19628 70084 19684 70094
rect 19628 69990 19684 70028
rect 19836 69020 20100 69030
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 19836 68954 20100 68964
rect 20748 68740 20804 68750
rect 20524 68684 20748 68740
rect 20300 68516 20356 68526
rect 19740 68514 20356 68516
rect 19740 68462 20302 68514
rect 20354 68462 20356 68514
rect 19740 68460 20356 68462
rect 19740 67954 19796 68460
rect 20300 68450 20356 68460
rect 19740 67902 19742 67954
rect 19794 67902 19796 67954
rect 19740 67890 19796 67902
rect 20188 67956 20244 67966
rect 20188 67862 20244 67900
rect 20524 67842 20580 68684
rect 20748 68646 20804 68684
rect 21084 68740 21140 71598
rect 21756 70308 21812 73892
rect 21868 71764 21924 71774
rect 21868 71670 21924 71708
rect 21756 70252 21924 70308
rect 21756 70084 21812 70094
rect 21084 68674 21140 68684
rect 21196 70082 21812 70084
rect 21196 70030 21758 70082
rect 21810 70030 21812 70082
rect 21196 70028 21812 70030
rect 21196 68738 21252 70028
rect 21756 70018 21812 70028
rect 21868 69860 21924 70252
rect 21196 68686 21198 68738
rect 21250 68686 21252 68738
rect 21196 68674 21252 68686
rect 21756 69804 21924 69860
rect 21084 68404 21140 68414
rect 20524 67790 20526 67842
rect 20578 67790 20580 67842
rect 20524 67778 20580 67790
rect 20636 68402 21140 68404
rect 20636 68350 21086 68402
rect 21138 68350 21140 68402
rect 20636 68348 21140 68350
rect 20636 67730 20692 68348
rect 21084 68338 21140 68348
rect 20636 67678 20638 67730
rect 20690 67678 20692 67730
rect 18732 67006 18734 67058
rect 18786 67006 18788 67058
rect 18732 66994 18788 67006
rect 18844 67228 19348 67284
rect 19404 67620 19460 67630
rect 18172 66948 18228 66958
rect 18172 66388 18228 66892
rect 17724 66274 17892 66276
rect 17724 66222 17726 66274
rect 17778 66222 17892 66274
rect 17724 66220 17892 66222
rect 17948 66274 18004 66286
rect 17948 66222 17950 66274
rect 18002 66222 18004 66274
rect 17724 66210 17780 66220
rect 17948 66164 18004 66222
rect 18172 66274 18228 66332
rect 18172 66222 18174 66274
rect 18226 66222 18228 66274
rect 18172 66210 18228 66222
rect 18620 66500 18676 66510
rect 17948 66098 18004 66108
rect 17500 65604 17556 65614
rect 17500 65510 17556 65548
rect 18620 64706 18676 66444
rect 18620 64654 18622 64706
rect 18674 64654 18676 64706
rect 18620 64642 18676 64654
rect 18732 66388 18788 66398
rect 18508 64482 18564 64494
rect 18508 64430 18510 64482
rect 18562 64430 18564 64482
rect 17948 64260 18004 64270
rect 17388 63870 17390 63922
rect 17442 63870 17444 63922
rect 17388 63858 17444 63870
rect 17500 64034 17556 64046
rect 17500 63982 17502 64034
rect 17554 63982 17556 64034
rect 17500 63924 17556 63982
rect 17500 63858 17556 63868
rect 17948 63140 18004 64204
rect 16660 63084 17108 63140
rect 17388 63138 18004 63140
rect 17388 63086 17950 63138
rect 18002 63086 18004 63138
rect 17388 63084 18004 63086
rect 16604 63026 16660 63084
rect 16604 62974 16606 63026
rect 16658 62974 16660 63026
rect 16492 62914 16548 62926
rect 16492 62862 16494 62914
rect 16546 62862 16548 62914
rect 16492 62354 16548 62862
rect 16492 62302 16494 62354
rect 16546 62302 16548 62354
rect 16492 62290 16548 62302
rect 16604 62244 16660 62974
rect 17276 63026 17332 63038
rect 17276 62974 17278 63026
rect 17330 62974 17332 63026
rect 16828 62916 16884 62926
rect 16716 62914 16884 62916
rect 16716 62862 16830 62914
rect 16882 62862 16884 62914
rect 16716 62860 16884 62862
rect 16716 62804 16772 62860
rect 16828 62850 16884 62860
rect 17052 62916 17108 62926
rect 17276 62916 17332 62974
rect 17052 62822 17108 62860
rect 17164 62860 17276 62916
rect 16716 62738 16772 62748
rect 16828 62692 16884 62702
rect 17164 62692 17220 62860
rect 17276 62850 17332 62860
rect 16884 62636 17220 62692
rect 16828 62578 16884 62636
rect 16828 62526 16830 62578
rect 16882 62526 16884 62578
rect 16828 62188 16884 62526
rect 17388 62188 17444 63084
rect 17948 63074 18004 63084
rect 18172 62804 18228 62814
rect 18172 62578 18228 62748
rect 18172 62526 18174 62578
rect 18226 62526 18228 62578
rect 18172 62356 18228 62526
rect 17724 62244 17780 62282
rect 16604 62178 16660 62188
rect 16268 62078 16270 62130
rect 16322 62078 16324 62130
rect 16268 62066 16324 62078
rect 16716 62132 16884 62188
rect 16940 62132 17444 62188
rect 17612 62188 17724 62244
rect 18172 62188 18228 62300
rect 16156 61794 16212 61806
rect 16156 61742 16158 61794
rect 16210 61742 16212 61794
rect 16156 61682 16212 61742
rect 16156 61630 16158 61682
rect 16210 61630 16212 61682
rect 16156 61618 16212 61630
rect 16716 61794 16772 62132
rect 16716 61742 16718 61794
rect 16770 61742 16772 61794
rect 16604 61348 16660 61358
rect 16492 61346 16660 61348
rect 16492 61294 16606 61346
rect 16658 61294 16660 61346
rect 16492 61292 16660 61294
rect 16492 61124 16548 61292
rect 16604 61282 16660 61292
rect 15820 61068 16548 61124
rect 16380 60116 16436 60126
rect 16156 60114 16436 60116
rect 16156 60062 16382 60114
rect 16434 60062 16436 60114
rect 16156 60060 16436 60062
rect 15484 59332 15540 59342
rect 15484 59238 15540 59276
rect 14588 59218 15092 59220
rect 14588 59166 14590 59218
rect 14642 59166 15092 59218
rect 14588 59164 15092 59166
rect 15708 59218 15764 59230
rect 15708 59166 15710 59218
rect 15762 59166 15764 59218
rect 14588 59154 14644 59164
rect 15148 59108 15204 59118
rect 15708 59108 15764 59166
rect 15148 59106 15764 59108
rect 15148 59054 15150 59106
rect 15202 59054 15764 59106
rect 15148 59052 15764 59054
rect 15148 59042 15204 59052
rect 14588 58996 14644 59006
rect 14812 58996 14868 59006
rect 14644 58994 14868 58996
rect 14644 58942 14814 58994
rect 14866 58942 14868 58994
rect 14644 58940 14868 58942
rect 14588 58930 14644 58940
rect 14476 58716 14756 58772
rect 14700 58546 14756 58716
rect 14700 58494 14702 58546
rect 14754 58494 14756 58546
rect 14700 58482 14756 58494
rect 14588 57876 14644 57886
rect 14588 56754 14644 57820
rect 14588 56702 14590 56754
rect 14642 56702 14644 56754
rect 14588 56690 14644 56702
rect 14700 56754 14756 56766
rect 14700 56702 14702 56754
rect 14754 56702 14756 56754
rect 14364 56644 14420 56654
rect 14364 56550 14420 56588
rect 14700 56420 14756 56702
rect 14140 56364 14756 56420
rect 14028 55300 14084 55310
rect 14140 55300 14196 56364
rect 14812 55412 14868 58940
rect 15036 58996 15092 59006
rect 15036 58436 15092 58940
rect 16044 58772 16100 58782
rect 15036 57538 15092 58380
rect 15036 57486 15038 57538
rect 15090 57486 15092 57538
rect 15036 57474 15092 57486
rect 15596 58660 15652 58670
rect 14812 55346 14868 55356
rect 15596 56642 15652 58604
rect 16044 57876 16100 58716
rect 16044 57782 16100 57820
rect 16156 57762 16212 60060
rect 16380 60050 16436 60060
rect 16492 59892 16548 61068
rect 16716 60676 16772 61742
rect 16156 57710 16158 57762
rect 16210 57710 16212 57762
rect 16156 57698 16212 57710
rect 16268 59836 16548 59892
rect 16604 60620 16772 60676
rect 16268 59220 16324 59836
rect 16268 57540 16324 59164
rect 16380 59108 16436 59118
rect 16380 59014 16436 59052
rect 16604 57876 16660 60620
rect 16828 59780 16884 59790
rect 16940 59780 16996 62132
rect 17612 61796 17668 62188
rect 17724 62178 17780 62188
rect 18060 62132 18228 62188
rect 18060 61796 18116 62132
rect 17164 61740 17668 61796
rect 17724 61740 18116 61796
rect 17052 61458 17108 61470
rect 17052 61406 17054 61458
rect 17106 61406 17108 61458
rect 17052 61348 17108 61406
rect 17164 61348 17220 61740
rect 17724 61684 17780 61740
rect 17052 61292 17164 61348
rect 17164 61282 17220 61292
rect 17276 61682 17780 61684
rect 17276 61630 17726 61682
rect 17778 61630 17780 61682
rect 17276 61628 17780 61630
rect 16828 59778 16996 59780
rect 16828 59726 16830 59778
rect 16882 59726 16996 59778
rect 16828 59724 16996 59726
rect 16828 59106 16884 59724
rect 16828 59054 16830 59106
rect 16882 59054 16884 59106
rect 16828 58772 16884 59054
rect 16716 58716 16884 58772
rect 16716 58660 16772 58716
rect 16716 58594 16772 58604
rect 16828 58546 16884 58558
rect 16828 58494 16830 58546
rect 16882 58494 16884 58546
rect 16828 58212 16884 58494
rect 16828 58146 16884 58156
rect 17276 58322 17332 61628
rect 17724 61618 17780 61628
rect 17948 61348 18004 61358
rect 17836 60340 17892 60350
rect 17724 60284 17836 60340
rect 17500 59332 17556 59342
rect 17500 59238 17556 59276
rect 17388 59220 17444 59230
rect 17388 59126 17444 59164
rect 17612 59218 17668 59230
rect 17612 59166 17614 59218
rect 17666 59166 17668 59218
rect 17612 58772 17668 59166
rect 17612 58706 17668 58716
rect 17276 58270 17278 58322
rect 17330 58270 17332 58322
rect 17276 58100 17332 58270
rect 17276 58034 17332 58044
rect 17612 58212 17668 58222
rect 16940 57988 16996 57998
rect 16828 57876 16884 57886
rect 16604 57874 16884 57876
rect 16604 57822 16830 57874
rect 16882 57822 16884 57874
rect 16604 57820 16884 57822
rect 16828 57764 16884 57820
rect 16828 57698 16884 57708
rect 15596 56590 15598 56642
rect 15650 56590 15652 56642
rect 14084 55244 14196 55300
rect 13804 53620 13860 53630
rect 13804 53526 13860 53564
rect 13804 49028 13860 49038
rect 13804 48934 13860 48972
rect 11900 48804 11956 48814
rect 11900 48354 11956 48748
rect 11900 48302 11902 48354
rect 11954 48302 11956 48354
rect 11900 48290 11956 48302
rect 12908 48804 12964 48814
rect 12348 48132 12404 48142
rect 12236 48076 12348 48132
rect 12236 45668 12292 48076
rect 12348 48038 12404 48076
rect 12796 48130 12852 48142
rect 12796 48078 12798 48130
rect 12850 48078 12852 48130
rect 12796 48020 12852 48078
rect 12796 47954 12852 47964
rect 12908 47570 12964 48748
rect 13020 48802 13076 48860
rect 13020 48750 13022 48802
rect 13074 48750 13076 48802
rect 13020 48132 13076 48750
rect 13020 48066 13076 48076
rect 13468 48860 13748 48916
rect 12908 47518 12910 47570
rect 12962 47518 12964 47570
rect 12908 47506 12964 47518
rect 13132 47348 13188 47358
rect 12908 45892 12964 45902
rect 12908 45798 12964 45836
rect 11900 44996 11956 45006
rect 11900 44902 11956 44940
rect 12236 44660 12292 45612
rect 11676 38612 11844 38668
rect 12012 44604 12292 44660
rect 12460 44996 12516 45006
rect 12012 38668 12068 44604
rect 12124 43428 12180 43438
rect 12124 43426 12404 43428
rect 12124 43374 12126 43426
rect 12178 43374 12404 43426
rect 12124 43372 12404 43374
rect 12124 43362 12180 43372
rect 12348 42642 12404 43372
rect 12348 42590 12350 42642
rect 12402 42590 12404 42642
rect 12348 42578 12404 42590
rect 12460 42084 12516 44940
rect 12572 42754 12628 42766
rect 12572 42702 12574 42754
rect 12626 42702 12628 42754
rect 12572 42194 12628 42702
rect 12572 42142 12574 42194
rect 12626 42142 12628 42194
rect 12572 42130 12628 42142
rect 12236 42028 12516 42084
rect 12236 39172 12292 42028
rect 13132 41970 13188 47292
rect 13468 46114 13524 48860
rect 13916 48468 13972 48478
rect 13916 48374 13972 48412
rect 13692 47572 13748 47582
rect 13580 47236 13636 47246
rect 13580 47142 13636 47180
rect 13468 46062 13470 46114
rect 13522 46062 13524 46114
rect 13468 46050 13524 46062
rect 13692 46116 13748 47516
rect 13804 46900 13860 46910
rect 14028 46900 14084 55244
rect 15148 54404 15204 54414
rect 14700 54402 15204 54404
rect 14700 54350 15150 54402
rect 15202 54350 15204 54402
rect 14700 54348 15204 54350
rect 14252 53508 14308 53518
rect 14252 53414 14308 53452
rect 14700 52274 14756 54348
rect 15148 54338 15204 54348
rect 15596 54402 15652 56590
rect 15596 54350 15598 54402
rect 15650 54350 15652 54402
rect 14700 52222 14702 52274
rect 14754 52222 14756 52274
rect 14700 52210 14756 52222
rect 14812 54068 14868 54078
rect 14588 51938 14644 51950
rect 14588 51886 14590 51938
rect 14642 51886 14644 51938
rect 14364 49812 14420 49822
rect 14588 49812 14644 51886
rect 14700 50708 14756 50718
rect 14812 50708 14868 54012
rect 15596 54068 15652 54350
rect 15596 54002 15652 54012
rect 16156 57484 16324 57540
rect 15820 53732 15876 53742
rect 15260 53172 15316 53182
rect 15148 53116 15260 53172
rect 15148 53058 15204 53116
rect 15260 53106 15316 53116
rect 15148 53006 15150 53058
rect 15202 53006 15204 53058
rect 15148 52994 15204 53006
rect 15820 52946 15876 53676
rect 15820 52894 15822 52946
rect 15874 52894 15876 52946
rect 15820 52882 15876 52894
rect 16044 52948 16100 52958
rect 15596 52164 15652 52174
rect 15596 52070 15652 52108
rect 16044 52050 16100 52892
rect 16044 51998 16046 52050
rect 16098 51998 16100 52050
rect 16044 51986 16100 51998
rect 15372 51940 15428 51950
rect 15820 51940 15876 51950
rect 15372 51938 15876 51940
rect 15372 51886 15374 51938
rect 15426 51886 15822 51938
rect 15874 51886 15876 51938
rect 15372 51884 15876 51886
rect 15372 51874 15428 51884
rect 15820 51716 15876 51884
rect 15820 51650 15876 51660
rect 15932 51938 15988 51950
rect 15932 51886 15934 51938
rect 15986 51886 15988 51938
rect 15932 51492 15988 51886
rect 15708 51436 15988 51492
rect 14700 50706 14980 50708
rect 14700 50654 14702 50706
rect 14754 50654 14980 50706
rect 14700 50652 14980 50654
rect 14700 50642 14756 50652
rect 14588 49756 14756 49812
rect 14140 48916 14196 48926
rect 14140 48822 14196 48860
rect 14252 48804 14308 48814
rect 14252 48710 14308 48748
rect 14364 48356 14420 49756
rect 14476 49700 14532 49710
rect 14476 49698 14644 49700
rect 14476 49646 14478 49698
rect 14530 49646 14644 49698
rect 14476 49644 14644 49646
rect 14476 49634 14532 49644
rect 14476 49252 14532 49262
rect 14476 49026 14532 49196
rect 14476 48974 14478 49026
rect 14530 48974 14532 49026
rect 14476 48962 14532 48974
rect 14364 48300 14532 48356
rect 14364 48130 14420 48142
rect 14364 48078 14366 48130
rect 14418 48078 14420 48130
rect 13804 46898 14084 46900
rect 13804 46846 13806 46898
rect 13858 46846 14084 46898
rect 13804 46844 14084 46846
rect 13804 46834 13860 46844
rect 14028 46788 14084 46844
rect 14252 47682 14308 47694
rect 14252 47630 14254 47682
rect 14306 47630 14308 47682
rect 14252 46898 14308 47630
rect 14364 47570 14420 48078
rect 14364 47518 14366 47570
rect 14418 47518 14420 47570
rect 14364 47236 14420 47518
rect 14364 47170 14420 47180
rect 14252 46846 14254 46898
rect 14306 46846 14308 46898
rect 14252 46834 14308 46846
rect 14140 46788 14196 46798
rect 14028 46786 14196 46788
rect 14028 46734 14142 46786
rect 14194 46734 14196 46786
rect 14028 46732 14196 46734
rect 14140 46722 14196 46732
rect 14252 46450 14308 46462
rect 14252 46398 14254 46450
rect 14306 46398 14308 46450
rect 13692 46060 14084 46116
rect 14028 46004 14084 46060
rect 14028 46002 14196 46004
rect 14028 45950 14030 46002
rect 14082 45950 14196 46002
rect 14028 45948 14196 45950
rect 14028 45938 14084 45948
rect 13804 45892 13860 45902
rect 13860 45836 13972 45892
rect 13804 45798 13860 45836
rect 13132 41918 13134 41970
rect 13186 41918 13188 41970
rect 12348 41860 12404 41870
rect 12908 41860 12964 41870
rect 12348 41858 12964 41860
rect 12348 41806 12350 41858
rect 12402 41806 12910 41858
rect 12962 41806 12964 41858
rect 12348 41804 12964 41806
rect 12348 41794 12404 41804
rect 12460 39396 12516 39406
rect 12460 39302 12516 39340
rect 12236 39116 12516 39172
rect 12012 38612 12180 38668
rect 11452 38052 11508 38062
rect 11452 37958 11508 37996
rect 11676 37156 11732 38612
rect 11676 37062 11732 37100
rect 12012 37044 12068 37054
rect 11788 37042 12068 37044
rect 11788 36990 12014 37042
rect 12066 36990 12068 37042
rect 11788 36988 12068 36990
rect 11788 36932 11844 36988
rect 12012 36978 12068 36988
rect 11676 36876 11844 36932
rect 11676 36482 11732 36876
rect 11676 36430 11678 36482
rect 11730 36430 11732 36482
rect 11676 36418 11732 36430
rect 12012 36596 12068 36606
rect 11452 36260 11508 36270
rect 11004 35868 11172 35924
rect 11228 36258 11508 36260
rect 11228 36206 11454 36258
rect 11506 36206 11508 36258
rect 11228 36204 11508 36206
rect 11004 30212 11060 35868
rect 11116 35700 11172 35710
rect 11116 35606 11172 35644
rect 11228 35474 11284 36204
rect 11452 36194 11508 36204
rect 12012 35698 12068 36540
rect 12012 35646 12014 35698
rect 12066 35646 12068 35698
rect 12012 35634 12068 35646
rect 11228 35422 11230 35474
rect 11282 35422 11284 35474
rect 11228 35410 11284 35422
rect 11564 34020 11620 34030
rect 11620 33964 11732 34020
rect 11564 33954 11620 33964
rect 11676 33572 11732 33964
rect 11676 32564 11732 33516
rect 11788 32564 11844 32574
rect 11676 32562 11844 32564
rect 11676 32510 11790 32562
rect 11842 32510 11844 32562
rect 11676 32508 11844 32510
rect 11788 32498 11844 32508
rect 11004 30146 11060 30156
rect 10780 30044 10948 30100
rect 10780 29988 10836 30044
rect 11004 29988 11060 29998
rect 10556 29426 10612 29596
rect 10556 29374 10558 29426
rect 10610 29374 10612 29426
rect 10556 29362 10612 29374
rect 10668 29932 10836 29988
rect 10892 29986 11060 29988
rect 10892 29934 11006 29986
rect 11058 29934 11060 29986
rect 10892 29932 11060 29934
rect 10556 27860 10612 27870
rect 10332 26852 10500 26908
rect 10332 24612 10388 24622
rect 10332 24518 10388 24556
rect 10108 22652 10276 22708
rect 9772 22596 9828 22606
rect 9828 22540 9940 22596
rect 9772 22530 9828 22540
rect 9324 22260 9380 22270
rect 9324 22258 9604 22260
rect 9324 22206 9326 22258
rect 9378 22206 9604 22258
rect 9324 22204 9604 22206
rect 9324 22194 9380 22204
rect 9548 21810 9604 22204
rect 9548 21758 9550 21810
rect 9602 21758 9604 21810
rect 9548 21746 9604 21758
rect 9772 21588 9828 21598
rect 8876 21422 8878 21474
rect 8930 21422 8932 21474
rect 8876 21410 8932 21422
rect 8988 21586 9828 21588
rect 8988 21534 9774 21586
rect 9826 21534 9828 21586
rect 8988 21532 9828 21534
rect 8988 21026 9044 21532
rect 9772 21522 9828 21532
rect 9884 21364 9940 22540
rect 8988 20974 8990 21026
rect 9042 20974 9044 21026
rect 8988 20962 9044 20974
rect 9548 21308 9940 21364
rect 9548 20914 9604 21308
rect 9548 20862 9550 20914
rect 9602 20862 9604 20914
rect 9548 20850 9604 20862
rect 8428 20750 8430 20802
rect 8482 20750 8484 20802
rect 8092 20578 8148 20590
rect 8092 20526 8094 20578
rect 8146 20526 8148 20578
rect 8092 20244 8148 20526
rect 8092 20178 8148 20188
rect 8428 18452 8484 20750
rect 8652 20802 8708 20814
rect 8652 20750 8654 20802
rect 8706 20750 8708 20802
rect 8652 20244 8708 20750
rect 8652 20178 8708 20188
rect 9548 18562 9604 18574
rect 9548 18510 9550 18562
rect 9602 18510 9604 18562
rect 8316 18396 8484 18452
rect 9324 18452 9380 18462
rect 7980 17948 8148 18004
rect 7980 17778 8036 17790
rect 7980 17726 7982 17778
rect 8034 17726 8036 17778
rect 7980 15988 8036 17726
rect 7980 15922 8036 15932
rect 8092 15540 8148 17948
rect 8204 16772 8260 16782
rect 8316 16772 8372 18396
rect 8204 16770 8372 16772
rect 8204 16718 8206 16770
rect 8258 16718 8372 16770
rect 8204 16716 8372 16718
rect 8652 17108 8708 17118
rect 8204 16706 8260 16716
rect 8652 16098 8708 17052
rect 9324 16210 9380 18396
rect 9548 17780 9604 18510
rect 9884 18452 9940 18462
rect 10108 18452 10164 22652
rect 10332 18562 10388 18574
rect 10332 18510 10334 18562
rect 10386 18510 10388 18562
rect 9884 18450 10164 18452
rect 9884 18398 9886 18450
rect 9938 18398 10164 18450
rect 9884 18396 10164 18398
rect 10220 18452 10276 18462
rect 10332 18452 10388 18510
rect 10276 18396 10388 18452
rect 9884 18386 9940 18396
rect 10220 18386 10276 18396
rect 10444 18340 10500 26852
rect 10556 23380 10612 27804
rect 10556 23286 10612 23324
rect 10668 21028 10724 29932
rect 10780 29540 10836 29550
rect 10780 29446 10836 29484
rect 10780 28756 10836 28766
rect 10892 28756 10948 29932
rect 11004 29922 11060 29932
rect 11340 29540 11396 29550
rect 11340 29314 11396 29484
rect 11340 29262 11342 29314
rect 11394 29262 11396 29314
rect 11340 29250 11396 29262
rect 10780 28754 10948 28756
rect 10780 28702 10782 28754
rect 10834 28702 10948 28754
rect 10780 28700 10948 28702
rect 10780 28690 10836 28700
rect 12124 26908 12180 38612
rect 11900 26852 12180 26908
rect 12236 37156 12292 37166
rect 12236 37044 12292 37100
rect 12348 37044 12404 37054
rect 12236 37042 12404 37044
rect 12236 36990 12350 37042
rect 12402 36990 12404 37042
rect 12236 36988 12404 36990
rect 12236 34018 12292 36988
rect 12348 36978 12404 36988
rect 12236 33966 12238 34018
rect 12290 33966 12292 34018
rect 12236 33908 12292 33966
rect 12236 31668 12292 33852
rect 11564 23266 11620 23278
rect 11564 23214 11566 23266
rect 11618 23214 11620 23266
rect 11004 23156 11060 23166
rect 11004 23042 11060 23100
rect 11004 22990 11006 23042
rect 11058 22990 11060 23042
rect 11004 22148 11060 22990
rect 11452 22484 11508 22494
rect 11452 22390 11508 22428
rect 11004 22082 11060 22092
rect 11564 21698 11620 23214
rect 11788 23154 11844 23166
rect 11788 23102 11790 23154
rect 11842 23102 11844 23154
rect 11788 22594 11844 23102
rect 11788 22542 11790 22594
rect 11842 22542 11844 22594
rect 11788 22530 11844 22542
rect 11564 21646 11566 21698
rect 11618 21646 11620 21698
rect 11564 21634 11620 21646
rect 10892 21588 10948 21598
rect 10892 21494 10948 21532
rect 10332 18284 10500 18340
rect 10556 20972 10724 21028
rect 10108 17780 10164 17790
rect 9548 17778 10164 17780
rect 9548 17726 10110 17778
rect 10162 17726 10164 17778
rect 9548 17724 10164 17726
rect 10108 17714 10164 17724
rect 9324 16158 9326 16210
rect 9378 16158 9380 16210
rect 9324 16146 9380 16158
rect 10220 16212 10276 16222
rect 8652 16046 8654 16098
rect 8706 16046 8708 16098
rect 8652 16034 8708 16046
rect 8092 15474 8148 15484
rect 8988 15540 9044 15550
rect 8988 15446 9044 15484
rect 10220 15540 10276 16156
rect 10220 15314 10276 15484
rect 10220 15262 10222 15314
rect 10274 15262 10276 15314
rect 10220 15250 10276 15262
rect 9884 15090 9940 15102
rect 9884 15038 9886 15090
rect 9938 15038 9940 15090
rect 8316 13860 8372 13870
rect 7980 13748 8036 13758
rect 7980 13654 8036 13692
rect 8316 13074 8372 13804
rect 9548 13860 9604 13870
rect 9548 13766 9604 13804
rect 9884 13858 9940 15038
rect 9884 13806 9886 13858
rect 9938 13806 9940 13858
rect 9884 13794 9940 13806
rect 8316 13022 8318 13074
rect 8370 13022 8372 13074
rect 8316 13010 8372 13022
rect 8092 12404 8148 12414
rect 8092 12310 8148 12348
rect 9884 12404 9940 12414
rect 8428 12178 8484 12190
rect 8428 12126 8430 12178
rect 8482 12126 8484 12178
rect 8428 12068 8484 12126
rect 9884 12178 9940 12348
rect 9884 12126 9886 12178
rect 9938 12126 9940 12178
rect 9884 12114 9940 12126
rect 8428 12002 8484 12012
rect 8988 12068 9044 12078
rect 8988 11974 9044 12012
rect 10108 12066 10164 12078
rect 10108 12014 10110 12066
rect 10162 12014 10164 12066
rect 9548 11954 9604 11966
rect 9548 11902 9550 11954
rect 9602 11902 9604 11954
rect 8988 11732 9044 11742
rect 8988 11396 9044 11676
rect 9100 11396 9156 11406
rect 8988 11394 9156 11396
rect 8988 11342 9102 11394
rect 9154 11342 9156 11394
rect 8988 11340 9156 11342
rect 8988 10834 9044 11340
rect 9100 11330 9156 11340
rect 8988 10782 8990 10834
rect 9042 10782 9044 10834
rect 8988 10770 9044 10782
rect 9548 10722 9604 11902
rect 9884 11282 9940 11294
rect 9884 11230 9886 11282
rect 9938 11230 9940 11282
rect 9884 10834 9940 11230
rect 10108 10948 10164 12014
rect 9884 10782 9886 10834
rect 9938 10782 9940 10834
rect 9884 10770 9940 10782
rect 9996 10892 10164 10948
rect 9548 10670 9550 10722
rect 9602 10670 9604 10722
rect 9548 10658 9604 10670
rect 8540 10498 8596 10510
rect 8540 10446 8542 10498
rect 8594 10446 8596 10498
rect 8540 10388 8596 10446
rect 8540 10322 8596 10332
rect 9996 10388 10052 10892
rect 9996 10322 10052 10332
rect 10108 10724 10164 10734
rect 8988 9268 9044 9278
rect 8988 9174 9044 9212
rect 9884 9268 9940 9278
rect 9884 9042 9940 9212
rect 9884 8990 9886 9042
rect 9938 8990 9940 9042
rect 9884 8978 9940 8990
rect 10108 9042 10164 10668
rect 10220 10612 10276 10622
rect 10220 10518 10276 10556
rect 10108 8990 10110 9042
rect 10162 8990 10164 9042
rect 10108 8978 10164 8990
rect 9548 8820 9604 8830
rect 9100 8818 9604 8820
rect 9100 8766 9550 8818
rect 9602 8766 9604 8818
rect 9100 8764 9604 8766
rect 8876 8260 8932 8270
rect 9100 8260 9156 8764
rect 9548 8754 9604 8764
rect 8876 8258 9156 8260
rect 8876 8206 8878 8258
rect 8930 8206 9156 8258
rect 8876 8204 9156 8206
rect 8876 8194 8932 8204
rect 8540 8036 8596 8046
rect 7980 8034 8596 8036
rect 7980 7982 8542 8034
rect 8594 7982 8596 8034
rect 7980 7980 8596 7982
rect 7980 6690 8036 7980
rect 8540 7970 8596 7980
rect 10220 7586 10276 7598
rect 10220 7534 10222 7586
rect 10274 7534 10276 7586
rect 9996 7474 10052 7486
rect 9996 7422 9998 7474
rect 10050 7422 10052 7474
rect 7980 6638 7982 6690
rect 8034 6638 8036 6690
rect 7980 6626 8036 6638
rect 8652 7252 8708 7262
rect 7868 6412 8148 6468
rect 5292 5170 5348 5180
rect 6412 5236 6468 5246
rect 5628 4900 5684 4910
rect 5628 4226 5684 4844
rect 5628 4174 5630 4226
rect 5682 4174 5684 4226
rect 5628 4162 5684 4174
rect 4732 2156 4900 2212
rect 6188 3442 6244 3454
rect 6188 3390 6190 3442
rect 6242 3390 6244 3442
rect 4396 1876 4452 1886
rect 4284 1874 4452 1876
rect 4284 1822 4398 1874
rect 4450 1822 4452 1874
rect 4284 1820 4452 1822
rect 4396 1810 4452 1820
rect 3388 1148 4116 1204
rect 3836 400 3892 1148
rect 4732 400 4788 2156
rect 5852 1876 5908 1886
rect 5628 1820 5852 1876
rect 5068 1764 5124 1774
rect 5068 1670 5124 1708
rect 5628 400 5684 1820
rect 5852 1782 5908 1820
rect 6188 1874 6244 3390
rect 6300 3444 6356 3482
rect 6300 3378 6356 3388
rect 6412 2882 6468 5180
rect 7980 4900 8036 4910
rect 7756 4898 8036 4900
rect 7756 4846 7982 4898
rect 8034 4846 8036 4898
rect 7756 4844 8036 4846
rect 7756 4450 7812 4844
rect 7980 4834 8036 4844
rect 7756 4398 7758 4450
rect 7810 4398 7812 4450
rect 7756 4386 7812 4398
rect 8092 4564 8148 6412
rect 8652 5572 8708 7196
rect 8988 7140 9044 7150
rect 8652 5122 8708 5516
rect 8652 5070 8654 5122
rect 8706 5070 8708 5122
rect 8652 5058 8708 5070
rect 8876 7084 8988 7140
rect 8316 5012 8372 5022
rect 8092 3666 8148 4508
rect 8204 5010 8372 5012
rect 8204 4958 8318 5010
rect 8370 4958 8372 5010
rect 8204 4956 8372 4958
rect 8204 4116 8260 4956
rect 8316 4946 8372 4956
rect 8764 4898 8820 4910
rect 8764 4846 8766 4898
rect 8818 4846 8820 4898
rect 8764 4676 8820 4846
rect 8204 4050 8260 4060
rect 8316 4620 8820 4676
rect 8092 3614 8094 3666
rect 8146 3614 8148 3666
rect 8092 3602 8148 3614
rect 7532 3556 7588 3566
rect 7420 3444 7476 3482
rect 7420 3378 7476 3388
rect 7532 3220 7588 3500
rect 8316 3556 8372 4620
rect 8876 4564 8932 7084
rect 8988 7074 9044 7084
rect 9996 6692 10052 7422
rect 10108 6804 10164 6814
rect 10108 6710 10164 6748
rect 9996 6626 10052 6636
rect 9660 6580 9716 6590
rect 9660 5906 9716 6524
rect 10220 6132 10276 7534
rect 10332 7140 10388 18284
rect 10444 15316 10500 15326
rect 10444 15222 10500 15260
rect 10556 15148 10612 20972
rect 11116 20244 11172 20254
rect 11116 19906 11172 20188
rect 11116 19854 11118 19906
rect 11170 19854 11172 19906
rect 11116 19796 11172 19854
rect 11452 19796 11508 19806
rect 11116 19730 11172 19740
rect 11228 19794 11508 19796
rect 11228 19742 11454 19794
rect 11506 19742 11508 19794
rect 11228 19740 11508 19742
rect 11228 19124 11284 19740
rect 11452 19730 11508 19740
rect 11788 19796 11844 19806
rect 11788 19702 11844 19740
rect 10668 19068 11284 19124
rect 10668 18562 10724 19068
rect 10668 18510 10670 18562
rect 10722 18510 10724 18562
rect 10668 18498 10724 18510
rect 10780 17666 10836 17678
rect 10780 17614 10782 17666
rect 10834 17614 10836 17666
rect 10780 17444 10836 17614
rect 11788 17556 11844 17566
rect 11340 17444 11396 17454
rect 11788 17444 11844 17500
rect 10780 17442 11844 17444
rect 10780 17390 11342 17442
rect 11394 17390 11844 17442
rect 10780 17388 11844 17390
rect 10780 17108 10836 17388
rect 11340 17378 11396 17388
rect 10780 17042 10836 17052
rect 11788 16884 11844 17388
rect 11676 16882 11844 16884
rect 11676 16830 11790 16882
rect 11842 16830 11844 16882
rect 11676 16828 11844 16830
rect 11452 16210 11508 16222
rect 11452 16158 11454 16210
rect 11506 16158 11508 16210
rect 11452 15876 11508 16158
rect 11452 15316 11508 15820
rect 11452 15250 11508 15260
rect 11676 15538 11732 16828
rect 11788 16818 11844 16828
rect 11900 16100 11956 26852
rect 12124 23044 12180 23054
rect 12124 22370 12180 22988
rect 12124 22318 12126 22370
rect 12178 22318 12180 22370
rect 12012 20916 12068 20926
rect 12012 20018 12068 20860
rect 12012 19966 12014 20018
rect 12066 19966 12068 20018
rect 12012 19954 12068 19966
rect 12124 19796 12180 22318
rect 12124 16212 12180 19740
rect 12236 16772 12292 31612
rect 12460 26908 12516 39116
rect 12572 37268 12628 37278
rect 12572 37174 12628 37212
rect 12684 37044 12740 41804
rect 12908 41794 12964 41804
rect 13132 41636 13188 41918
rect 12796 41580 13188 41636
rect 13244 41972 13300 41982
rect 12796 40290 12852 41580
rect 12908 41300 12964 41310
rect 12908 41206 12964 41244
rect 12796 40238 12798 40290
rect 12850 40238 12852 40290
rect 12796 40226 12852 40238
rect 13020 40628 13076 40638
rect 12908 39620 12964 39630
rect 12908 39526 12964 39564
rect 13020 39058 13076 40572
rect 13244 40628 13300 41916
rect 13580 40964 13636 40974
rect 13580 40962 13748 40964
rect 13580 40910 13582 40962
rect 13634 40910 13748 40962
rect 13580 40908 13748 40910
rect 13580 40898 13636 40908
rect 13692 40628 13748 40908
rect 13244 40626 13636 40628
rect 13244 40574 13246 40626
rect 13298 40574 13636 40626
rect 13244 40572 13636 40574
rect 13244 40562 13300 40572
rect 13580 40516 13636 40572
rect 13692 40516 13748 40572
rect 13804 40516 13860 40526
rect 13692 40460 13804 40516
rect 13580 40422 13636 40460
rect 13804 40450 13860 40460
rect 13020 39006 13022 39058
rect 13074 39006 13076 39058
rect 13020 38994 13076 39006
rect 13804 39618 13860 39630
rect 13804 39566 13806 39618
rect 13858 39566 13860 39618
rect 13356 38722 13412 38734
rect 13356 38670 13358 38722
rect 13410 38670 13412 38722
rect 13356 38164 13412 38670
rect 13804 38668 13860 39566
rect 13356 38098 13412 38108
rect 13692 38612 13860 38668
rect 13468 37380 13524 37390
rect 12684 36978 12740 36988
rect 12796 37378 13524 37380
rect 12796 37326 13470 37378
rect 13522 37326 13524 37378
rect 12796 37324 13524 37326
rect 12796 35810 12852 37324
rect 13468 37314 13524 37324
rect 13020 37156 13076 37166
rect 13020 37062 13076 37100
rect 12796 35758 12798 35810
rect 12850 35758 12852 35810
rect 12796 35746 12852 35758
rect 12908 35700 12964 35710
rect 12908 35028 12964 35644
rect 12908 35026 13188 35028
rect 12908 34974 12910 35026
rect 12962 34974 13188 35026
rect 12908 34972 13188 34974
rect 12908 34962 12964 34972
rect 13132 34130 13188 34972
rect 13132 34078 13134 34130
rect 13186 34078 13188 34130
rect 13132 34066 13188 34078
rect 13580 34690 13636 34702
rect 13580 34638 13582 34690
rect 13634 34638 13636 34690
rect 12572 33906 12628 33918
rect 12572 33854 12574 33906
rect 12626 33854 12628 33906
rect 12572 33346 12628 33854
rect 12684 33908 12740 33918
rect 12908 33908 12964 33918
rect 12740 33906 12964 33908
rect 12740 33854 12910 33906
rect 12962 33854 12964 33906
rect 12740 33852 12964 33854
rect 12684 33842 12740 33852
rect 12908 33842 12964 33852
rect 12572 33294 12574 33346
rect 12626 33294 12628 33346
rect 12572 33282 12628 33294
rect 13580 33572 13636 34638
rect 12796 33124 12852 33134
rect 12572 33122 12852 33124
rect 12572 33070 12798 33122
rect 12850 33070 12852 33122
rect 12572 33068 12852 33070
rect 12572 32674 12628 33068
rect 12796 33058 12852 33068
rect 12572 32622 12574 32674
rect 12626 32622 12628 32674
rect 12572 32610 12628 32622
rect 13580 32564 13636 33516
rect 13580 32498 13636 32508
rect 12684 30210 12740 30222
rect 12684 30158 12686 30210
rect 12738 30158 12740 30210
rect 12684 28868 12740 30158
rect 12908 29988 12964 29998
rect 12908 29986 13524 29988
rect 12908 29934 12910 29986
rect 12962 29934 13524 29986
rect 12908 29932 13524 29934
rect 12908 29922 12964 29932
rect 12684 28802 12740 28812
rect 13244 29652 13300 29662
rect 12908 28754 12964 28766
rect 12908 28702 12910 28754
rect 12962 28702 12964 28754
rect 12908 28196 12964 28702
rect 12908 28130 12964 28140
rect 13244 28082 13300 29596
rect 13468 29538 13524 29932
rect 13468 29486 13470 29538
rect 13522 29486 13524 29538
rect 13468 29474 13524 29486
rect 13468 28868 13524 28878
rect 13468 28774 13524 28812
rect 13244 28030 13246 28082
rect 13298 28030 13300 28082
rect 13244 28018 13300 28030
rect 13580 28644 13636 28654
rect 13580 28082 13636 28588
rect 13580 28030 13582 28082
rect 13634 28030 13636 28082
rect 13580 28018 13636 28030
rect 13468 27748 13524 27758
rect 13468 27186 13524 27692
rect 13468 27134 13470 27186
rect 13522 27134 13524 27186
rect 13468 27122 13524 27134
rect 12460 26852 13412 26908
rect 12684 25396 12740 25406
rect 12684 25302 12740 25340
rect 13244 25396 13300 25406
rect 13020 25172 13076 25182
rect 13020 24724 13076 25116
rect 12460 24722 13076 24724
rect 12460 24670 13022 24722
rect 13074 24670 13076 24722
rect 12460 24668 13076 24670
rect 12460 24610 12516 24668
rect 13020 24658 13076 24668
rect 12460 24558 12462 24610
rect 12514 24558 12516 24610
rect 12460 24546 12516 24558
rect 13244 24500 13300 25340
rect 13132 24498 13300 24500
rect 13132 24446 13246 24498
rect 13298 24446 13300 24498
rect 13132 24444 13300 24446
rect 12796 24164 12852 24174
rect 12796 24070 12852 24108
rect 12684 23826 12740 23838
rect 12684 23774 12686 23826
rect 12738 23774 12740 23826
rect 12348 23714 12404 23726
rect 12348 23662 12350 23714
rect 12402 23662 12404 23714
rect 12348 23604 12404 23662
rect 12348 23538 12404 23548
rect 12684 23604 12740 23774
rect 12684 23538 12740 23548
rect 12796 23714 12852 23726
rect 12796 23662 12798 23714
rect 12850 23662 12852 23714
rect 12348 23044 12404 23054
rect 12348 22950 12404 22988
rect 12796 22820 12852 23662
rect 12348 22764 12852 22820
rect 12348 22484 12404 22764
rect 12348 22390 12404 22428
rect 12796 22596 12852 22606
rect 12796 22482 12852 22540
rect 12796 22430 12798 22482
rect 12850 22430 12852 22482
rect 12796 22418 12852 22430
rect 13132 22484 13188 24444
rect 13244 24434 13300 24444
rect 13356 23380 13412 26852
rect 13692 25172 13748 38612
rect 13916 37828 13972 45836
rect 14028 45108 14084 45118
rect 14028 45014 14084 45052
rect 14140 43428 14196 45948
rect 14252 43652 14308 46398
rect 14364 45332 14420 45342
rect 14364 45238 14420 45276
rect 14476 44436 14532 48300
rect 14588 48354 14644 49644
rect 14700 49028 14756 49756
rect 14812 49810 14868 49822
rect 14812 49758 14814 49810
rect 14866 49758 14868 49810
rect 14812 49252 14868 49758
rect 14924 49812 14980 50652
rect 15372 50484 15428 50522
rect 15372 50418 15428 50428
rect 15596 50482 15652 50494
rect 15596 50430 15598 50482
rect 15650 50430 15652 50482
rect 14924 49746 14980 49756
rect 15260 49812 15316 49822
rect 15260 49810 15540 49812
rect 15260 49758 15262 49810
rect 15314 49758 15540 49810
rect 15260 49756 15540 49758
rect 15260 49746 15316 49756
rect 14812 49186 14868 49196
rect 15260 49588 15316 49598
rect 15260 49138 15316 49532
rect 15260 49086 15262 49138
rect 15314 49086 15316 49138
rect 15260 49074 15316 49086
rect 14700 48962 14756 48972
rect 14588 48302 14590 48354
rect 14642 48302 14644 48354
rect 14588 48290 14644 48302
rect 14924 48804 14980 48814
rect 14700 48244 14756 48254
rect 14700 48018 14756 48188
rect 14700 47966 14702 48018
rect 14754 47966 14756 48018
rect 14700 47682 14756 47966
rect 14700 47630 14702 47682
rect 14754 47630 14756 47682
rect 14700 47618 14756 47630
rect 14812 47796 14868 47806
rect 14812 47570 14868 47740
rect 14812 47518 14814 47570
rect 14866 47518 14868 47570
rect 14812 47506 14868 47518
rect 14924 47124 14980 48748
rect 15372 48244 15428 48254
rect 15372 48150 15428 48188
rect 15484 47570 15540 49756
rect 15596 49364 15652 50430
rect 15708 50482 15764 51436
rect 15932 51268 15988 51278
rect 16156 51268 16212 57484
rect 16940 56978 16996 57932
rect 17612 57874 17668 58156
rect 17612 57822 17614 57874
rect 17666 57822 17668 57874
rect 17612 57810 17668 57822
rect 17388 57764 17444 57774
rect 17388 57670 17444 57708
rect 16940 56926 16942 56978
rect 16994 56926 16996 56978
rect 16940 56914 16996 56926
rect 17164 56866 17220 56878
rect 17164 56814 17166 56866
rect 17218 56814 17220 56866
rect 16604 56642 16660 56654
rect 16604 56590 16606 56642
rect 16658 56590 16660 56642
rect 16604 56532 16660 56590
rect 16604 56466 16660 56476
rect 17164 56532 17220 56814
rect 17164 56466 17220 56476
rect 17500 56642 17556 56654
rect 17500 56590 17502 56642
rect 17554 56590 17556 56642
rect 17500 56194 17556 56590
rect 17500 56142 17502 56194
rect 17554 56142 17556 56194
rect 17500 56130 17556 56142
rect 16716 55076 16772 55086
rect 16716 53730 16772 55020
rect 16716 53678 16718 53730
rect 16770 53678 16772 53730
rect 16380 53506 16436 53518
rect 16380 53454 16382 53506
rect 16434 53454 16436 53506
rect 16268 53172 16324 53182
rect 16268 53078 16324 53116
rect 16268 52724 16324 52734
rect 16268 52162 16324 52668
rect 16380 52612 16436 53454
rect 16604 53060 16660 53070
rect 16604 52966 16660 53004
rect 16380 52546 16436 52556
rect 16268 52110 16270 52162
rect 16322 52110 16324 52162
rect 16268 52098 16324 52110
rect 16604 51604 16660 51614
rect 16380 51380 16436 51390
rect 16380 51286 16436 51324
rect 15932 51266 16212 51268
rect 15932 51214 15934 51266
rect 15986 51214 16212 51266
rect 15932 51212 16212 51214
rect 15932 51202 15988 51212
rect 15708 50430 15710 50482
rect 15762 50430 15764 50482
rect 15708 50418 15764 50430
rect 16044 50428 16100 51212
rect 16268 50932 16324 50942
rect 15932 50372 15988 50382
rect 16044 50372 16212 50428
rect 15932 50278 15988 50316
rect 15596 49298 15652 49308
rect 15932 49810 15988 49822
rect 15932 49758 15934 49810
rect 15986 49758 15988 49810
rect 15932 49028 15988 49758
rect 16156 49700 16212 50372
rect 16268 49922 16324 50876
rect 16604 50706 16660 51548
rect 16716 51380 16772 53678
rect 16828 54516 16884 54526
rect 17388 54516 17444 54526
rect 16828 54514 17444 54516
rect 16828 54462 16830 54514
rect 16882 54462 17390 54514
rect 17442 54462 17444 54514
rect 16828 54460 17444 54462
rect 16828 53732 16884 54460
rect 17388 54450 17444 54460
rect 17724 54180 17780 60284
rect 17836 60274 17892 60284
rect 17836 58660 17892 58670
rect 17836 58434 17892 58604
rect 17836 58382 17838 58434
rect 17890 58382 17892 58434
rect 17836 58370 17892 58382
rect 17836 58100 17892 58110
rect 17836 57874 17892 58044
rect 17836 57822 17838 57874
rect 17890 57822 17892 57874
rect 17836 56980 17892 57822
rect 17948 57652 18004 61292
rect 18172 59778 18228 59790
rect 18172 59726 18174 59778
rect 18226 59726 18228 59778
rect 18060 59218 18116 59230
rect 18060 59166 18062 59218
rect 18114 59166 18116 59218
rect 18060 57874 18116 59166
rect 18172 59220 18228 59726
rect 18172 59154 18228 59164
rect 18060 57822 18062 57874
rect 18114 57822 18116 57874
rect 18060 57810 18116 57822
rect 18060 57652 18116 57662
rect 17948 57650 18116 57652
rect 17948 57598 18062 57650
rect 18114 57598 18116 57650
rect 17948 57596 18116 57598
rect 17948 56980 18004 56990
rect 17836 56924 17948 56980
rect 17948 56886 18004 56924
rect 18060 56420 18116 57596
rect 18508 57428 18564 64430
rect 18620 64484 18676 64494
rect 18620 63250 18676 64428
rect 18620 63198 18622 63250
rect 18674 63198 18676 63250
rect 18620 63186 18676 63198
rect 18620 62580 18676 62590
rect 18620 62486 18676 62524
rect 18732 62132 18788 66332
rect 18844 66052 18900 67228
rect 18956 67060 19012 67070
rect 18956 66274 19012 67004
rect 19292 67058 19348 67070
rect 19292 67006 19294 67058
rect 19346 67006 19348 67058
rect 18956 66222 18958 66274
rect 19010 66222 19012 66274
rect 18956 66210 19012 66222
rect 19068 66834 19124 66846
rect 19068 66782 19070 66834
rect 19122 66782 19124 66834
rect 18844 65996 19012 66052
rect 18732 60676 18788 62076
rect 18732 60114 18788 60620
rect 18732 60062 18734 60114
rect 18786 60062 18788 60114
rect 18732 59668 18788 60062
rect 18620 59612 18788 59668
rect 18844 65828 18900 65838
rect 18620 58884 18676 59612
rect 18844 59556 18900 65772
rect 18956 63140 19012 65996
rect 19068 65490 19124 66782
rect 19180 66500 19236 66510
rect 19180 66406 19236 66444
rect 19292 66276 19348 67006
rect 19404 66500 19460 67564
rect 19404 66434 19460 66444
rect 19628 67618 19684 67630
rect 19628 67566 19630 67618
rect 19682 67566 19684 67618
rect 19292 66210 19348 66220
rect 19404 66276 19460 66286
rect 19628 66276 19684 67566
rect 19836 67452 20100 67462
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 19836 67386 20100 67396
rect 20076 67172 20132 67182
rect 20076 67058 20132 67116
rect 20076 67006 20078 67058
rect 20130 67006 20132 67058
rect 20076 66994 20132 67006
rect 19404 66274 19684 66276
rect 19404 66222 19406 66274
rect 19458 66222 19684 66274
rect 19404 66220 19684 66222
rect 20412 66276 20468 66286
rect 19068 65438 19070 65490
rect 19122 65438 19124 65490
rect 19068 65426 19124 65438
rect 18956 62580 19012 63084
rect 19180 65378 19236 65390
rect 19180 65326 19182 65378
rect 19234 65326 19236 65378
rect 19068 62580 19124 62590
rect 19012 62578 19124 62580
rect 19012 62526 19070 62578
rect 19122 62526 19124 62578
rect 19012 62524 19124 62526
rect 18956 62486 19012 62524
rect 19068 62514 19124 62524
rect 19180 62188 19236 65326
rect 19404 65380 19460 66220
rect 19836 65884 20100 65894
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 19836 65818 20100 65828
rect 19404 65314 19460 65324
rect 19516 65716 19572 65726
rect 19516 64594 19572 65660
rect 19516 64542 19518 64594
rect 19570 64542 19572 64594
rect 19516 64530 19572 64542
rect 19836 64316 20100 64326
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 19836 64250 20100 64260
rect 19964 64036 20020 64046
rect 19964 63942 20020 63980
rect 19628 63810 19684 63822
rect 19628 63758 19630 63810
rect 19682 63758 19684 63810
rect 19404 62580 19460 62590
rect 19404 62354 19460 62524
rect 19404 62302 19406 62354
rect 19458 62302 19460 62354
rect 19404 62290 19460 62302
rect 19180 62132 19348 62188
rect 18956 61572 19012 61582
rect 18956 61012 19012 61516
rect 18956 60918 19012 60956
rect 18732 59500 18900 59556
rect 18956 60788 19012 60798
rect 18956 60002 19012 60732
rect 19180 60786 19236 60798
rect 19180 60734 19182 60786
rect 19234 60734 19236 60786
rect 18956 59950 18958 60002
rect 19010 59950 19012 60002
rect 18732 59444 18788 59500
rect 18956 59444 19012 59950
rect 18732 59350 18788 59388
rect 18844 59388 19012 59444
rect 19068 60226 19124 60238
rect 19068 60174 19070 60226
rect 19122 60174 19124 60226
rect 18620 58828 18788 58884
rect 18620 58660 18676 58670
rect 18620 58546 18676 58604
rect 18620 58494 18622 58546
rect 18674 58494 18676 58546
rect 18620 58482 18676 58494
rect 18508 57362 18564 57372
rect 18060 56354 18116 56364
rect 18284 57204 18340 57214
rect 18284 56866 18340 57148
rect 18396 56980 18452 56990
rect 18452 56924 18564 56980
rect 18396 56914 18452 56924
rect 18284 56814 18286 56866
rect 18338 56814 18340 56866
rect 17836 56196 17892 56206
rect 17836 56194 18228 56196
rect 17836 56142 17838 56194
rect 17890 56142 18228 56194
rect 17836 56140 18228 56142
rect 17836 56130 17892 56140
rect 17276 54124 17780 54180
rect 17948 55972 18004 55982
rect 17948 55074 18004 55916
rect 17948 55022 17950 55074
rect 18002 55022 18004 55074
rect 17052 53844 17108 53854
rect 17052 53750 17108 53788
rect 16828 53666 16884 53676
rect 16828 52276 16884 52286
rect 16828 52182 16884 52220
rect 17164 52276 17220 52286
rect 16828 52052 16884 52062
rect 16828 51602 16884 51996
rect 16828 51550 16830 51602
rect 16882 51550 16884 51602
rect 16828 51538 16884 51550
rect 16716 51324 16884 51380
rect 16604 50654 16606 50706
rect 16658 50654 16660 50706
rect 16604 50642 16660 50654
rect 16716 51044 16772 51054
rect 16268 49870 16270 49922
rect 16322 49870 16324 49922
rect 16268 49858 16324 49870
rect 16492 49810 16548 49822
rect 16492 49758 16494 49810
rect 16546 49758 16548 49810
rect 16492 49700 16548 49758
rect 16156 49644 16548 49700
rect 16492 49364 16548 49644
rect 15932 48962 15988 48972
rect 16044 49140 16100 49150
rect 16044 49026 16100 49084
rect 16156 49140 16212 49150
rect 16156 49138 16436 49140
rect 16156 49086 16158 49138
rect 16210 49086 16436 49138
rect 16156 49084 16436 49086
rect 16156 49074 16212 49084
rect 16044 48974 16046 49026
rect 16098 48974 16100 49026
rect 16044 48962 16100 48974
rect 15484 47518 15486 47570
rect 15538 47518 15540 47570
rect 15484 47506 15540 47518
rect 15596 48914 15652 48926
rect 15596 48862 15598 48914
rect 15650 48862 15652 48914
rect 15596 47572 15652 48862
rect 15820 48804 15876 48814
rect 15820 48710 15876 48748
rect 16156 48802 16212 48814
rect 16156 48750 16158 48802
rect 16210 48750 16212 48802
rect 16156 48580 16212 48750
rect 16268 48580 16324 48590
rect 15596 47506 15652 47516
rect 15708 48524 16268 48580
rect 15708 47458 15764 48524
rect 16268 48514 16324 48524
rect 15820 48356 15876 48366
rect 15820 48130 15876 48300
rect 15820 48078 15822 48130
rect 15874 48078 15876 48130
rect 15820 47796 15876 48078
rect 15820 47730 15876 47740
rect 16156 48242 16212 48254
rect 16156 48190 16158 48242
rect 16210 48190 16212 48242
rect 15708 47406 15710 47458
rect 15762 47406 15764 47458
rect 15036 47348 15092 47358
rect 15036 47254 15092 47292
rect 15484 47348 15540 47358
rect 15484 47254 15540 47292
rect 15260 47234 15316 47246
rect 15260 47182 15262 47234
rect 15314 47182 15316 47234
rect 15260 47124 15316 47182
rect 15708 47236 15764 47406
rect 15708 47170 15764 47180
rect 14924 47068 15316 47124
rect 16156 47068 16212 48190
rect 16380 48242 16436 49084
rect 16492 48356 16548 49308
rect 16492 48290 16548 48300
rect 16380 48190 16382 48242
rect 16434 48190 16436 48242
rect 16380 48178 16436 48190
rect 16492 48130 16548 48142
rect 16492 48078 16494 48130
rect 16546 48078 16548 48130
rect 16492 47458 16548 48078
rect 16492 47406 16494 47458
rect 16546 47406 16548 47458
rect 16492 47394 16548 47406
rect 16268 47236 16324 47246
rect 16268 47142 16324 47180
rect 15036 46562 15092 47068
rect 16156 47012 16324 47068
rect 15036 46510 15038 46562
rect 15090 46510 15092 46562
rect 14812 45666 14868 45678
rect 14812 45614 14814 45666
rect 14866 45614 14868 45666
rect 14812 44994 14868 45614
rect 14812 44942 14814 44994
rect 14866 44942 14868 44994
rect 14476 44434 14644 44436
rect 14476 44382 14478 44434
rect 14530 44382 14644 44434
rect 14476 44380 14644 44382
rect 14476 44370 14532 44380
rect 14252 43596 14532 43652
rect 14252 43428 14308 43438
rect 14140 43426 14308 43428
rect 14140 43374 14254 43426
rect 14306 43374 14308 43426
rect 14140 43372 14308 43374
rect 14252 43362 14308 43372
rect 14364 42530 14420 42542
rect 14364 42478 14366 42530
rect 14418 42478 14420 42530
rect 14364 42308 14420 42478
rect 14364 42242 14420 42252
rect 14364 40516 14420 40526
rect 14364 40422 14420 40460
rect 14028 39396 14084 39406
rect 14028 39302 14084 39340
rect 14476 38668 14532 43596
rect 14588 41972 14644 44380
rect 14812 42530 14868 44942
rect 15036 42644 15092 46510
rect 15596 46564 15652 46574
rect 15596 46470 15652 46508
rect 15932 46562 15988 46574
rect 15932 46510 15934 46562
rect 15986 46510 15988 46562
rect 15932 46340 15988 46510
rect 16268 46564 16324 47012
rect 15932 46274 15988 46284
rect 16044 46450 16100 46462
rect 16044 46398 16046 46450
rect 16098 46398 16100 46450
rect 15932 45892 15988 45902
rect 16044 45892 16100 46398
rect 15932 45890 16100 45892
rect 15932 45838 15934 45890
rect 15986 45838 16100 45890
rect 15932 45836 16100 45838
rect 15932 45826 15988 45836
rect 16156 45778 16212 45790
rect 16156 45726 16158 45778
rect 16210 45726 16212 45778
rect 15148 45666 15204 45678
rect 15148 45614 15150 45666
rect 15202 45614 15204 45666
rect 15148 45332 15204 45614
rect 15596 45668 15652 45678
rect 15596 45666 15764 45668
rect 15596 45614 15598 45666
rect 15650 45614 15764 45666
rect 15596 45612 15764 45614
rect 15596 45602 15652 45612
rect 15148 44996 15204 45276
rect 15372 45108 15428 45118
rect 15372 45014 15428 45052
rect 15260 44996 15316 45006
rect 15148 44994 15316 44996
rect 15148 44942 15262 44994
rect 15314 44942 15316 44994
rect 15148 44940 15316 44942
rect 15148 44100 15204 44940
rect 15260 44930 15316 44940
rect 15260 44212 15316 44222
rect 15260 44100 15316 44156
rect 15596 44100 15652 44110
rect 15148 44098 15540 44100
rect 15148 44046 15150 44098
rect 15202 44046 15540 44098
rect 15148 44044 15540 44046
rect 15148 44034 15204 44044
rect 15148 43652 15204 43662
rect 15148 43538 15204 43596
rect 15148 43486 15150 43538
rect 15202 43486 15204 43538
rect 15148 43474 15204 43486
rect 15484 43540 15540 44044
rect 15596 44006 15652 44044
rect 15484 43484 15652 43540
rect 15372 43314 15428 43326
rect 15372 43262 15374 43314
rect 15426 43262 15428 43314
rect 15372 43204 15428 43262
rect 15372 43138 15428 43148
rect 15484 43316 15540 43326
rect 15148 42756 15204 42766
rect 15148 42754 15316 42756
rect 15148 42702 15150 42754
rect 15202 42702 15316 42754
rect 15148 42700 15316 42702
rect 15148 42690 15204 42700
rect 15036 42578 15092 42588
rect 14812 42478 14814 42530
rect 14866 42478 14868 42530
rect 14812 42196 14868 42478
rect 14812 42130 14868 42140
rect 14588 41906 14644 41916
rect 15036 41860 15092 41870
rect 15036 41766 15092 41804
rect 15148 41300 15204 41310
rect 14812 41188 14868 41198
rect 15036 41188 15092 41198
rect 14812 41094 14868 41132
rect 14924 41186 15092 41188
rect 14924 41134 15038 41186
rect 15090 41134 15092 41186
rect 14924 41132 15092 41134
rect 14924 40292 14980 41132
rect 15036 41122 15092 41132
rect 15148 40516 15204 41244
rect 14924 40226 14980 40236
rect 15036 40514 15204 40516
rect 15036 40462 15150 40514
rect 15202 40462 15204 40514
rect 15036 40460 15204 40462
rect 15036 39506 15092 40460
rect 15148 40422 15204 40460
rect 15148 39620 15204 39630
rect 15148 39526 15204 39564
rect 15036 39454 15038 39506
rect 15090 39454 15092 39506
rect 15036 39442 15092 39454
rect 14924 39396 14980 39406
rect 14924 39302 14980 39340
rect 14364 38612 14532 38668
rect 15036 39284 15092 39294
rect 14252 37828 14308 37838
rect 13916 37734 13972 37772
rect 14028 37826 14308 37828
rect 14028 37774 14254 37826
rect 14306 37774 14308 37826
rect 14028 37772 14308 37774
rect 14028 37492 14084 37772
rect 14252 37762 14308 37772
rect 13804 37436 14084 37492
rect 13804 37378 13860 37436
rect 13804 37326 13806 37378
rect 13858 37326 13860 37378
rect 13804 37314 13860 37326
rect 13804 30436 13860 30446
rect 13804 29652 13860 30380
rect 13804 28866 13860 29596
rect 14252 29876 14308 29886
rect 13804 28814 13806 28866
rect 13858 28814 13860 28866
rect 13804 28802 13860 28814
rect 14140 29428 14196 29438
rect 14028 28756 14084 28766
rect 14028 28662 14084 28700
rect 14140 28644 14196 29372
rect 14140 28578 14196 28588
rect 14252 28420 14308 29820
rect 13692 25106 13748 25116
rect 14028 28364 14308 28420
rect 14028 24948 14084 28364
rect 14364 26908 14420 38612
rect 14812 38164 14868 38174
rect 14812 38070 14868 38108
rect 14588 38050 14644 38062
rect 14588 37998 14590 38050
rect 14642 37998 14644 38050
rect 14588 37828 14644 37998
rect 14588 35140 14644 37772
rect 14924 35586 14980 35598
rect 14924 35534 14926 35586
rect 14978 35534 14980 35586
rect 14924 35476 14980 35534
rect 14924 35410 14980 35420
rect 15036 35308 15092 39228
rect 15260 38668 15316 42700
rect 15372 42644 15428 42654
rect 15484 42644 15540 43260
rect 15372 42642 15540 42644
rect 15372 42590 15374 42642
rect 15426 42590 15540 42642
rect 15372 42588 15540 42590
rect 15372 42578 15428 42588
rect 15596 42308 15652 43484
rect 15708 42868 15764 45612
rect 16044 45556 16100 45566
rect 15932 45500 16044 45556
rect 15932 44322 15988 45500
rect 16044 45490 16100 45500
rect 15932 44270 15934 44322
rect 15986 44270 15988 44322
rect 15932 44212 15988 44270
rect 15932 44146 15988 44156
rect 16156 43540 16212 45726
rect 16268 45668 16324 46508
rect 16492 46562 16548 46574
rect 16492 46510 16494 46562
rect 16546 46510 16548 46562
rect 16380 46004 16436 46014
rect 16380 45890 16436 45948
rect 16380 45838 16382 45890
rect 16434 45838 16436 45890
rect 16380 45826 16436 45838
rect 16492 45892 16548 46510
rect 16716 46450 16772 50988
rect 16828 49588 16884 51324
rect 17164 50428 17220 52220
rect 17276 52276 17332 54124
rect 17836 53618 17892 53630
rect 17836 53566 17838 53618
rect 17890 53566 17892 53618
rect 17836 53508 17892 53566
rect 17836 53442 17892 53452
rect 17500 53058 17556 53070
rect 17500 53006 17502 53058
rect 17554 53006 17556 53058
rect 17388 52724 17444 52734
rect 17388 52630 17444 52668
rect 17500 52612 17556 53006
rect 17724 52724 17780 52734
rect 17948 52724 18004 55022
rect 18172 54626 18228 56140
rect 18172 54574 18174 54626
rect 18226 54574 18228 54626
rect 18172 54562 18228 54574
rect 18172 53508 18228 53518
rect 17780 52668 18004 52724
rect 18060 52948 18116 52958
rect 17724 52630 17780 52668
rect 17500 52546 17556 52556
rect 18060 52276 18116 52892
rect 17276 52274 17668 52276
rect 17276 52222 17278 52274
rect 17330 52222 17668 52274
rect 17276 52220 17668 52222
rect 17276 52210 17332 52220
rect 17612 50484 17668 52220
rect 17052 50370 17108 50382
rect 17164 50372 17444 50428
rect 17052 50318 17054 50370
rect 17106 50318 17108 50370
rect 17052 50036 17108 50318
rect 17052 49970 17108 49980
rect 16828 49522 16884 49532
rect 17052 48802 17108 48814
rect 17052 48750 17054 48802
rect 17106 48750 17108 48802
rect 17052 48692 17108 48750
rect 17052 48626 17108 48636
rect 17388 48468 17444 50372
rect 17612 49924 17668 50428
rect 17612 49858 17668 49868
rect 17724 52162 17780 52174
rect 17724 52110 17726 52162
rect 17778 52110 17780 52162
rect 17724 50596 17780 52110
rect 17948 52052 18004 52062
rect 17836 51716 17892 51726
rect 17836 51602 17892 51660
rect 17836 51550 17838 51602
rect 17890 51550 17892 51602
rect 17836 51538 17892 51550
rect 17948 51492 18004 51996
rect 18060 52050 18116 52220
rect 18060 51998 18062 52050
rect 18114 51998 18116 52050
rect 18060 51986 18116 51998
rect 18172 51604 18228 53452
rect 18284 53060 18340 56814
rect 18508 56866 18564 56924
rect 18508 56814 18510 56866
rect 18562 56814 18564 56866
rect 18508 56532 18564 56814
rect 18508 56466 18564 56476
rect 18508 56196 18564 56206
rect 18508 56102 18564 56140
rect 18732 55972 18788 58828
rect 18844 57092 18900 59388
rect 18956 59220 19012 59230
rect 19068 59220 19124 60174
rect 18956 59218 19124 59220
rect 18956 59166 18958 59218
rect 19010 59166 19124 59218
rect 18956 59164 19124 59166
rect 18956 59154 19012 59164
rect 19180 58660 19236 60734
rect 19180 58594 19236 58604
rect 18844 57026 18900 57036
rect 19180 57762 19236 57774
rect 19180 57710 19182 57762
rect 19234 57710 19236 57762
rect 18844 56868 18900 56878
rect 18844 56644 18900 56812
rect 19180 56868 19236 57710
rect 19292 57092 19348 62132
rect 19516 62132 19572 62142
rect 19516 62038 19572 62076
rect 19404 61348 19460 61358
rect 19404 60898 19460 61292
rect 19404 60846 19406 60898
rect 19458 60846 19460 60898
rect 19404 60002 19460 60846
rect 19516 61012 19572 61022
rect 19516 60898 19572 60956
rect 19516 60846 19518 60898
rect 19570 60846 19572 60898
rect 19516 60834 19572 60846
rect 19404 59950 19406 60002
rect 19458 59950 19460 60002
rect 19404 59938 19460 59950
rect 19516 59332 19572 59342
rect 19516 59238 19572 59276
rect 19292 57026 19348 57036
rect 19404 59108 19460 59118
rect 19404 57204 19460 59052
rect 19180 56802 19236 56812
rect 19292 56868 19348 56878
rect 19404 56868 19460 57148
rect 19292 56866 19460 56868
rect 19292 56814 19294 56866
rect 19346 56814 19460 56866
rect 19292 56812 19460 56814
rect 19292 56802 19348 56812
rect 18844 56642 19012 56644
rect 18844 56590 18846 56642
rect 18898 56590 19012 56642
rect 18844 56588 19012 56590
rect 18844 56578 18900 56588
rect 18732 55906 18788 55916
rect 18508 55074 18564 55086
rect 18508 55022 18510 55074
rect 18562 55022 18564 55074
rect 18508 53956 18564 55022
rect 18508 53890 18564 53900
rect 18844 53170 18900 53182
rect 18844 53118 18846 53170
rect 18898 53118 18900 53170
rect 18508 53060 18564 53070
rect 18284 53058 18564 53060
rect 18284 53006 18510 53058
rect 18562 53006 18564 53058
rect 18284 53004 18564 53006
rect 18172 51538 18228 51548
rect 18284 52836 18340 52846
rect 18060 51492 18116 51502
rect 17948 51490 18116 51492
rect 17948 51438 18062 51490
rect 18114 51438 18116 51490
rect 17948 51436 18116 51438
rect 18060 51380 18116 51436
rect 18060 51324 18228 51380
rect 17500 49810 17556 49822
rect 17500 49758 17502 49810
rect 17554 49758 17556 49810
rect 17500 49588 17556 49758
rect 17500 49522 17556 49532
rect 17612 48916 17668 48926
rect 17724 48916 17780 50540
rect 18060 50482 18116 50494
rect 18060 50430 18062 50482
rect 18114 50430 18116 50482
rect 18060 50034 18116 50430
rect 18060 49982 18062 50034
rect 18114 49982 18116 50034
rect 17612 48914 17780 48916
rect 17612 48862 17614 48914
rect 17666 48862 17780 48914
rect 17612 48860 17780 48862
rect 17836 49812 17892 49822
rect 17836 49476 17892 49756
rect 17612 48850 17668 48860
rect 17388 48242 17444 48412
rect 17388 48190 17390 48242
rect 17442 48190 17444 48242
rect 17052 47346 17108 47358
rect 17052 47294 17054 47346
rect 17106 47294 17108 47346
rect 16716 46398 16718 46450
rect 16770 46398 16772 46450
rect 16716 46386 16772 46398
rect 16828 46562 16884 46574
rect 16828 46510 16830 46562
rect 16882 46510 16884 46562
rect 16828 46004 16884 46510
rect 16492 45826 16548 45836
rect 16716 45948 16884 46004
rect 16268 45612 16548 45668
rect 16156 43446 16212 43484
rect 16268 44884 16324 44894
rect 15820 43316 15876 43326
rect 15820 43314 16212 43316
rect 15820 43262 15822 43314
rect 15874 43262 16212 43314
rect 15820 43260 16212 43262
rect 15820 43250 15876 43260
rect 15708 42812 16100 42868
rect 15932 42642 15988 42654
rect 15932 42590 15934 42642
rect 15986 42590 15988 42642
rect 15932 42308 15988 42590
rect 15596 42252 15764 42308
rect 15484 42196 15540 42206
rect 15484 42102 15540 42140
rect 15708 42084 15764 42252
rect 15932 42242 15988 42252
rect 15932 42084 15988 42094
rect 15708 42082 15988 42084
rect 15708 42030 15934 42082
rect 15986 42030 15988 42082
rect 15708 42028 15988 42030
rect 15932 42018 15988 42028
rect 15372 41412 15428 41422
rect 15372 40628 15428 41356
rect 15596 41084 15652 41096
rect 15596 41032 15598 41084
rect 15650 41076 15652 41084
rect 15708 41076 15764 41086
rect 15650 41032 15708 41076
rect 15596 41020 15708 41032
rect 15708 41010 15764 41020
rect 15372 40290 15428 40572
rect 15372 40238 15374 40290
rect 15426 40238 15428 40290
rect 15372 40226 15428 40238
rect 15596 40404 15652 40414
rect 15596 39842 15652 40348
rect 15932 40404 15988 40414
rect 15708 40180 15764 40190
rect 15708 40086 15764 40124
rect 15596 39790 15598 39842
rect 15650 39790 15652 39842
rect 15596 39778 15652 39790
rect 15932 38836 15988 40348
rect 15932 38770 15988 38780
rect 15484 38722 15540 38734
rect 15484 38670 15486 38722
rect 15538 38670 15540 38722
rect 15484 38668 15540 38670
rect 15260 38612 15428 38668
rect 15484 38612 15764 38668
rect 15260 38276 15316 38286
rect 15260 37940 15316 38220
rect 15372 38164 15428 38612
rect 15372 38108 15540 38164
rect 15372 37940 15428 37950
rect 15260 37938 15428 37940
rect 15260 37886 15374 37938
rect 15426 37886 15428 37938
rect 15260 37884 15428 37886
rect 15372 37492 15428 37884
rect 15372 37426 15428 37436
rect 15148 36596 15204 36606
rect 15148 36502 15204 36540
rect 15372 35476 15428 35486
rect 15036 35252 15316 35308
rect 14588 35084 15204 35140
rect 15148 34914 15204 35084
rect 15148 34862 15150 34914
rect 15202 34862 15204 34914
rect 14812 34692 14868 34702
rect 15148 34692 15204 34862
rect 14812 34690 15092 34692
rect 14812 34638 14814 34690
rect 14866 34638 15092 34690
rect 14812 34636 15092 34638
rect 14812 34626 14868 34636
rect 15036 34242 15092 34636
rect 15148 34626 15204 34636
rect 15036 34190 15038 34242
rect 15090 34190 15092 34242
rect 15036 34178 15092 34190
rect 15260 33684 15316 35252
rect 15372 35026 15428 35420
rect 15484 35308 15540 38108
rect 15596 37828 15652 37838
rect 15596 35924 15652 37772
rect 15708 37490 15764 38612
rect 15932 38164 15988 38174
rect 15932 38070 15988 38108
rect 15820 38052 15876 38062
rect 15820 37958 15876 37996
rect 15932 37828 15988 37838
rect 15708 37438 15710 37490
rect 15762 37438 15764 37490
rect 15708 37426 15764 37438
rect 15820 37772 15932 37828
rect 15820 36148 15876 37772
rect 15932 37734 15988 37772
rect 16044 37604 16100 42812
rect 16156 39508 16212 43260
rect 16268 42866 16324 44828
rect 16380 44212 16436 44222
rect 16380 43650 16436 44156
rect 16380 43598 16382 43650
rect 16434 43598 16436 43650
rect 16380 43586 16436 43598
rect 16268 42814 16270 42866
rect 16322 42814 16324 42866
rect 16268 42802 16324 42814
rect 16380 43092 16436 43102
rect 16380 42194 16436 43036
rect 16380 42142 16382 42194
rect 16434 42142 16436 42194
rect 16380 42130 16436 42142
rect 16380 41188 16436 41198
rect 16380 40740 16436 41132
rect 16492 41086 16548 45612
rect 16716 45108 16772 45948
rect 16716 44324 16772 45052
rect 16828 45778 16884 45790
rect 16828 45726 16830 45778
rect 16882 45726 16884 45778
rect 16828 44996 16884 45726
rect 16940 45668 16996 45678
rect 16940 45574 16996 45612
rect 16828 44902 16884 44940
rect 17052 44884 17108 47294
rect 17052 44818 17108 44828
rect 17164 47236 17220 47246
rect 16716 44268 16884 44324
rect 16716 44100 16772 44110
rect 16716 43538 16772 44044
rect 16716 43486 16718 43538
rect 16770 43486 16772 43538
rect 16716 43092 16772 43486
rect 16716 43026 16772 43036
rect 16828 43428 16884 44268
rect 17052 44212 17108 44222
rect 17052 44118 17108 44156
rect 16716 42532 16772 42542
rect 16716 42438 16772 42476
rect 16828 42194 16884 43372
rect 16828 42142 16830 42194
rect 16882 42142 16884 42194
rect 16828 42130 16884 42142
rect 16940 43652 16996 43662
rect 16940 43538 16996 43596
rect 16940 43486 16942 43538
rect 16994 43486 16996 43538
rect 16940 42196 16996 43486
rect 16940 42130 16996 42140
rect 16940 41972 16996 41982
rect 16492 41030 16660 41086
rect 16380 40626 16436 40684
rect 16380 40574 16382 40626
rect 16434 40574 16436 40626
rect 16380 40562 16436 40574
rect 16492 40962 16548 40974
rect 16492 40910 16494 40962
rect 16546 40910 16548 40962
rect 16492 40852 16548 40910
rect 16156 39442 16212 39452
rect 16268 40516 16324 40526
rect 16268 38834 16324 40460
rect 16492 40516 16548 40796
rect 16492 40450 16548 40460
rect 16268 38782 16270 38834
rect 16322 38782 16324 38834
rect 16268 38668 16324 38782
rect 16156 38612 16324 38668
rect 16380 39394 16436 39406
rect 16380 39342 16382 39394
rect 16434 39342 16436 39394
rect 16380 38612 16436 39342
rect 16156 37716 16212 38612
rect 16380 38546 16436 38556
rect 16492 38836 16548 38846
rect 16492 38388 16548 38780
rect 16156 37650 16212 37660
rect 16268 38332 16548 38388
rect 15932 37548 16100 37604
rect 15932 36932 15988 37548
rect 16044 37380 16100 37390
rect 16268 37380 16324 38332
rect 16604 38276 16660 41030
rect 16940 40626 16996 41916
rect 17052 40964 17108 40974
rect 17052 40870 17108 40908
rect 16940 40574 16942 40626
rect 16994 40574 16996 40626
rect 16940 40562 16996 40574
rect 16828 40516 16884 40526
rect 16828 40404 16884 40460
rect 16828 40348 16996 40404
rect 16828 38724 16884 38762
rect 16828 38500 16884 38668
rect 16828 38434 16884 38444
rect 16492 38220 16660 38276
rect 16380 38164 16436 38174
rect 16380 38070 16436 38108
rect 16044 37378 16324 37380
rect 16044 37326 16046 37378
rect 16098 37326 16324 37378
rect 16044 37324 16324 37326
rect 16044 37314 16100 37324
rect 15932 36876 16436 36932
rect 15820 36092 16212 36148
rect 15708 35924 15764 35934
rect 15596 35922 16100 35924
rect 15596 35870 15710 35922
rect 15762 35870 16100 35922
rect 15596 35868 16100 35870
rect 15708 35858 15764 35868
rect 15596 35700 15652 35710
rect 15596 35606 15652 35644
rect 15932 35698 15988 35710
rect 15932 35646 15934 35698
rect 15986 35646 15988 35698
rect 15820 35588 15876 35598
rect 15820 35494 15876 35532
rect 15932 35476 15988 35646
rect 15932 35410 15988 35420
rect 15484 35252 15764 35308
rect 15372 34974 15374 35026
rect 15426 34974 15428 35026
rect 15372 34962 15428 34974
rect 15148 33628 15316 33684
rect 15372 34242 15428 34254
rect 15372 34190 15374 34242
rect 15426 34190 15428 34242
rect 14588 33346 14644 33358
rect 14588 33294 14590 33346
rect 14642 33294 14644 33346
rect 14588 32900 14644 33294
rect 14812 32900 14868 32910
rect 14588 32844 14812 32900
rect 14700 32452 14756 32462
rect 14700 32358 14756 32396
rect 14700 29428 14756 29438
rect 14812 29428 14868 32844
rect 15148 32788 15204 33628
rect 15260 33460 15316 33470
rect 15372 33460 15428 34190
rect 15260 33458 15428 33460
rect 15260 33406 15262 33458
rect 15314 33406 15428 33458
rect 15260 33404 15428 33406
rect 15260 33394 15316 33404
rect 15596 32788 15652 32798
rect 15148 32732 15428 32788
rect 15148 32564 15204 32574
rect 15148 29876 15204 32508
rect 15260 31668 15316 31678
rect 15260 31574 15316 31612
rect 15148 29810 15204 29820
rect 14756 29372 14868 29428
rect 14700 29334 14756 29372
rect 13804 24946 14084 24948
rect 13804 24894 14030 24946
rect 14082 24894 14084 24946
rect 13804 24892 14084 24894
rect 13580 24498 13636 24510
rect 13580 24446 13582 24498
rect 13634 24446 13636 24498
rect 13580 23938 13636 24446
rect 13580 23886 13582 23938
rect 13634 23886 13636 23938
rect 13580 23874 13636 23886
rect 13132 20804 13188 22428
rect 13132 20738 13188 20748
rect 13244 23324 13412 23380
rect 12572 17444 12628 17454
rect 12572 16994 12628 17388
rect 12572 16942 12574 16994
rect 12626 16942 12628 16994
rect 12572 16930 12628 16942
rect 12236 16706 12292 16716
rect 12124 16146 12180 16156
rect 12908 16212 12964 16222
rect 12908 16118 12964 16156
rect 12012 16100 12068 16110
rect 11900 16044 12012 16100
rect 11788 15988 11844 15998
rect 11788 15894 11844 15932
rect 11676 15486 11678 15538
rect 11730 15486 11732 15538
rect 11676 15316 11732 15486
rect 10556 15092 11508 15148
rect 10444 13076 10500 13086
rect 10444 13074 10724 13076
rect 10444 13022 10446 13074
rect 10498 13022 10724 13074
rect 10444 13020 10724 13022
rect 10444 13010 10500 13020
rect 10668 10834 10724 13020
rect 10892 12740 10948 12750
rect 10780 12738 10948 12740
rect 10780 12686 10894 12738
rect 10946 12686 10948 12738
rect 10780 12684 10948 12686
rect 10780 11732 10836 12684
rect 10892 12674 10948 12684
rect 11340 12404 11396 12414
rect 11004 11844 11060 11854
rect 10780 11666 10836 11676
rect 10892 11788 11004 11844
rect 10668 10782 10670 10834
rect 10722 10782 10724 10834
rect 10668 10724 10724 10782
rect 10780 10836 10836 10846
rect 10780 10742 10836 10780
rect 10668 10658 10724 10668
rect 10444 10612 10500 10622
rect 10444 10610 10612 10612
rect 10444 10558 10446 10610
rect 10498 10558 10612 10610
rect 10444 10556 10612 10558
rect 10444 10546 10500 10556
rect 10444 10388 10500 10398
rect 10444 9826 10500 10332
rect 10556 9940 10612 10556
rect 10668 10498 10724 10510
rect 10668 10446 10670 10498
rect 10722 10446 10724 10498
rect 10668 10388 10724 10446
rect 10892 10388 10948 11788
rect 11004 11778 11060 11788
rect 11340 10834 11396 12348
rect 11340 10782 11342 10834
rect 11394 10782 11396 10834
rect 10668 10332 10948 10388
rect 11004 10612 11060 10622
rect 10668 9940 10724 9950
rect 10556 9884 10668 9940
rect 10444 9774 10446 9826
rect 10498 9774 10500 9826
rect 10444 9762 10500 9774
rect 10668 9826 10724 9884
rect 11004 9938 11060 10556
rect 11340 10386 11396 10782
rect 11340 10334 11342 10386
rect 11394 10334 11396 10386
rect 11340 10322 11396 10334
rect 11340 10052 11396 10062
rect 11004 9886 11006 9938
rect 11058 9886 11060 9938
rect 11004 9874 11060 9886
rect 11116 10050 11396 10052
rect 11116 9998 11342 10050
rect 11394 9998 11396 10050
rect 11116 9996 11396 9998
rect 10668 9774 10670 9826
rect 10722 9774 10724 9826
rect 10668 9762 10724 9774
rect 11116 9826 11172 9996
rect 11340 9986 11396 9996
rect 11452 9828 11508 15092
rect 11676 11732 11732 15260
rect 12012 15148 12068 16044
rect 12460 16098 12516 16110
rect 12460 16046 12462 16098
rect 12514 16046 12516 16098
rect 12124 15874 12180 15886
rect 12124 15822 12126 15874
rect 12178 15822 12180 15874
rect 12124 15428 12180 15822
rect 12236 15876 12292 15886
rect 12236 15782 12292 15820
rect 12460 15652 12516 16046
rect 12684 15652 12740 15662
rect 12460 15596 12684 15652
rect 12124 15362 12180 15372
rect 12684 15538 12740 15596
rect 12684 15486 12686 15538
rect 12738 15486 12740 15538
rect 12012 15092 12292 15148
rect 12236 12404 12292 15092
rect 12236 12310 12292 12348
rect 11676 11666 11732 11676
rect 12012 12292 12068 12302
rect 11788 11508 11844 11518
rect 11788 10836 11844 11452
rect 12012 11506 12068 12236
rect 12460 12178 12516 12190
rect 12460 12126 12462 12178
rect 12514 12126 12516 12178
rect 12348 12066 12404 12078
rect 12348 12014 12350 12066
rect 12402 12014 12404 12066
rect 12012 11454 12014 11506
rect 12066 11454 12068 11506
rect 12012 11442 12068 11454
rect 12124 11732 12180 11742
rect 12124 11172 12180 11676
rect 12348 11620 12404 12014
rect 12348 11554 12404 11564
rect 12460 11396 12516 12126
rect 12684 12180 12740 15486
rect 13132 15316 13188 15326
rect 13132 15222 13188 15260
rect 13244 15148 13300 23324
rect 13468 23156 13524 23166
rect 13468 21588 13524 23100
rect 13804 22596 13860 24892
rect 14028 24882 14084 24892
rect 14252 26852 14420 26908
rect 15036 26964 15092 26974
rect 13916 23716 13972 23726
rect 13916 23714 14196 23716
rect 13916 23662 13918 23714
rect 13970 23662 14196 23714
rect 13916 23660 14196 23662
rect 13916 23650 13972 23660
rect 14140 23266 14196 23660
rect 14140 23214 14142 23266
rect 14194 23214 14196 23266
rect 14140 23202 14196 23214
rect 13804 22530 13860 22540
rect 13468 21522 13524 21532
rect 14140 21588 14196 21598
rect 14140 21494 14196 21532
rect 13692 21474 13748 21486
rect 13692 21422 13694 21474
rect 13746 21422 13748 21474
rect 13692 21252 13748 21422
rect 13692 20916 13748 21196
rect 13692 20850 13748 20860
rect 14252 19348 14308 26852
rect 15036 26514 15092 26908
rect 15036 26462 15038 26514
rect 15090 26462 15092 26514
rect 15036 26450 15092 26462
rect 14812 26292 14868 26302
rect 14812 26198 14868 26236
rect 15148 23492 15204 23502
rect 14924 22372 14980 22382
rect 14924 22278 14980 22316
rect 15148 22372 15204 23436
rect 15260 22372 15316 22382
rect 15204 22370 15316 22372
rect 15204 22318 15262 22370
rect 15314 22318 15316 22370
rect 15204 22316 15316 22318
rect 15148 22306 15204 22316
rect 15260 22306 15316 22316
rect 14252 19254 14308 19292
rect 13468 19236 13524 19246
rect 13468 17668 13524 19180
rect 15372 18340 15428 32732
rect 15596 32452 15652 32732
rect 15596 31890 15652 32396
rect 15596 31838 15598 31890
rect 15650 31838 15652 31890
rect 15596 31826 15652 31838
rect 15708 29650 15764 35252
rect 15820 34692 15876 34702
rect 15820 33684 15876 34636
rect 16044 33908 16100 35868
rect 16156 35698 16212 36092
rect 16156 35646 16158 35698
rect 16210 35646 16212 35698
rect 16156 34020 16212 35646
rect 16156 33954 16212 33964
rect 16044 33842 16100 33852
rect 15820 33618 15876 33628
rect 15820 31778 15876 31790
rect 15820 31726 15822 31778
rect 15874 31726 15876 31778
rect 15820 31668 15876 31726
rect 15820 31602 15876 31612
rect 16156 31554 16212 31566
rect 16156 31502 16158 31554
rect 16210 31502 16212 31554
rect 16156 31108 16212 31502
rect 16268 31108 16324 31118
rect 16156 31106 16324 31108
rect 16156 31054 16270 31106
rect 16322 31054 16324 31106
rect 16156 31052 16324 31054
rect 16268 31042 16324 31052
rect 15708 29598 15710 29650
rect 15762 29598 15764 29650
rect 15708 29586 15764 29598
rect 15820 30996 15876 31006
rect 15484 29540 15540 29550
rect 15484 29446 15540 29484
rect 15820 29426 15876 30940
rect 15932 30210 15988 30222
rect 15932 30158 15934 30210
rect 15986 30158 15988 30210
rect 15932 29876 15988 30158
rect 16380 29988 16436 36876
rect 16492 30100 16548 38220
rect 16604 37938 16660 37950
rect 16604 37886 16606 37938
rect 16658 37886 16660 37938
rect 16604 37828 16660 37886
rect 16604 37762 16660 37772
rect 16828 37938 16884 37950
rect 16828 37886 16830 37938
rect 16882 37886 16884 37938
rect 16716 37716 16772 37726
rect 16604 37492 16660 37502
rect 16604 37398 16660 37436
rect 16604 36596 16660 36606
rect 16716 36596 16772 37660
rect 16828 37492 16884 37886
rect 16828 37426 16884 37436
rect 16604 36594 16772 36596
rect 16604 36542 16606 36594
rect 16658 36542 16772 36594
rect 16604 36540 16772 36542
rect 16828 36596 16884 36606
rect 16604 36530 16660 36540
rect 16828 32900 16884 36540
rect 16828 32786 16884 32844
rect 16828 32734 16830 32786
rect 16882 32734 16884 32786
rect 16828 32722 16884 32734
rect 16604 31106 16660 31118
rect 16604 31054 16606 31106
rect 16658 31054 16660 31106
rect 16604 30324 16660 31054
rect 16716 30324 16772 30334
rect 16604 30322 16772 30324
rect 16604 30270 16718 30322
rect 16770 30270 16772 30322
rect 16604 30268 16772 30270
rect 16716 30258 16772 30268
rect 16492 30044 16772 30100
rect 16380 29932 16548 29988
rect 15932 29810 15988 29820
rect 15820 29374 15822 29426
rect 15874 29374 15876 29426
rect 15820 29362 15876 29374
rect 16268 29426 16324 29438
rect 16268 29374 16270 29426
rect 16322 29374 16324 29426
rect 16156 28532 16212 28542
rect 16156 27076 16212 28476
rect 16268 28084 16324 29374
rect 16268 28018 16324 28028
rect 16380 27860 16436 27870
rect 16268 27076 16324 27086
rect 16156 27020 16268 27076
rect 15596 26964 15652 27002
rect 16268 26982 16324 27020
rect 15596 26898 15652 26908
rect 15820 26292 15876 26302
rect 15820 26198 15876 26236
rect 15484 26178 15540 26190
rect 15484 26126 15486 26178
rect 15538 26126 15540 26178
rect 15484 26068 15540 26126
rect 16380 26180 16436 27804
rect 16492 26292 16548 29932
rect 16604 29652 16660 29662
rect 16604 29558 16660 29596
rect 16604 27858 16660 27870
rect 16604 27806 16606 27858
rect 16658 27806 16660 27858
rect 16604 26516 16660 27806
rect 16716 26852 16772 30044
rect 16940 28756 16996 40348
rect 17052 38050 17108 38062
rect 17052 37998 17054 38050
rect 17106 37998 17108 38050
rect 17052 37156 17108 37998
rect 17052 37090 17108 37100
rect 17052 35700 17108 35710
rect 17052 29428 17108 35644
rect 17052 29362 17108 29372
rect 17052 28756 17108 28766
rect 16940 28754 17108 28756
rect 16940 28702 17054 28754
rect 17106 28702 17108 28754
rect 16940 28700 17108 28702
rect 17052 28532 17108 28700
rect 17052 28466 17108 28476
rect 16828 27970 16884 27982
rect 16828 27918 16830 27970
rect 16882 27918 16884 27970
rect 16828 27412 16884 27918
rect 16828 27346 16884 27356
rect 17164 27188 17220 47180
rect 17388 45556 17444 48190
rect 17836 46898 17892 49420
rect 17836 46846 17838 46898
rect 17890 46846 17892 46898
rect 17836 46834 17892 46846
rect 17948 48356 18004 48366
rect 18060 48356 18116 49982
rect 17948 48354 18116 48356
rect 17948 48302 17950 48354
rect 18002 48302 18116 48354
rect 17948 48300 18116 48302
rect 17388 45490 17444 45500
rect 17500 46228 17556 46238
rect 17500 45330 17556 46172
rect 17500 45278 17502 45330
rect 17554 45278 17556 45330
rect 17500 45266 17556 45278
rect 17612 45780 17668 45790
rect 17500 45106 17556 45118
rect 17500 45054 17502 45106
rect 17554 45054 17556 45106
rect 17500 44996 17556 45054
rect 17388 44436 17444 44446
rect 17388 42084 17444 44380
rect 17500 42644 17556 44940
rect 17612 43650 17668 45724
rect 17948 45220 18004 48300
rect 18172 46340 18228 51324
rect 18284 51154 18340 52780
rect 18396 52162 18452 53004
rect 18508 52994 18564 53004
rect 18844 53060 18900 53118
rect 18844 52994 18900 53004
rect 18956 52836 19012 56588
rect 19180 53956 19236 53966
rect 19180 52946 19236 53900
rect 19180 52894 19182 52946
rect 19234 52894 19236 52946
rect 19180 52882 19236 52894
rect 19292 53618 19348 53630
rect 19292 53566 19294 53618
rect 19346 53566 19348 53618
rect 18956 52770 19012 52780
rect 19292 52276 19348 53566
rect 19404 53060 19460 53070
rect 19404 52966 19460 53004
rect 18396 52110 18398 52162
rect 18450 52110 18452 52162
rect 18396 51380 18452 52110
rect 18732 52274 19348 52276
rect 18732 52222 19294 52274
rect 19346 52222 19348 52274
rect 18732 52220 19348 52222
rect 18396 51314 18452 51324
rect 18620 51492 18676 51502
rect 18284 51102 18286 51154
rect 18338 51102 18340 51154
rect 18284 51044 18340 51102
rect 18284 50978 18340 50988
rect 18620 51154 18676 51436
rect 18620 51102 18622 51154
rect 18674 51102 18676 51154
rect 18620 51044 18676 51102
rect 18620 50978 18676 50988
rect 18620 50820 18676 50830
rect 18620 50594 18676 50764
rect 18620 50542 18622 50594
rect 18674 50542 18676 50594
rect 18620 50530 18676 50542
rect 18508 50372 18564 50382
rect 18508 47458 18564 50316
rect 18620 49924 18676 49934
rect 18620 49830 18676 49868
rect 18620 49028 18676 49038
rect 18620 48934 18676 48972
rect 18508 47406 18510 47458
rect 18562 47406 18564 47458
rect 18508 47394 18564 47406
rect 18732 46788 18788 52220
rect 19292 52210 19348 52220
rect 18396 46564 18452 46574
rect 18172 46274 18228 46284
rect 18284 46452 18340 46462
rect 17612 43598 17614 43650
rect 17666 43598 17668 43650
rect 17612 43586 17668 43598
rect 17724 45218 18004 45220
rect 17724 45166 17950 45218
rect 18002 45166 18004 45218
rect 17724 45164 18004 45166
rect 17724 44212 17780 45164
rect 17948 45154 18004 45164
rect 18060 44324 18116 44334
rect 17724 43652 17780 44156
rect 17836 44322 18116 44324
rect 17836 44270 18062 44322
rect 18114 44270 18116 44322
rect 17836 44268 18116 44270
rect 17836 44100 17892 44268
rect 18060 44258 18116 44268
rect 17836 44034 17892 44044
rect 18172 44098 18228 44110
rect 18172 44046 18174 44098
rect 18226 44046 18228 44098
rect 17836 43652 17892 43662
rect 17724 43650 17892 43652
rect 17724 43598 17838 43650
rect 17890 43598 17892 43650
rect 17724 43596 17892 43598
rect 17612 42644 17668 42654
rect 17500 42642 17668 42644
rect 17500 42590 17614 42642
rect 17666 42590 17668 42642
rect 17500 42588 17668 42590
rect 17500 42084 17556 42094
rect 17388 42082 17556 42084
rect 17388 42030 17502 42082
rect 17554 42030 17556 42082
rect 17388 42028 17556 42030
rect 17388 40404 17444 42028
rect 17500 42018 17556 42028
rect 17500 41076 17556 41086
rect 17612 41076 17668 42588
rect 17500 41074 17668 41076
rect 17500 41022 17502 41074
rect 17554 41022 17668 41074
rect 17500 41020 17668 41022
rect 17500 41010 17556 41020
rect 17276 40402 17444 40404
rect 17276 40350 17390 40402
rect 17442 40350 17444 40402
rect 17276 40348 17444 40350
rect 17276 40292 17332 40348
rect 17388 40338 17444 40348
rect 17500 40626 17556 40638
rect 17500 40574 17502 40626
rect 17554 40574 17556 40626
rect 17500 40404 17556 40574
rect 17612 40516 17668 41020
rect 17836 41076 17892 43596
rect 18060 42754 18116 42766
rect 18060 42702 18062 42754
rect 18114 42702 18116 42754
rect 18060 41972 18116 42702
rect 18060 41906 18116 41916
rect 17836 40516 17892 41020
rect 18172 40740 18228 44046
rect 18060 40684 18228 40740
rect 17948 40516 18004 40526
rect 17612 40450 17668 40460
rect 17724 40514 18004 40516
rect 17724 40462 17950 40514
rect 18002 40462 18004 40514
rect 17724 40460 18004 40462
rect 17500 40338 17556 40348
rect 17276 40226 17332 40236
rect 17388 40180 17444 40190
rect 17388 38946 17444 40124
rect 17724 39506 17780 40460
rect 17948 40450 18004 40460
rect 17724 39454 17726 39506
rect 17778 39454 17780 39506
rect 17724 39442 17780 39454
rect 17388 38894 17390 38946
rect 17442 38894 17444 38946
rect 17388 38882 17444 38894
rect 17724 38946 17780 38958
rect 17724 38894 17726 38946
rect 17778 38894 17780 38946
rect 17612 38724 17668 38734
rect 17388 37828 17444 37838
rect 17388 37734 17444 37772
rect 17276 36820 17332 36830
rect 17276 36596 17332 36764
rect 17276 36502 17332 36540
rect 17500 35812 17556 35822
rect 17500 35718 17556 35756
rect 17388 35588 17444 35598
rect 17388 35494 17444 35532
rect 17612 35140 17668 38668
rect 17724 38668 17780 38894
rect 17724 38612 18004 38668
rect 17948 38610 18004 38612
rect 17948 38558 17950 38610
rect 18002 38558 18004 38610
rect 17948 38546 18004 38558
rect 17724 38052 17780 38062
rect 17724 38050 17892 38052
rect 17724 37998 17726 38050
rect 17778 37998 17892 38050
rect 17724 37996 17892 37998
rect 17724 37986 17780 37996
rect 17388 35084 17668 35140
rect 17724 37156 17780 37166
rect 17724 35140 17780 37100
rect 17836 36820 17892 37996
rect 17836 36754 17892 36764
rect 17836 36596 17892 36606
rect 17836 35810 17892 36540
rect 17836 35758 17838 35810
rect 17890 35758 17892 35810
rect 17836 35746 17892 35758
rect 17948 35700 18004 35710
rect 17948 35606 18004 35644
rect 18060 35476 18116 40684
rect 18172 40516 18228 40526
rect 18172 39618 18228 40460
rect 18172 39566 18174 39618
rect 18226 39566 18228 39618
rect 18172 39554 18228 39566
rect 18060 35410 18116 35420
rect 18172 39394 18228 39406
rect 18172 39342 18174 39394
rect 18226 39342 18228 39394
rect 17388 34580 17444 35084
rect 17724 35074 17780 35084
rect 18172 35028 18228 39342
rect 18284 38500 18340 46396
rect 18396 45890 18452 46508
rect 18396 45838 18398 45890
rect 18450 45838 18452 45890
rect 18396 45780 18452 45838
rect 18396 45714 18452 45724
rect 18508 44884 18564 44894
rect 18508 44210 18564 44828
rect 18732 44436 18788 46732
rect 18732 44370 18788 44380
rect 18844 51940 18900 51950
rect 19628 51940 19684 63758
rect 19836 62748 20100 62758
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 19836 62682 20100 62692
rect 20076 62468 20132 62478
rect 20076 62374 20132 62412
rect 20188 61572 20244 61582
rect 20188 61570 20356 61572
rect 20188 61518 20190 61570
rect 20242 61518 20356 61570
rect 20188 61516 20356 61518
rect 20188 61506 20244 61516
rect 20300 61458 20356 61516
rect 20300 61406 20302 61458
rect 20354 61406 20356 61458
rect 20300 61394 20356 61406
rect 20076 61348 20132 61386
rect 20076 61282 20132 61292
rect 19836 61180 20100 61190
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 19836 61114 20100 61124
rect 20300 60674 20356 60686
rect 20300 60622 20302 60674
rect 20354 60622 20356 60674
rect 20300 60562 20356 60622
rect 20300 60510 20302 60562
rect 20354 60510 20356 60562
rect 19836 59612 20100 59622
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 19836 59546 20100 59556
rect 20300 58548 20356 60510
rect 20300 58482 20356 58492
rect 20412 60002 20468 66220
rect 20636 66274 20692 67678
rect 21420 67956 21476 67966
rect 20860 67618 20916 67630
rect 20860 67566 20862 67618
rect 20914 67566 20916 67618
rect 20748 67172 20804 67182
rect 20860 67172 20916 67566
rect 20748 67170 20916 67172
rect 20748 67118 20750 67170
rect 20802 67118 20916 67170
rect 20748 67116 20916 67118
rect 20748 67106 20804 67116
rect 21420 66388 21476 67900
rect 21644 67732 21700 67742
rect 21532 67620 21588 67630
rect 21532 67526 21588 67564
rect 21420 66294 21476 66332
rect 20636 66222 20638 66274
rect 20690 66222 20692 66274
rect 20636 66210 20692 66222
rect 20524 66052 20580 66062
rect 20524 65602 20580 65996
rect 20524 65550 20526 65602
rect 20578 65550 20580 65602
rect 20524 65538 20580 65550
rect 21196 65492 21252 65502
rect 21196 65398 21252 65436
rect 21308 65380 21364 65390
rect 20748 64708 20804 64718
rect 20748 64614 20804 64652
rect 21308 64706 21364 65324
rect 21308 64654 21310 64706
rect 21362 64654 21364 64706
rect 21308 64642 21364 64654
rect 21644 64596 21700 67676
rect 21756 65604 21812 69804
rect 21980 69412 22036 74732
rect 22204 74004 22260 74844
rect 22428 74834 22484 74844
rect 22540 74340 22596 77980
rect 22540 73948 22596 74284
rect 22204 72658 22260 73948
rect 22204 72606 22206 72658
rect 22258 72606 22260 72658
rect 22204 72594 22260 72606
rect 22428 73892 22596 73948
rect 22652 75794 22708 78764
rect 23436 78708 23492 78718
rect 23436 78614 23492 78652
rect 22764 78596 22820 78606
rect 22764 78502 22820 78540
rect 22876 78594 22932 78606
rect 22876 78542 22878 78594
rect 22930 78542 22932 78594
rect 22652 75742 22654 75794
rect 22706 75742 22708 75794
rect 22652 73948 22708 75742
rect 22876 75124 22932 78542
rect 22988 78596 23044 78606
rect 22988 78594 23156 78596
rect 22988 78542 22990 78594
rect 23042 78542 23156 78594
rect 22988 78540 23156 78542
rect 22988 78530 23044 78540
rect 23100 76468 23156 78540
rect 23548 78034 23604 82574
rect 23660 82180 23716 86044
rect 23884 85988 23940 88284
rect 23660 82114 23716 82124
rect 23772 85932 23940 85988
rect 23996 88284 24164 88340
rect 24556 88898 24612 88910
rect 24556 88846 24558 88898
rect 24610 88846 24612 88898
rect 23772 81732 23828 85932
rect 23884 84532 23940 84542
rect 23884 84438 23940 84476
rect 23660 81676 23828 81732
rect 23660 80388 23716 81676
rect 23996 81620 24052 88284
rect 24108 88116 24164 88126
rect 24108 87668 24164 88060
rect 24556 87892 24612 88846
rect 24892 88338 24948 89180
rect 25116 89570 25172 89582
rect 25116 89518 25118 89570
rect 25170 89518 25172 89570
rect 25116 88788 25172 89518
rect 25228 89124 25284 89134
rect 25228 89010 25284 89068
rect 25228 88958 25230 89010
rect 25282 88958 25284 89010
rect 25228 88946 25284 88958
rect 25116 88722 25172 88732
rect 25004 88452 25060 88462
rect 25004 88450 25172 88452
rect 25004 88398 25006 88450
rect 25058 88398 25172 88450
rect 25004 88396 25172 88398
rect 25004 88386 25060 88396
rect 24892 88286 24894 88338
rect 24946 88286 24948 88338
rect 24556 87826 24612 87836
rect 24780 88226 24836 88238
rect 24780 88174 24782 88226
rect 24834 88174 24836 88226
rect 24780 88004 24836 88174
rect 24108 87612 24388 87668
rect 24332 87554 24388 87612
rect 24332 87502 24334 87554
rect 24386 87502 24388 87554
rect 24332 87490 24388 87502
rect 24556 87556 24612 87566
rect 24556 87462 24612 87500
rect 24220 87444 24276 87454
rect 24108 87442 24276 87444
rect 24108 87390 24222 87442
rect 24274 87390 24276 87442
rect 24108 87388 24276 87390
rect 24108 86772 24164 87388
rect 24220 87378 24276 87388
rect 24668 87444 24724 87454
rect 24668 87350 24724 87388
rect 24668 86884 24724 86894
rect 24668 86790 24724 86828
rect 24108 86716 24276 86772
rect 24108 86546 24164 86558
rect 24108 86494 24110 86546
rect 24162 86494 24164 86546
rect 24108 86436 24164 86494
rect 24108 86370 24164 86380
rect 24220 85708 24276 86716
rect 24332 86658 24388 86670
rect 24780 86660 24836 87948
rect 24332 86606 24334 86658
rect 24386 86606 24388 86658
rect 24332 86212 24388 86606
rect 24332 86146 24388 86156
rect 24556 86604 24836 86660
rect 24892 86660 24948 88286
rect 24108 85652 24276 85708
rect 24108 82404 24164 85652
rect 24220 84644 24276 84654
rect 24220 84418 24276 84588
rect 24220 84366 24222 84418
rect 24274 84366 24276 84418
rect 24220 84354 24276 84366
rect 24444 84308 24500 84318
rect 24444 84214 24500 84252
rect 24108 82338 24164 82348
rect 24220 84196 24276 84206
rect 23772 81564 24052 81620
rect 24108 82180 24164 82190
rect 23772 80500 23828 81564
rect 23772 80434 23828 80444
rect 23996 81284 24052 81294
rect 23996 80946 24052 81228
rect 23996 80894 23998 80946
rect 24050 80894 24052 80946
rect 23660 79828 23716 80332
rect 23660 79772 23828 79828
rect 23660 79602 23716 79614
rect 23660 79550 23662 79602
rect 23714 79550 23716 79602
rect 23660 79492 23716 79550
rect 23660 79426 23716 79436
rect 23548 77982 23550 78034
rect 23602 77982 23604 78034
rect 23548 77970 23604 77982
rect 23772 77924 23828 79772
rect 23884 79604 23940 79614
rect 23884 79510 23940 79548
rect 23996 79380 24052 80894
rect 24108 80500 24164 82124
rect 24108 80434 24164 80444
rect 23884 79324 24052 79380
rect 23884 78932 23940 79324
rect 23884 78866 23940 78876
rect 23996 78820 24052 78830
rect 23996 78726 24052 78764
rect 23100 76412 23716 76468
rect 22876 75058 22932 75068
rect 22876 74898 22932 74910
rect 22876 74846 22878 74898
rect 22930 74846 22932 74898
rect 22652 73892 22820 73948
rect 22428 71090 22484 73892
rect 22540 72772 22596 72782
rect 22540 71874 22596 72716
rect 22540 71822 22542 71874
rect 22594 71822 22596 71874
rect 22540 71810 22596 71822
rect 22428 71038 22430 71090
rect 22482 71038 22484 71090
rect 22316 70196 22372 70206
rect 22092 69412 22148 69422
rect 21980 69410 22148 69412
rect 21980 69358 22094 69410
rect 22146 69358 22148 69410
rect 21980 69356 22148 69358
rect 22092 69346 22148 69356
rect 22316 67732 22372 70140
rect 22428 67956 22484 71038
rect 22764 70308 22820 73892
rect 22876 71652 22932 74846
rect 22988 74900 23044 74910
rect 22988 74806 23044 74844
rect 23100 74900 23156 74910
rect 23324 74900 23380 74910
rect 23100 74898 23380 74900
rect 23100 74846 23102 74898
rect 23154 74846 23326 74898
rect 23378 74846 23380 74898
rect 23100 74844 23380 74846
rect 23100 74116 23156 74844
rect 23324 74834 23380 74844
rect 23100 73442 23156 74060
rect 23100 73390 23102 73442
rect 23154 73390 23156 73442
rect 23100 73378 23156 73390
rect 23548 74786 23604 74798
rect 23548 74734 23550 74786
rect 23602 74734 23604 74786
rect 23548 72772 23604 74734
rect 23660 74226 23716 76412
rect 23772 76132 23828 77868
rect 24108 78706 24164 78718
rect 24108 78654 24110 78706
rect 24162 78654 24164 78706
rect 24108 76580 24164 78654
rect 24108 76514 24164 76524
rect 24220 76468 24276 84140
rect 24556 82348 24612 86604
rect 24892 86594 24948 86604
rect 25004 87892 25060 87902
rect 24444 82292 24612 82348
rect 24668 86436 24724 86446
rect 24332 81170 24388 81182
rect 24332 81118 24334 81170
rect 24386 81118 24388 81170
rect 24332 79044 24388 81118
rect 24444 79716 24500 82292
rect 24556 81172 24612 81182
rect 24668 81172 24724 86380
rect 24892 86100 24948 86110
rect 24556 81170 24724 81172
rect 24556 81118 24558 81170
rect 24610 81118 24724 81170
rect 24556 81116 24724 81118
rect 24780 83522 24836 83534
rect 24780 83470 24782 83522
rect 24834 83470 24836 83522
rect 24556 81106 24612 81116
rect 24780 80724 24836 83470
rect 24892 82068 24948 86044
rect 25004 84308 25060 87836
rect 25116 86996 25172 88396
rect 25340 87780 25396 90636
rect 25676 90578 25732 92092
rect 25676 90526 25678 90578
rect 25730 90526 25732 90578
rect 25676 90514 25732 90526
rect 25116 86930 25172 86940
rect 25228 87724 25396 87780
rect 25452 90468 25508 90478
rect 25116 86772 25172 86782
rect 25116 86658 25172 86716
rect 25116 86606 25118 86658
rect 25170 86606 25172 86658
rect 25116 86594 25172 86606
rect 25228 86100 25284 87724
rect 25452 87668 25508 90412
rect 25788 89570 25844 89582
rect 25788 89518 25790 89570
rect 25842 89518 25844 89570
rect 25788 88900 25844 89518
rect 25900 89572 25956 92204
rect 26124 92194 26180 92204
rect 26124 92034 26180 92046
rect 26124 91982 26126 92034
rect 26178 91982 26180 92034
rect 26124 91924 26180 91982
rect 26124 91858 26180 91868
rect 26012 90692 26068 90702
rect 26236 90692 26292 92764
rect 26012 90690 26292 90692
rect 26012 90638 26014 90690
rect 26066 90638 26292 90690
rect 26012 90636 26292 90638
rect 26012 90626 26068 90636
rect 26236 90354 26292 90366
rect 26236 90302 26238 90354
rect 26290 90302 26292 90354
rect 26012 89572 26068 89582
rect 25900 89570 26068 89572
rect 25900 89518 26014 89570
rect 26066 89518 26068 89570
rect 25900 89516 26068 89518
rect 25564 88004 25620 88014
rect 25564 87910 25620 87948
rect 25452 87602 25508 87612
rect 25116 86044 25284 86100
rect 25340 87556 25396 87566
rect 25116 85708 25172 86044
rect 25340 85986 25396 87500
rect 25340 85934 25342 85986
rect 25394 85934 25396 85986
rect 25340 85922 25396 85934
rect 25676 87442 25732 87454
rect 25676 87390 25678 87442
rect 25730 87390 25732 87442
rect 25228 85876 25284 85886
rect 25228 85782 25284 85820
rect 25676 85708 25732 87390
rect 25116 85652 25396 85708
rect 25228 84308 25284 84318
rect 25004 84306 25284 84308
rect 25004 84254 25230 84306
rect 25282 84254 25284 84306
rect 25004 84252 25284 84254
rect 25228 84242 25284 84252
rect 25228 82740 25284 82750
rect 25228 82646 25284 82684
rect 24892 82002 24948 82012
rect 25004 81956 25060 81966
rect 24780 80658 24836 80668
rect 24892 81732 24948 81742
rect 24444 79660 24612 79716
rect 24444 79490 24500 79502
rect 24444 79438 24446 79490
rect 24498 79438 24500 79490
rect 24444 79378 24500 79438
rect 24444 79326 24446 79378
rect 24498 79326 24500 79378
rect 24444 79314 24500 79326
rect 24556 78988 24612 79660
rect 24892 79492 24948 81676
rect 25004 81284 25060 81900
rect 25004 81218 25060 81228
rect 25228 81170 25284 81182
rect 25228 81118 25230 81170
rect 25282 81118 25284 81170
rect 24780 79436 24948 79492
rect 25004 79492 25060 79502
rect 24780 79378 24836 79436
rect 24780 79326 24782 79378
rect 24834 79326 24836 79378
rect 24780 79314 24836 79326
rect 24332 78978 24388 78988
rect 24444 78932 24612 78988
rect 24332 78596 24388 78606
rect 24332 78502 24388 78540
rect 24220 76402 24276 76412
rect 24332 76692 24388 76702
rect 24444 76692 24500 78932
rect 25004 78930 25060 79436
rect 25004 78878 25006 78930
rect 25058 78878 25060 78930
rect 25004 78866 25060 78878
rect 24332 76690 24500 76692
rect 24332 76638 24334 76690
rect 24386 76638 24500 76690
rect 24332 76636 24500 76638
rect 24556 78818 24612 78830
rect 24556 78766 24558 78818
rect 24610 78766 24612 78818
rect 24556 76692 24612 78766
rect 24780 78706 24836 78718
rect 24780 78654 24782 78706
rect 24834 78654 24836 78706
rect 24780 78596 24836 78654
rect 24780 78530 24836 78540
rect 25228 78036 25284 81118
rect 25340 78930 25396 85652
rect 25564 85652 25732 85708
rect 25788 85708 25844 88844
rect 25900 88788 25956 88798
rect 25900 86658 25956 88732
rect 26012 86882 26068 89516
rect 26124 89572 26180 89582
rect 26124 89478 26180 89516
rect 26236 89570 26292 90302
rect 26236 89518 26238 89570
rect 26290 89518 26292 89570
rect 26236 89460 26292 89518
rect 26236 89394 26292 89404
rect 26012 86830 26014 86882
rect 26066 86830 26068 86882
rect 26012 86818 26068 86830
rect 26236 87668 26292 87678
rect 25900 86606 25902 86658
rect 25954 86606 25956 86658
rect 25900 86436 25956 86606
rect 26124 86770 26180 86782
rect 26124 86718 26126 86770
rect 26178 86718 26180 86770
rect 26124 86660 26180 86718
rect 26124 86594 26180 86604
rect 25900 86380 26180 86436
rect 25788 85652 25956 85708
rect 25564 84978 25620 85652
rect 25564 84926 25566 84978
rect 25618 84926 25620 84978
rect 25452 84194 25508 84206
rect 25452 84142 25454 84194
rect 25506 84142 25508 84194
rect 25452 82516 25508 84142
rect 25452 82450 25508 82460
rect 25564 81954 25620 84926
rect 25676 84532 25732 84542
rect 25676 84438 25732 84476
rect 25900 84530 25956 85596
rect 25900 84478 25902 84530
rect 25954 84478 25956 84530
rect 25900 84466 25956 84478
rect 25788 84196 25844 84206
rect 25788 84102 25844 84140
rect 26012 83410 26068 83422
rect 26012 83358 26014 83410
rect 26066 83358 26068 83410
rect 25900 83188 25956 83198
rect 25900 82964 25956 83132
rect 25900 82738 25956 82908
rect 25900 82686 25902 82738
rect 25954 82686 25956 82738
rect 25900 82674 25956 82686
rect 25564 81902 25566 81954
rect 25618 81902 25620 81954
rect 25564 81890 25620 81902
rect 25788 82404 25844 82414
rect 25452 81844 25508 81854
rect 25452 81284 25508 81788
rect 25788 81732 25844 82348
rect 25452 81190 25508 81228
rect 25564 81676 25844 81732
rect 25900 82292 25956 82302
rect 25452 81060 25508 81070
rect 25564 81060 25620 81676
rect 25452 81058 25620 81060
rect 25452 81006 25454 81058
rect 25506 81006 25620 81058
rect 25452 81004 25620 81006
rect 25676 81170 25732 81182
rect 25676 81118 25678 81170
rect 25730 81118 25732 81170
rect 25452 80994 25508 81004
rect 25676 80948 25732 81118
rect 25676 80882 25732 80892
rect 25900 81170 25956 82236
rect 25900 81118 25902 81170
rect 25954 81118 25956 81170
rect 25340 78878 25342 78930
rect 25394 78878 25396 78930
rect 25340 78866 25396 78878
rect 25452 80724 25508 80734
rect 25452 80274 25508 80668
rect 25900 80724 25956 81118
rect 25900 80658 25956 80668
rect 26012 80612 26068 83358
rect 26124 81396 26180 86380
rect 26236 84756 26292 87612
rect 26236 84532 26292 84700
rect 26236 84466 26292 84476
rect 26236 83300 26292 83310
rect 26236 82626 26292 83244
rect 26236 82574 26238 82626
rect 26290 82574 26292 82626
rect 26236 82562 26292 82574
rect 26348 81956 26404 97412
rect 26796 97412 26852 97422
rect 26460 95954 26516 95966
rect 26460 95902 26462 95954
rect 26514 95902 26516 95954
rect 26460 95844 26516 95902
rect 26796 95954 26852 97356
rect 28476 97412 28532 99600
rect 28476 97346 28532 97356
rect 30156 96628 30212 96638
rect 30156 96626 30324 96628
rect 30156 96574 30158 96626
rect 30210 96574 30324 96626
rect 30156 96572 30324 96574
rect 30156 96562 30212 96572
rect 26796 95902 26798 95954
rect 26850 95902 26852 95954
rect 26796 95890 26852 95902
rect 29260 96066 29316 96078
rect 29260 96014 29262 96066
rect 29314 96014 29316 96066
rect 26460 95778 26516 95788
rect 27356 95844 27412 95854
rect 27412 95788 27524 95844
rect 27356 95750 27412 95788
rect 27356 95058 27412 95070
rect 27356 95006 27358 95058
rect 27410 95006 27412 95058
rect 27356 94612 27412 95006
rect 27356 93940 27412 94556
rect 27468 94276 27524 95788
rect 27804 95284 27860 95294
rect 27804 94498 27860 95228
rect 27804 94446 27806 94498
rect 27858 94446 27860 94498
rect 27468 94220 27636 94276
rect 27468 93940 27524 93950
rect 27356 93884 27468 93940
rect 27356 93490 27412 93884
rect 27468 93874 27524 93884
rect 27356 93438 27358 93490
rect 27410 93438 27412 93490
rect 27356 93426 27412 93438
rect 26684 92820 26740 92830
rect 26684 92726 26740 92764
rect 27468 92820 27524 92830
rect 27468 92726 27524 92764
rect 26460 92484 26516 92494
rect 26460 82852 26516 92428
rect 27356 92148 27412 92158
rect 27356 92054 27412 92092
rect 26572 90466 26628 90478
rect 26572 90414 26574 90466
rect 26626 90414 26628 90466
rect 26572 90354 26628 90414
rect 26572 90302 26574 90354
rect 26626 90302 26628 90354
rect 26572 90290 26628 90302
rect 27020 90468 27076 90478
rect 27468 90468 27524 90478
rect 27020 90466 27524 90468
rect 27020 90414 27022 90466
rect 27074 90414 27470 90466
rect 27522 90414 27524 90466
rect 27020 90412 27524 90414
rect 27020 89794 27076 90412
rect 27468 90402 27524 90412
rect 27020 89742 27022 89794
rect 27074 89742 27076 89794
rect 26572 89682 26628 89694
rect 26572 89630 26574 89682
rect 26626 89630 26628 89682
rect 26572 87444 26628 89630
rect 26572 87378 26628 87388
rect 26908 89124 26964 89134
rect 26908 86548 26964 89068
rect 27020 88004 27076 89742
rect 27020 87938 27076 87948
rect 27356 89906 27412 89918
rect 27356 89854 27358 89906
rect 27410 89854 27412 89906
rect 27356 88676 27412 89854
rect 27356 87892 27412 88620
rect 27356 87826 27412 87836
rect 27468 89012 27524 89022
rect 27244 87556 27300 87566
rect 27244 87462 27300 87500
rect 27132 87220 27188 87230
rect 27132 86658 27188 87164
rect 27132 86606 27134 86658
rect 27186 86606 27188 86658
rect 27132 86594 27188 86606
rect 26908 86454 26964 86492
rect 27020 86434 27076 86446
rect 27020 86382 27022 86434
rect 27074 86382 27076 86434
rect 26908 84308 26964 84318
rect 26908 84214 26964 84252
rect 27020 82852 27076 86382
rect 27356 86434 27412 86446
rect 27356 86382 27358 86434
rect 27410 86382 27412 86434
rect 27356 85652 27412 86382
rect 27468 85986 27524 88956
rect 27468 85934 27470 85986
rect 27522 85934 27524 85986
rect 27468 85922 27524 85934
rect 27356 85586 27412 85596
rect 27468 84980 27524 84990
rect 27356 84532 27412 84542
rect 27244 84476 27356 84532
rect 27132 84194 27188 84206
rect 27132 84142 27134 84194
rect 27186 84142 27188 84194
rect 27132 82964 27188 84142
rect 27132 82898 27188 82908
rect 26460 82758 26516 82796
rect 26796 82796 27076 82852
rect 26348 81890 26404 81900
rect 26572 82740 26628 82750
rect 26124 81340 26404 81396
rect 26348 80836 26404 81340
rect 26572 81394 26628 82684
rect 26684 82180 26740 82190
rect 26684 81508 26740 82124
rect 26796 81620 26852 82796
rect 27244 82738 27300 84476
rect 27356 84466 27412 84476
rect 27244 82686 27246 82738
rect 27298 82686 27300 82738
rect 27020 82628 27076 82638
rect 26908 82516 26964 82526
rect 26908 82068 26964 82460
rect 27020 82514 27076 82572
rect 27020 82462 27022 82514
rect 27074 82462 27076 82514
rect 27020 82450 27076 82462
rect 27132 82626 27188 82638
rect 27132 82574 27134 82626
rect 27186 82574 27188 82626
rect 27132 82516 27188 82574
rect 27020 82068 27076 82078
rect 26908 82066 27076 82068
rect 26908 82014 27022 82066
rect 27074 82014 27076 82066
rect 26908 82012 27076 82014
rect 27132 82068 27188 82460
rect 27244 82404 27300 82686
rect 27356 84308 27412 84318
rect 27356 82628 27412 84252
rect 27468 84196 27524 84924
rect 27468 84102 27524 84140
rect 27356 82562 27412 82572
rect 27244 82338 27300 82348
rect 27356 82180 27412 82190
rect 27356 82086 27412 82124
rect 27132 82012 27300 82068
rect 27020 82002 27076 82012
rect 26908 81844 26964 81854
rect 26908 81750 26964 81788
rect 27132 81842 27188 81854
rect 27132 81790 27134 81842
rect 27186 81790 27188 81842
rect 27132 81732 27188 81790
rect 27132 81666 27188 81676
rect 26796 81564 26964 81620
rect 26684 81452 26852 81508
rect 26572 81342 26574 81394
rect 26626 81342 26628 81394
rect 26572 81330 26628 81342
rect 26460 81172 26516 81182
rect 26460 81170 26628 81172
rect 26460 81118 26462 81170
rect 26514 81118 26628 81170
rect 26460 81116 26628 81118
rect 26460 81106 26516 81116
rect 26572 80836 26628 81116
rect 26348 80780 26516 80836
rect 26012 80546 26068 80556
rect 26348 80612 26404 80622
rect 25452 80222 25454 80274
rect 25506 80222 25508 80274
rect 25228 77980 25396 78036
rect 23772 76076 23940 76132
rect 23884 75908 23940 76076
rect 23884 75852 24052 75908
rect 23772 75012 23828 75022
rect 23772 74918 23828 74956
rect 23884 74900 23940 74910
rect 23884 74806 23940 74844
rect 23660 74174 23662 74226
rect 23714 74174 23716 74226
rect 23660 74162 23716 74174
rect 23548 72706 23604 72716
rect 23996 72212 24052 75852
rect 23996 72146 24052 72156
rect 24332 75012 24388 76636
rect 24556 76626 24612 76636
rect 24780 77922 24836 77934
rect 24780 77870 24782 77922
rect 24834 77870 24836 77922
rect 24668 76468 24724 76478
rect 24780 76468 24836 77870
rect 25228 77812 25284 77822
rect 24724 76412 24836 76468
rect 24892 77810 25284 77812
rect 24892 77758 25230 77810
rect 25282 77758 25284 77810
rect 24892 77756 25284 77758
rect 24556 75908 24612 75918
rect 24332 73444 24388 74956
rect 24444 75684 24500 75694
rect 24444 75010 24500 75628
rect 24556 75122 24612 75852
rect 24556 75070 24558 75122
rect 24610 75070 24612 75122
rect 24556 75058 24612 75070
rect 24444 74958 24446 75010
rect 24498 74958 24500 75010
rect 24444 74946 24500 74958
rect 22876 71586 22932 71596
rect 23884 70978 23940 70990
rect 23884 70926 23886 70978
rect 23938 70926 23940 70978
rect 23884 70756 23940 70926
rect 24332 70980 24388 73388
rect 24668 73220 24724 76412
rect 24780 75684 24836 75694
rect 24892 75684 24948 77756
rect 25228 77746 25284 77756
rect 25228 77588 25284 77598
rect 25228 76466 25284 77532
rect 25340 77028 25396 77980
rect 25452 77250 25508 80222
rect 25788 80500 25844 80510
rect 25564 79044 25620 79054
rect 25564 78036 25620 78988
rect 25788 78930 25844 80444
rect 25788 78878 25790 78930
rect 25842 78878 25844 78930
rect 25788 78866 25844 78878
rect 25900 79602 25956 79614
rect 25900 79550 25902 79602
rect 25954 79550 25956 79602
rect 25676 78706 25732 78718
rect 25676 78654 25678 78706
rect 25730 78654 25732 78706
rect 25676 78596 25732 78654
rect 25788 78596 25844 78606
rect 25676 78540 25788 78596
rect 25788 78530 25844 78540
rect 25788 78148 25844 78158
rect 25564 77980 25732 78036
rect 25564 77810 25620 77822
rect 25564 77758 25566 77810
rect 25618 77758 25620 77810
rect 25564 77700 25620 77758
rect 25564 77634 25620 77644
rect 25452 77198 25454 77250
rect 25506 77198 25508 77250
rect 25452 77186 25508 77198
rect 25340 76972 25508 77028
rect 25340 76692 25396 76702
rect 25340 76598 25396 76636
rect 25228 76414 25230 76466
rect 25282 76414 25284 76466
rect 25228 76132 25284 76414
rect 25228 76076 25396 76132
rect 24780 75682 24948 75684
rect 24780 75630 24782 75682
rect 24834 75630 24948 75682
rect 24780 75628 24948 75630
rect 24780 75618 24836 75628
rect 25228 75124 25284 75134
rect 25228 75030 25284 75068
rect 25340 75012 25396 76076
rect 25340 74946 25396 74956
rect 24668 73154 24724 73164
rect 24780 74898 24836 74910
rect 24780 74846 24782 74898
rect 24834 74846 24836 74898
rect 24780 72772 24836 74846
rect 24780 72706 24836 72716
rect 25228 74900 25284 74910
rect 25228 72660 25284 74844
rect 25004 72434 25060 72446
rect 25004 72382 25006 72434
rect 25058 72382 25060 72434
rect 25004 72212 25060 72382
rect 24668 71652 24724 71662
rect 24668 71558 24724 71596
rect 25004 71090 25060 72156
rect 25004 71038 25006 71090
rect 25058 71038 25060 71090
rect 25004 71026 25060 71038
rect 24332 70914 24388 70924
rect 25228 70978 25284 72604
rect 25228 70926 25230 70978
rect 25282 70926 25284 70978
rect 25228 70914 25284 70926
rect 24332 70756 24388 70766
rect 23884 70754 24388 70756
rect 23884 70702 24334 70754
rect 24386 70702 24388 70754
rect 23884 70700 24388 70702
rect 22764 70252 23268 70308
rect 22428 67890 22484 67900
rect 23100 67732 23156 67742
rect 22316 67730 23156 67732
rect 22316 67678 23102 67730
rect 23154 67678 23156 67730
rect 22316 67676 23156 67678
rect 22316 67172 22372 67676
rect 23100 67666 23156 67676
rect 22316 67106 22372 67116
rect 22876 66946 22932 66958
rect 22876 66894 22878 66946
rect 22930 66894 22932 66946
rect 22092 66724 22148 66734
rect 22092 66274 22148 66668
rect 22092 66222 22094 66274
rect 22146 66222 22148 66274
rect 22092 66210 22148 66222
rect 22316 66388 22372 66398
rect 21756 65548 22148 65604
rect 21868 65378 21924 65390
rect 21868 65326 21870 65378
rect 21922 65326 21924 65378
rect 21532 64484 21588 64494
rect 21532 64390 21588 64428
rect 21644 64260 21700 64540
rect 21308 64204 21700 64260
rect 21756 65266 21812 65278
rect 21756 65214 21758 65266
rect 21810 65214 21812 65266
rect 20860 64036 20916 64046
rect 20748 63252 20804 63262
rect 20524 63250 20804 63252
rect 20524 63198 20750 63250
rect 20802 63198 20804 63250
rect 20524 63196 20804 63198
rect 20524 61458 20580 63196
rect 20748 63186 20804 63196
rect 20860 62188 20916 63980
rect 21196 63924 21252 63934
rect 21196 63830 21252 63868
rect 21196 62466 21252 62478
rect 21196 62414 21198 62466
rect 21250 62414 21252 62466
rect 20748 62132 20916 62188
rect 21084 62356 21140 62366
rect 20748 61684 20804 62132
rect 20524 61406 20526 61458
rect 20578 61406 20580 61458
rect 20524 61394 20580 61406
rect 20636 61682 20804 61684
rect 20636 61630 20750 61682
rect 20802 61630 20804 61682
rect 20636 61628 20804 61630
rect 20412 59950 20414 60002
rect 20466 59950 20468 60002
rect 19836 58044 20100 58054
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 19836 57978 20100 57988
rect 20188 57764 20244 57774
rect 19964 57652 20020 57662
rect 19964 57558 20020 57596
rect 19836 56476 20100 56486
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 19836 56410 20100 56420
rect 19740 56308 19796 56318
rect 19740 55412 19796 56252
rect 19740 55318 19796 55356
rect 19836 54908 20100 54918
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 19836 54842 20100 54852
rect 19836 53340 20100 53350
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 19836 53274 20100 53284
rect 20188 53284 20244 57708
rect 20412 57538 20468 59950
rect 20524 60562 20580 60574
rect 20524 60510 20526 60562
rect 20578 60510 20580 60562
rect 20524 59780 20580 60510
rect 20636 60340 20692 61628
rect 20748 61618 20804 61628
rect 20748 60676 20804 60686
rect 20748 60582 20804 60620
rect 21084 60452 21140 62300
rect 21196 62244 21252 62414
rect 21196 62178 21252 62188
rect 21308 61124 21364 64204
rect 21420 63140 21476 63150
rect 21420 63046 21476 63084
rect 21420 62916 21476 62926
rect 21420 62822 21476 62860
rect 21756 62188 21812 65214
rect 21868 65268 21924 65326
rect 21980 65268 22036 65278
rect 21868 65212 21980 65268
rect 21980 65202 22036 65212
rect 22092 64820 22148 65548
rect 22316 65490 22372 66332
rect 22764 66164 22820 66174
rect 22652 66162 22820 66164
rect 22652 66110 22766 66162
rect 22818 66110 22820 66162
rect 22652 66108 22820 66110
rect 22652 65714 22708 66108
rect 22764 66098 22820 66108
rect 22652 65662 22654 65714
rect 22706 65662 22708 65714
rect 22652 65650 22708 65662
rect 22316 65438 22318 65490
rect 22370 65438 22372 65490
rect 22316 65380 22372 65438
rect 22316 65314 22372 65324
rect 22876 65268 22932 66894
rect 23212 66948 23268 70252
rect 24332 69300 24388 70700
rect 25452 70754 25508 76972
rect 25564 76468 25620 76478
rect 25564 76374 25620 76412
rect 25676 75124 25732 77980
rect 25788 78034 25844 78092
rect 25788 77982 25790 78034
rect 25842 77982 25844 78034
rect 25788 77970 25844 77982
rect 25900 77476 25956 79550
rect 26124 79604 26180 79614
rect 26124 78818 26180 79548
rect 26124 78766 26126 78818
rect 26178 78766 26180 78818
rect 26012 78708 26068 78718
rect 26012 78614 26068 78652
rect 26124 78148 26180 78766
rect 26348 78260 26404 80556
rect 26124 78054 26180 78092
rect 26236 78204 26404 78260
rect 25900 77420 26180 77476
rect 25788 76466 25844 76478
rect 25788 76414 25790 76466
rect 25842 76414 25844 76466
rect 25788 76356 25844 76414
rect 26012 76356 26068 76366
rect 25788 76300 26012 76356
rect 25676 75058 25732 75068
rect 25788 75348 25844 75358
rect 25788 74898 25844 75292
rect 25788 74846 25790 74898
rect 25842 74846 25844 74898
rect 25788 74834 25844 74846
rect 25564 74674 25620 74686
rect 25564 74622 25566 74674
rect 25618 74622 25620 74674
rect 25564 73948 25620 74622
rect 25564 73892 25956 73948
rect 25564 72772 25620 72782
rect 25900 72772 25956 73892
rect 26012 73556 26068 76300
rect 26124 75794 26180 77420
rect 26124 75742 26126 75794
rect 26178 75742 26180 75794
rect 26124 74114 26180 75742
rect 26236 76690 26292 78204
rect 26348 78036 26404 78046
rect 26348 77942 26404 77980
rect 26460 77812 26516 80780
rect 26572 80770 26628 80780
rect 26684 81060 26740 81070
rect 26684 78596 26740 81004
rect 26796 80948 26852 81452
rect 26908 81396 26964 81564
rect 26908 81340 27076 81396
rect 26908 80948 26964 80958
rect 26796 80946 26964 80948
rect 26796 80894 26910 80946
rect 26962 80894 26964 80946
rect 26796 80892 26964 80894
rect 26908 79604 26964 80892
rect 26908 79538 26964 79548
rect 27020 78820 27076 81340
rect 27132 81172 27188 81182
rect 27132 81078 27188 81116
rect 27244 80276 27300 82012
rect 27468 81956 27524 81966
rect 27356 81954 27524 81956
rect 27356 81902 27470 81954
rect 27522 81902 27524 81954
rect 27356 81900 27524 81902
rect 27356 80948 27412 81900
rect 27468 81890 27524 81900
rect 27468 81508 27524 81518
rect 27468 81170 27524 81452
rect 27468 81118 27470 81170
rect 27522 81118 27524 81170
rect 27468 81106 27524 81118
rect 27356 80892 27524 80948
rect 27132 80220 27300 80276
rect 27132 79156 27188 80220
rect 27244 79492 27300 79502
rect 27244 79398 27300 79436
rect 27132 79090 27188 79100
rect 27468 79044 27524 80892
rect 27580 80724 27636 94220
rect 27804 92034 27860 94446
rect 28252 95282 28308 95294
rect 28252 95230 28254 95282
rect 28306 95230 28308 95282
rect 28252 94500 28308 95230
rect 29148 95284 29204 95294
rect 29148 95190 29204 95228
rect 28588 94500 28644 94510
rect 28252 94498 28644 94500
rect 28252 94446 28590 94498
rect 28642 94446 28644 94498
rect 28252 94444 28644 94446
rect 28588 93716 28644 94444
rect 29260 94498 29316 96014
rect 30156 96068 30212 96078
rect 29260 94446 29262 94498
rect 29314 94446 29316 94498
rect 28812 93716 28868 93726
rect 29260 93716 29316 94446
rect 28588 93714 29316 93716
rect 28588 93662 28814 93714
rect 28866 93662 29316 93714
rect 28588 93660 29316 93662
rect 28812 93650 28868 93660
rect 29260 92930 29316 93660
rect 29596 95284 29652 95294
rect 29596 93714 29652 95228
rect 29596 93662 29598 93714
rect 29650 93662 29652 93714
rect 29596 93650 29652 93662
rect 30156 95284 30212 96012
rect 30156 94498 30212 95228
rect 30268 95172 30324 96572
rect 30940 95732 30996 99600
rect 31276 96850 31332 96862
rect 31276 96798 31278 96850
rect 31330 96798 31332 96850
rect 31276 96068 31332 96798
rect 32284 96852 32340 96862
rect 32284 96758 32340 96796
rect 32956 96852 33012 96862
rect 31276 96002 31332 96012
rect 32956 96066 33012 96796
rect 32956 96014 32958 96066
rect 33010 96014 33012 96066
rect 30940 95666 30996 95676
rect 31500 95842 31556 95854
rect 31500 95790 31502 95842
rect 31554 95790 31556 95842
rect 30492 95172 30548 95182
rect 30268 95170 30548 95172
rect 30268 95118 30494 95170
rect 30546 95118 30548 95170
rect 30268 95116 30548 95118
rect 30156 94446 30158 94498
rect 30210 94446 30212 94498
rect 29260 92878 29262 92930
rect 29314 92878 29316 92930
rect 29260 92820 29316 92878
rect 30156 92932 30212 94446
rect 30492 93940 30548 95116
rect 30492 93492 30548 93884
rect 31500 94274 31556 95790
rect 32956 95284 33012 96014
rect 33180 96626 33236 96638
rect 33180 96574 33182 96626
rect 33234 96574 33236 96626
rect 33180 95844 33236 96574
rect 33404 95956 33460 99600
rect 35196 98028 35460 98038
rect 35252 97972 35300 98028
rect 35356 97972 35404 98028
rect 35196 97962 35460 97972
rect 34300 96850 34356 96862
rect 34300 96798 34302 96850
rect 34354 96798 34356 96850
rect 33404 95890 33460 95900
rect 33852 96068 33908 96078
rect 34300 96068 34356 96798
rect 35196 96852 35252 96862
rect 35196 96758 35252 96796
rect 35196 96460 35460 96470
rect 35252 96404 35300 96460
rect 35356 96404 35404 96460
rect 35196 96394 35460 96404
rect 35868 96180 35924 99600
rect 35868 96114 35924 96124
rect 33852 96066 34356 96068
rect 33852 96014 33854 96066
rect 33906 96014 34356 96066
rect 33852 96012 34356 96014
rect 33180 95778 33236 95788
rect 33068 95284 33124 95294
rect 32956 95228 33068 95284
rect 31500 94222 31502 94274
rect 31554 94222 31556 94274
rect 30828 93492 30884 93502
rect 30492 93490 30996 93492
rect 30492 93438 30830 93490
rect 30882 93438 30996 93490
rect 30492 93436 30996 93438
rect 30828 93426 30884 93436
rect 30940 93156 30996 93436
rect 30940 93090 30996 93100
rect 31500 93156 31556 94222
rect 32844 94500 32900 94510
rect 33068 94500 33124 95228
rect 32844 94498 33124 94500
rect 32844 94446 32846 94498
rect 32898 94446 33124 94498
rect 32844 94444 33124 94446
rect 33852 95172 33908 96012
rect 35196 95844 35252 95854
rect 34076 95282 34132 95294
rect 34076 95230 34078 95282
rect 34130 95230 34132 95282
rect 34076 95172 34132 95230
rect 33852 95116 34076 95172
rect 33852 94498 33908 95116
rect 34076 95106 34132 95116
rect 35196 95060 35252 95788
rect 35644 95284 35700 95294
rect 35644 95190 35700 95228
rect 36428 95282 36484 95294
rect 36428 95230 36430 95282
rect 36482 95230 36484 95282
rect 36428 95172 36484 95230
rect 36428 95106 36484 95116
rect 34972 95004 35196 95060
rect 34972 94722 35028 95004
rect 34972 94670 34974 94722
rect 35026 94670 35028 94722
rect 34972 94658 35028 94670
rect 33852 94446 33854 94498
rect 33906 94446 33908 94498
rect 31500 93042 31556 93100
rect 31500 92990 31502 93042
rect 31554 92990 31556 93042
rect 31500 92978 31556 92990
rect 31836 94052 31892 94062
rect 30156 92838 30212 92876
rect 31836 92930 31892 93996
rect 32844 94052 32900 94444
rect 32844 93986 32900 93996
rect 33180 93714 33236 93726
rect 33180 93662 33182 93714
rect 33234 93662 33236 93714
rect 31836 92878 31838 92930
rect 31890 92878 31892 92930
rect 29260 92754 29316 92764
rect 31836 92820 31892 92878
rect 31836 92754 31892 92764
rect 32508 93044 32564 93054
rect 32508 92708 32564 92988
rect 32732 92932 32788 92942
rect 32732 92838 32788 92876
rect 27804 91982 27806 92034
rect 27858 91982 27860 92034
rect 27804 91970 27860 91982
rect 28364 92036 28420 92046
rect 27692 91362 27748 91374
rect 27692 91310 27694 91362
rect 27746 91310 27748 91362
rect 27692 88900 27748 91310
rect 28364 90748 28420 91980
rect 32508 91586 32564 92652
rect 32508 91534 32510 91586
rect 32562 91534 32564 91586
rect 32508 91522 32564 91534
rect 33180 92820 33236 93662
rect 33180 92146 33236 92764
rect 33180 92094 33182 92146
rect 33234 92094 33236 92146
rect 33180 91364 33236 92094
rect 33180 91298 33236 91308
rect 33852 93714 33908 94446
rect 33852 93662 33854 93714
rect 33906 93662 33908 93714
rect 33852 92932 33908 93662
rect 33852 92146 33908 92876
rect 35084 93492 35140 95004
rect 35196 94994 35252 95004
rect 37772 95060 37828 95070
rect 37772 94966 37828 95004
rect 35196 94892 35460 94902
rect 35252 94836 35300 94892
rect 35356 94836 35404 94892
rect 35196 94826 35460 94836
rect 35196 93492 35252 93502
rect 35084 93490 35252 93492
rect 35084 93438 35198 93490
rect 35250 93438 35252 93490
rect 35084 93436 35252 93438
rect 34076 92708 34132 92718
rect 34076 92614 34132 92652
rect 35084 92708 35140 93436
rect 35196 93426 35252 93436
rect 35196 93324 35460 93334
rect 35252 93268 35300 93324
rect 35356 93268 35404 93324
rect 35196 93258 35460 93268
rect 33852 92094 33854 92146
rect 33906 92094 33908 92146
rect 33852 91362 33908 92094
rect 35084 91924 35140 92652
rect 37884 92258 37940 92270
rect 37884 92206 37886 92258
rect 37938 92206 37940 92258
rect 37660 92036 37716 92046
rect 37660 91942 37716 91980
rect 35196 91924 35252 91934
rect 35084 91922 35252 91924
rect 35084 91870 35198 91922
rect 35250 91870 35252 91922
rect 35084 91868 35252 91870
rect 35196 91858 35252 91868
rect 35196 91756 35460 91766
rect 35252 91700 35300 91756
rect 35356 91700 35404 91756
rect 35196 91690 35460 91700
rect 33852 91310 33854 91362
rect 33906 91310 33908 91362
rect 33852 91298 33908 91310
rect 34524 91364 34580 91374
rect 34524 91270 34580 91308
rect 28364 90692 28532 90748
rect 27916 90468 27972 90478
rect 28252 90468 28308 90478
rect 27916 90466 28084 90468
rect 27916 90414 27918 90466
rect 27970 90414 28084 90466
rect 27916 90412 28084 90414
rect 27916 90402 27972 90412
rect 28028 89570 28084 90412
rect 28252 90374 28308 90412
rect 28028 89518 28030 89570
rect 28082 89518 28084 89570
rect 28028 89124 28084 89518
rect 28028 89058 28084 89068
rect 28476 89570 28532 90692
rect 29708 90692 29764 90702
rect 29708 90598 29764 90636
rect 30156 90692 30212 90702
rect 30156 90598 30212 90636
rect 35084 90692 35140 90702
rect 30268 90578 30324 90590
rect 30268 90526 30270 90578
rect 30322 90526 30324 90578
rect 30156 90356 30212 90366
rect 30044 90354 30212 90356
rect 30044 90302 30158 90354
rect 30210 90302 30212 90354
rect 30044 90300 30212 90302
rect 28476 89518 28478 89570
rect 28530 89518 28532 89570
rect 27692 88834 27748 88844
rect 27804 88116 27860 88126
rect 27804 88022 27860 88060
rect 28028 86996 28084 87006
rect 28476 86996 28532 89518
rect 29260 89570 29316 89582
rect 29260 89518 29262 89570
rect 29314 89518 29316 89570
rect 29260 89124 29316 89518
rect 29260 89058 29316 89068
rect 29932 88340 29988 88350
rect 30044 88340 30100 90300
rect 30156 90290 30212 90300
rect 30268 90018 30324 90526
rect 30268 89966 30270 90018
rect 30322 89966 30324 90018
rect 30268 89954 30324 89966
rect 30492 89906 30548 89918
rect 30492 89854 30494 89906
rect 30546 89854 30548 89906
rect 30380 89794 30436 89806
rect 30380 89742 30382 89794
rect 30434 89742 30436 89794
rect 30156 88900 30212 88910
rect 30212 88844 30324 88900
rect 30156 88806 30212 88844
rect 29932 88338 30100 88340
rect 29932 88286 29934 88338
rect 29986 88286 30100 88338
rect 29932 88284 30100 88286
rect 29932 88274 29988 88284
rect 28588 88228 28644 88238
rect 28588 88134 28644 88172
rect 29260 88228 29316 88238
rect 29260 88134 29316 88172
rect 28084 86940 28532 86996
rect 29148 88004 29204 88014
rect 28028 86658 28084 86940
rect 29148 86770 29204 87948
rect 29148 86718 29150 86770
rect 29202 86718 29204 86770
rect 28028 86606 28030 86658
rect 28082 86606 28084 86658
rect 28028 86594 28084 86606
rect 28476 86658 28532 86670
rect 28476 86606 28478 86658
rect 28530 86606 28532 86658
rect 27692 86548 27748 86558
rect 27692 86436 27748 86492
rect 27804 86436 27860 86446
rect 27692 86434 27860 86436
rect 27692 86382 27806 86434
rect 27858 86382 27860 86434
rect 27692 86380 27860 86382
rect 27692 82292 27748 86380
rect 27804 86370 27860 86380
rect 27916 86436 27972 86446
rect 27916 86342 27972 86380
rect 28476 85652 28532 86606
rect 28924 85764 28980 85774
rect 28924 85652 29092 85708
rect 28364 84866 28420 84878
rect 28364 84814 28366 84866
rect 28418 84814 28420 84866
rect 28028 84532 28084 84542
rect 28028 84418 28084 84476
rect 28028 84366 28030 84418
rect 28082 84366 28084 84418
rect 28028 84354 28084 84366
rect 27804 84306 27860 84318
rect 27804 84254 27806 84306
rect 27858 84254 27860 84306
rect 27804 83748 27860 84254
rect 28252 84084 28308 84094
rect 27804 83682 27860 83692
rect 28140 84082 28308 84084
rect 28140 84030 28254 84082
rect 28306 84030 28308 84082
rect 28140 84028 28308 84030
rect 27692 82226 27748 82236
rect 27916 82738 27972 82750
rect 27916 82686 27918 82738
rect 27970 82686 27972 82738
rect 27804 82068 27860 82078
rect 27804 81394 27860 82012
rect 27804 81342 27806 81394
rect 27858 81342 27860 81394
rect 27804 81330 27860 81342
rect 27916 81954 27972 82686
rect 28028 82516 28084 82526
rect 28140 82516 28196 84028
rect 28252 84018 28308 84028
rect 28364 83636 28420 84814
rect 28476 84420 28532 85596
rect 29036 84756 29092 85652
rect 29148 85204 29204 86718
rect 29484 87892 29540 87902
rect 29260 86436 29316 86446
rect 29260 86434 29428 86436
rect 29260 86382 29262 86434
rect 29314 86382 29428 86434
rect 29260 86380 29428 86382
rect 29260 86370 29316 86380
rect 29148 85138 29204 85148
rect 29372 85090 29428 86380
rect 29484 85202 29540 87836
rect 29596 86772 29652 86782
rect 29596 86678 29652 86716
rect 29484 85150 29486 85202
rect 29538 85150 29540 85202
rect 29484 85138 29540 85150
rect 29932 85876 29988 85886
rect 29932 85202 29988 85820
rect 30268 85874 30324 88844
rect 30380 87444 30436 89742
rect 30492 87668 30548 89854
rect 31052 88898 31108 88910
rect 31052 88846 31054 88898
rect 31106 88846 31108 88898
rect 31052 88228 31108 88846
rect 31052 88162 31108 88172
rect 32060 88338 32116 88350
rect 32060 88286 32062 88338
rect 32114 88286 32116 88338
rect 32060 87668 32116 88286
rect 30492 87612 31220 87668
rect 31164 87554 31220 87612
rect 32060 87602 32116 87612
rect 32508 88228 32564 88238
rect 32508 88002 32564 88172
rect 32508 87950 32510 88002
rect 32562 87950 32564 88002
rect 31164 87502 31166 87554
rect 31218 87502 31220 87554
rect 30380 87378 30436 87388
rect 30828 87442 30884 87454
rect 30828 87390 30830 87442
rect 30882 87390 30884 87442
rect 30268 85822 30270 85874
rect 30322 85822 30324 85874
rect 30268 85810 30324 85822
rect 30828 86772 30884 87390
rect 29932 85150 29934 85202
rect 29986 85150 29988 85202
rect 29932 85138 29988 85150
rect 30716 85764 30772 85774
rect 30828 85764 30884 86716
rect 30772 85708 30884 85764
rect 31052 87444 31108 87454
rect 31052 85708 31108 87388
rect 31164 85876 31220 87502
rect 32060 87444 32116 87454
rect 31612 87220 31668 87230
rect 31612 87218 32004 87220
rect 31612 87166 31614 87218
rect 31666 87166 32004 87218
rect 31612 87164 32004 87166
rect 31612 87154 31668 87164
rect 31724 86546 31780 86558
rect 31724 86494 31726 86546
rect 31778 86494 31780 86546
rect 31164 85782 31220 85820
rect 31388 86268 31668 86324
rect 31388 85708 31444 86268
rect 29372 85038 29374 85090
rect 29426 85038 29428 85090
rect 29372 85026 29428 85038
rect 30380 84866 30436 84878
rect 30380 84814 30382 84866
rect 30434 84814 30436 84866
rect 30156 84756 30212 84766
rect 29036 84700 29316 84756
rect 28588 84532 28644 84542
rect 29148 84532 29204 84542
rect 28588 84530 29204 84532
rect 28588 84478 28590 84530
rect 28642 84478 29150 84530
rect 29202 84478 29204 84530
rect 28588 84476 29204 84478
rect 28588 84466 28644 84476
rect 29148 84466 29204 84476
rect 28476 84354 28532 84364
rect 28476 84084 28532 84094
rect 28476 83748 28532 84028
rect 29260 83972 29316 84700
rect 29148 83916 29316 83972
rect 29372 84644 29428 84654
rect 28476 83692 28756 83748
rect 28420 83580 28532 83636
rect 28364 83570 28420 83580
rect 28364 83300 28420 83310
rect 28084 82460 28196 82516
rect 28252 82962 28308 82974
rect 28252 82910 28254 82962
rect 28306 82910 28308 82962
rect 28028 82450 28084 82460
rect 27916 81902 27918 81954
rect 27970 81902 27972 81954
rect 27692 81284 27748 81294
rect 27692 81190 27748 81228
rect 27916 81170 27972 81902
rect 28140 81730 28196 81742
rect 28140 81678 28142 81730
rect 28194 81678 28196 81730
rect 28140 81508 28196 81678
rect 28140 81442 28196 81452
rect 27916 81118 27918 81170
rect 27970 81118 27972 81170
rect 27580 80668 27860 80724
rect 27692 80498 27748 80510
rect 27692 80446 27694 80498
rect 27746 80446 27748 80498
rect 27692 79716 27748 80446
rect 27692 79650 27748 79660
rect 27692 79380 27748 79390
rect 27580 79044 27636 79054
rect 27468 78988 27580 79044
rect 27580 78978 27636 78988
rect 27020 78754 27076 78764
rect 27132 78932 27188 78942
rect 27132 78706 27188 78876
rect 27356 78930 27412 78942
rect 27356 78878 27358 78930
rect 27410 78878 27412 78930
rect 27244 78820 27300 78830
rect 27244 78726 27300 78764
rect 27132 78654 27134 78706
rect 27186 78654 27188 78706
rect 27132 78642 27188 78654
rect 26684 78034 26740 78540
rect 26684 77982 26686 78034
rect 26738 77982 26740 78034
rect 26348 77756 26516 77812
rect 26572 77922 26628 77934
rect 26572 77870 26574 77922
rect 26626 77870 26628 77922
rect 26348 76916 26404 77756
rect 26572 77252 26628 77870
rect 26684 77588 26740 77982
rect 27020 77922 27076 77934
rect 27020 77870 27022 77922
rect 27074 77870 27076 77922
rect 27020 77700 27076 77870
rect 27244 77812 27300 77822
rect 27020 77634 27076 77644
rect 27132 77756 27244 77812
rect 26684 77522 26740 77532
rect 27020 77476 27076 77486
rect 26908 77252 26964 77262
rect 26572 77250 26964 77252
rect 26572 77198 26910 77250
rect 26962 77198 26964 77250
rect 26572 77196 26964 77198
rect 26908 77186 26964 77196
rect 27020 77028 27076 77420
rect 26348 76850 26404 76860
rect 26908 76972 27076 77028
rect 27132 77026 27188 77756
rect 27244 77718 27300 77756
rect 27356 77588 27412 78878
rect 27692 78818 27748 79324
rect 27692 78766 27694 78818
rect 27746 78766 27748 78818
rect 27692 78754 27748 78766
rect 27244 77532 27412 77588
rect 27468 78596 27524 78606
rect 27804 78596 27860 80668
rect 27916 80500 27972 81118
rect 28252 81170 28308 82910
rect 28364 82850 28420 83244
rect 28364 82798 28366 82850
rect 28418 82798 28420 82850
rect 28364 82786 28420 82798
rect 28364 81956 28420 81966
rect 28476 81956 28532 83580
rect 28364 81954 28532 81956
rect 28364 81902 28366 81954
rect 28418 81902 28532 81954
rect 28364 81900 28532 81902
rect 28588 82738 28644 82750
rect 28588 82686 28590 82738
rect 28642 82686 28644 82738
rect 28588 81954 28644 82686
rect 28588 81902 28590 81954
rect 28642 81902 28644 81954
rect 28364 81732 28420 81900
rect 28588 81844 28644 81902
rect 28588 81778 28644 81788
rect 28364 81666 28420 81676
rect 28700 81620 28756 83692
rect 29036 83524 29092 83534
rect 28924 83522 29092 83524
rect 28924 83470 29038 83522
rect 29090 83470 29092 83522
rect 28924 83468 29092 83470
rect 28812 82738 28868 82750
rect 28812 82686 28814 82738
rect 28866 82686 28868 82738
rect 28812 82180 28868 82686
rect 28924 82628 28980 83468
rect 29036 83458 29092 83468
rect 29148 83076 29204 83916
rect 29260 83748 29316 83758
rect 29260 83654 29316 83692
rect 29372 83300 29428 84588
rect 30156 84530 30212 84700
rect 30156 84478 30158 84530
rect 30210 84478 30212 84530
rect 30156 84466 30212 84478
rect 29708 84420 29764 84430
rect 29708 84326 29764 84364
rect 29596 83412 29652 83422
rect 29596 83318 29652 83356
rect 30044 83300 30100 83310
rect 29372 83298 29540 83300
rect 29372 83246 29374 83298
rect 29426 83246 29540 83298
rect 29372 83244 29540 83246
rect 29372 83234 29428 83244
rect 29148 83020 29316 83076
rect 29036 82964 29092 82974
rect 29036 82870 29092 82908
rect 29148 82852 29204 82862
rect 29148 82738 29204 82796
rect 29148 82686 29150 82738
rect 29202 82686 29204 82738
rect 29148 82674 29204 82686
rect 28924 82562 28980 82572
rect 28812 82114 28868 82124
rect 28476 81564 28756 81620
rect 28476 81396 28532 81564
rect 28252 81118 28254 81170
rect 28306 81118 28308 81170
rect 28252 81106 28308 81118
rect 28364 81340 28532 81396
rect 27916 80444 28308 80500
rect 27916 80274 27972 80286
rect 27916 80222 27918 80274
rect 27970 80222 27972 80274
rect 27916 78932 27972 80222
rect 28140 80274 28196 80286
rect 28140 80222 28142 80274
rect 28194 80222 28196 80274
rect 27916 78866 27972 78876
rect 28028 78930 28084 78942
rect 28028 78878 28030 78930
rect 28082 78878 28084 78930
rect 28028 78820 28084 78878
rect 28140 78932 28196 80222
rect 28140 78866 28196 78876
rect 28252 80162 28308 80444
rect 28252 80110 28254 80162
rect 28306 80110 28308 80162
rect 28028 78754 28084 78764
rect 27244 77250 27300 77532
rect 27468 77476 27524 78540
rect 27692 78540 27860 78596
rect 28252 78596 28308 80110
rect 28364 79044 28420 81340
rect 28700 81282 28756 81294
rect 28700 81230 28702 81282
rect 28754 81230 28756 81282
rect 28476 81172 28532 81210
rect 28476 81106 28532 81116
rect 28476 80948 28532 80958
rect 28476 80386 28532 80892
rect 28476 80334 28478 80386
rect 28530 80334 28532 80386
rect 28476 80322 28532 80334
rect 28364 78988 28532 79044
rect 27580 78260 27636 78270
rect 27692 78260 27748 78540
rect 28252 78530 28308 78540
rect 28364 78820 28420 78830
rect 27580 78258 27748 78260
rect 27580 78206 27582 78258
rect 27634 78206 27748 78258
rect 27580 78204 27748 78206
rect 27580 78194 27636 78204
rect 28028 77924 28084 77934
rect 28028 77830 28084 77868
rect 27468 77420 27972 77476
rect 27244 77198 27246 77250
rect 27298 77198 27300 77250
rect 27244 77186 27300 77198
rect 27356 77250 27412 77262
rect 27356 77198 27358 77250
rect 27410 77198 27412 77250
rect 27132 76974 27134 77026
rect 27186 76974 27188 77026
rect 26236 76638 26238 76690
rect 26290 76638 26292 76690
rect 26236 75348 26292 76638
rect 26796 76692 26852 76702
rect 26796 76580 26852 76636
rect 26684 76578 26852 76580
rect 26684 76526 26798 76578
rect 26850 76526 26852 76578
rect 26684 76524 26852 76526
rect 26236 75282 26292 75292
rect 26348 75908 26404 75918
rect 26124 74062 26126 74114
rect 26178 74062 26180 74114
rect 26124 74050 26180 74062
rect 26236 73556 26292 73566
rect 26012 73554 26292 73556
rect 26012 73502 26238 73554
rect 26290 73502 26292 73554
rect 26012 73500 26292 73502
rect 26236 73490 26292 73500
rect 26124 73330 26180 73342
rect 26124 73278 26126 73330
rect 26178 73278 26180 73330
rect 26124 73108 26180 73278
rect 26236 73220 26292 73230
rect 26236 73126 26292 73164
rect 26124 73042 26180 73052
rect 25900 72716 26180 72772
rect 25564 71762 25620 72716
rect 26124 71986 26180 72716
rect 26124 71934 26126 71986
rect 26178 71934 26180 71986
rect 26124 71922 26180 71934
rect 26236 71988 26292 71998
rect 26348 71988 26404 75852
rect 26684 75908 26740 76524
rect 26796 76514 26852 76524
rect 26684 75842 26740 75852
rect 26796 76244 26852 76254
rect 26460 75010 26516 75022
rect 26460 74958 26462 75010
rect 26514 74958 26516 75010
rect 26460 74900 26516 74958
rect 26460 74834 26516 74844
rect 26796 74898 26852 76188
rect 26796 74846 26798 74898
rect 26850 74846 26852 74898
rect 26796 74834 26852 74846
rect 26908 73948 26964 76972
rect 27132 76962 27188 76974
rect 27356 77028 27412 77198
rect 27804 77028 27860 77038
rect 27356 76962 27412 76972
rect 27692 77026 27860 77028
rect 27692 76974 27806 77026
rect 27858 76974 27860 77026
rect 27692 76972 27860 76974
rect 27692 76804 27748 76972
rect 27804 76962 27860 76972
rect 27020 76748 27748 76804
rect 27804 76804 27860 76814
rect 27020 76578 27076 76748
rect 27804 76690 27860 76748
rect 27804 76638 27806 76690
rect 27858 76638 27860 76690
rect 27020 76526 27022 76578
rect 27074 76526 27076 76578
rect 27020 76514 27076 76526
rect 27132 76578 27188 76590
rect 27132 76526 27134 76578
rect 27186 76526 27188 76578
rect 27132 76356 27188 76526
rect 27244 76580 27300 76590
rect 27244 76486 27300 76524
rect 27468 76580 27524 76590
rect 27356 76468 27412 76478
rect 27356 76374 27412 76412
rect 27020 76300 27132 76356
rect 27020 74900 27076 76300
rect 27132 76262 27188 76300
rect 27468 75122 27524 76524
rect 27580 76466 27636 76478
rect 27580 76414 27582 76466
rect 27634 76414 27636 76466
rect 27580 75684 27636 76414
rect 27804 75796 27860 76638
rect 27916 76466 27972 77420
rect 28140 77364 28196 77374
rect 28364 77364 28420 78764
rect 28476 78260 28532 78988
rect 28700 78820 28756 81230
rect 29260 81284 29316 83020
rect 29372 82740 29428 82750
rect 29372 82646 29428 82684
rect 29484 82628 29540 83244
rect 30044 83206 30100 83244
rect 30156 83076 30212 83086
rect 29820 82628 29876 82638
rect 29484 82626 29876 82628
rect 29484 82574 29822 82626
rect 29874 82574 29876 82626
rect 29484 82572 29876 82574
rect 29596 81730 29652 81742
rect 29596 81678 29598 81730
rect 29650 81678 29652 81730
rect 29596 81284 29652 81678
rect 29708 81732 29764 82572
rect 29820 82562 29876 82572
rect 30156 82628 30212 83020
rect 30156 82626 30324 82628
rect 30156 82574 30158 82626
rect 30210 82574 30324 82626
rect 30156 82572 30324 82574
rect 30156 82562 30212 82572
rect 29708 81666 29764 81676
rect 29820 82404 29876 82414
rect 29260 81228 29428 81284
rect 28812 81172 28868 81182
rect 29036 81172 29092 81182
rect 28812 81170 29092 81172
rect 28812 81118 28814 81170
rect 28866 81118 29038 81170
rect 29090 81118 29092 81170
rect 28812 81116 29092 81118
rect 28812 81106 28868 81116
rect 29036 81106 29092 81116
rect 29260 81060 29316 81070
rect 29260 80966 29316 81004
rect 29260 80500 29316 80510
rect 29372 80500 29428 81228
rect 29596 81218 29652 81228
rect 29596 80948 29652 80958
rect 29596 80946 29764 80948
rect 29596 80894 29598 80946
rect 29650 80894 29764 80946
rect 29596 80892 29764 80894
rect 29596 80882 29652 80892
rect 29708 80610 29764 80892
rect 29708 80558 29710 80610
rect 29762 80558 29764 80610
rect 29708 80546 29764 80558
rect 28700 78754 28756 78764
rect 28812 80498 29428 80500
rect 28812 80446 29262 80498
rect 29314 80446 29428 80498
rect 28812 80444 29428 80446
rect 28588 78706 28644 78718
rect 28588 78654 28590 78706
rect 28642 78654 28644 78706
rect 28588 78596 28644 78654
rect 28812 78596 28868 80444
rect 29260 80434 29316 80444
rect 29372 79492 29428 79502
rect 29148 78932 29204 78942
rect 29148 78838 29204 78876
rect 28588 78540 28868 78596
rect 28812 78260 28868 78540
rect 28476 78204 28644 78260
rect 28476 78036 28532 78046
rect 28476 77942 28532 77980
rect 28588 77812 28644 78204
rect 28812 78194 28868 78204
rect 29148 78596 29204 78606
rect 29148 78258 29204 78540
rect 29148 78206 29150 78258
rect 29202 78206 29204 78258
rect 29148 78194 29204 78206
rect 29260 78260 29316 78270
rect 29260 78166 29316 78204
rect 29372 78258 29428 79436
rect 29708 78932 29764 78942
rect 29708 78838 29764 78876
rect 29484 78820 29540 78830
rect 29484 78726 29540 78764
rect 29372 78206 29374 78258
rect 29426 78206 29428 78258
rect 29372 78194 29428 78206
rect 29484 78036 29540 78046
rect 27916 76414 27918 76466
rect 27970 76414 27972 76466
rect 27916 76356 27972 76414
rect 27916 76290 27972 76300
rect 28028 77362 28420 77364
rect 28028 77310 28142 77362
rect 28194 77310 28420 77362
rect 28028 77308 28420 77310
rect 28476 77756 28644 77812
rect 29372 78034 29540 78036
rect 29372 77982 29486 78034
rect 29538 77982 29540 78034
rect 29372 77980 29540 77982
rect 27804 75730 27860 75740
rect 27580 75618 27636 75628
rect 27468 75070 27470 75122
rect 27522 75070 27524 75122
rect 27468 75058 27524 75070
rect 27804 75348 27860 75358
rect 27020 74834 27076 74844
rect 27132 75012 27188 75022
rect 27132 73948 27188 74956
rect 27580 74898 27636 74910
rect 27580 74846 27582 74898
rect 27634 74846 27636 74898
rect 26908 73892 27076 73948
rect 27132 73892 27300 73948
rect 26908 73330 26964 73342
rect 26908 73278 26910 73330
rect 26962 73278 26964 73330
rect 26908 73108 26964 73278
rect 26908 73042 26964 73052
rect 26236 71986 26404 71988
rect 26236 71934 26238 71986
rect 26290 71934 26404 71986
rect 26236 71932 26404 71934
rect 26796 72436 26852 72446
rect 26236 71922 26292 71932
rect 25564 71710 25566 71762
rect 25618 71710 25620 71762
rect 25564 71698 25620 71710
rect 26012 71762 26068 71774
rect 26012 71710 26014 71762
rect 26066 71710 26068 71762
rect 25788 71652 25844 71662
rect 26012 71652 26068 71710
rect 25788 71650 25956 71652
rect 25788 71598 25790 71650
rect 25842 71598 25956 71650
rect 25788 71596 25956 71598
rect 25788 71586 25844 71596
rect 25452 70702 25454 70754
rect 25506 70702 25508 70754
rect 25452 70690 25508 70702
rect 25564 70980 25620 70990
rect 25564 70588 25620 70924
rect 25788 70866 25844 70878
rect 25788 70814 25790 70866
rect 25842 70814 25844 70866
rect 25564 70532 25732 70588
rect 25340 70420 25396 70430
rect 25228 70364 25340 70420
rect 24444 69300 24500 69310
rect 24332 69298 24500 69300
rect 24332 69246 24446 69298
rect 24498 69246 24500 69298
rect 24332 69244 24500 69246
rect 24108 67954 24164 67966
rect 24108 67902 24110 67954
rect 24162 67902 24164 67954
rect 23212 65716 23268 66892
rect 23100 65660 23268 65716
rect 23436 66946 23492 66958
rect 23884 66948 23940 66958
rect 23436 66894 23438 66946
rect 23490 66894 23492 66946
rect 22876 65202 22932 65212
rect 22988 65490 23044 65502
rect 22988 65438 22990 65490
rect 23042 65438 23044 65490
rect 22988 64930 23044 65438
rect 22988 64878 22990 64930
rect 23042 64878 23044 64930
rect 22988 64866 23044 64878
rect 21868 64818 22148 64820
rect 21868 64766 22094 64818
rect 22146 64766 22148 64818
rect 21868 64764 22148 64766
rect 21868 64036 21924 64764
rect 22092 64754 22148 64764
rect 22540 64596 22596 64606
rect 22540 64502 22596 64540
rect 21868 63026 21924 63980
rect 22988 63922 23044 63934
rect 22988 63870 22990 63922
rect 23042 63870 23044 63922
rect 22876 63140 22932 63150
rect 21868 62974 21870 63026
rect 21922 62974 21924 63026
rect 21868 62962 21924 62974
rect 22204 63028 22260 63038
rect 21532 62132 21812 62188
rect 21420 61684 21476 61694
rect 21420 61590 21476 61628
rect 21308 61068 21476 61124
rect 21420 60898 21476 61068
rect 21420 60846 21422 60898
rect 21474 60846 21476 60898
rect 21420 60834 21476 60846
rect 21196 60788 21252 60798
rect 21196 60694 21252 60732
rect 21084 60386 21140 60396
rect 20636 60274 20692 60284
rect 21532 60116 21588 62132
rect 21756 61684 21812 61694
rect 21756 61570 21812 61628
rect 21756 61518 21758 61570
rect 21810 61518 21812 61570
rect 21756 61506 21812 61518
rect 21644 60674 21700 60686
rect 21644 60622 21646 60674
rect 21698 60622 21700 60674
rect 21644 60452 21700 60622
rect 21700 60396 21924 60452
rect 21644 60358 21700 60396
rect 20636 60060 21588 60116
rect 20636 60002 20692 60060
rect 20636 59950 20638 60002
rect 20690 59950 20692 60002
rect 20636 59938 20692 59950
rect 21308 59890 21364 59902
rect 21308 59838 21310 59890
rect 21362 59838 21364 59890
rect 21308 59780 21364 59838
rect 21532 59890 21588 60060
rect 21644 60116 21700 60126
rect 21644 60114 21812 60116
rect 21644 60062 21646 60114
rect 21698 60062 21812 60114
rect 21644 60060 21812 60062
rect 21644 60050 21700 60060
rect 21532 59838 21534 59890
rect 21586 59838 21588 59890
rect 21532 59826 21588 59838
rect 20524 59724 21364 59780
rect 20972 59106 21028 59118
rect 20972 59054 20974 59106
rect 21026 59054 21028 59106
rect 20748 58548 20804 58558
rect 20412 57486 20414 57538
rect 20466 57486 20468 57538
rect 20412 57474 20468 57486
rect 20524 58546 20804 58548
rect 20524 58494 20750 58546
rect 20802 58494 20804 58546
rect 20524 58492 20804 58494
rect 20300 54402 20356 54414
rect 20300 54350 20302 54402
rect 20354 54350 20356 54402
rect 20300 53620 20356 54350
rect 20412 53732 20468 53742
rect 20412 53638 20468 53676
rect 20300 53554 20356 53564
rect 20188 53228 20356 53284
rect 20076 52948 20132 52958
rect 19964 52946 20132 52948
rect 19964 52894 20078 52946
rect 20130 52894 20132 52946
rect 19964 52892 20132 52894
rect 19964 52500 20020 52892
rect 20076 52882 20132 52892
rect 19964 52052 20020 52444
rect 20076 52164 20132 52174
rect 20076 52070 20132 52108
rect 20188 52162 20244 52174
rect 20188 52110 20190 52162
rect 20242 52110 20244 52162
rect 19964 51986 20020 51996
rect 18508 44158 18510 44210
rect 18562 44158 18564 44210
rect 18508 41412 18564 44158
rect 18844 44100 18900 51884
rect 19068 51884 19684 51940
rect 19068 47572 19124 51884
rect 19836 51772 20100 51782
rect 19180 51716 19236 51726
rect 19180 51378 19236 51660
rect 19628 51716 19684 51726
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 19836 51706 20100 51716
rect 19516 51604 19572 51614
rect 19180 51326 19182 51378
rect 19234 51326 19236 51378
rect 19180 51156 19236 51326
rect 19180 51090 19236 51100
rect 19292 51490 19348 51502
rect 19292 51438 19294 51490
rect 19346 51438 19348 51490
rect 19292 50428 19348 51438
rect 18396 41356 18564 41412
rect 18620 44044 18900 44100
rect 18956 47516 19124 47572
rect 19180 50372 19348 50428
rect 19404 51380 19460 51390
rect 19180 49698 19236 50372
rect 19404 50036 19460 51324
rect 19516 50484 19572 51548
rect 19516 50418 19572 50428
rect 19404 49942 19460 49980
rect 19180 49646 19182 49698
rect 19234 49646 19236 49698
rect 18396 40852 18452 41356
rect 18508 41186 18564 41198
rect 18508 41134 18510 41186
rect 18562 41134 18564 41186
rect 18508 41076 18564 41134
rect 18508 41010 18564 41020
rect 18396 40796 18564 40852
rect 18508 40740 18564 40796
rect 18508 40516 18564 40684
rect 18508 39730 18564 40460
rect 18508 39678 18510 39730
rect 18562 39678 18564 39730
rect 18508 39666 18564 39678
rect 18620 39396 18676 44044
rect 18956 43988 19012 47516
rect 19068 47346 19124 47358
rect 19068 47294 19070 47346
rect 19122 47294 19124 47346
rect 19068 47236 19124 47294
rect 19068 47170 19124 47180
rect 18508 39340 18676 39396
rect 18732 43932 19012 43988
rect 19068 46004 19124 46014
rect 19068 45780 19124 45948
rect 19068 45108 19124 45724
rect 19180 45332 19236 49646
rect 19404 49252 19460 49262
rect 19404 48580 19460 49196
rect 19404 48466 19460 48524
rect 19404 48414 19406 48466
rect 19458 48414 19460 48466
rect 19404 48402 19460 48414
rect 19404 46786 19460 46798
rect 19404 46734 19406 46786
rect 19458 46734 19460 46786
rect 19404 46340 19460 46734
rect 19516 46676 19572 46686
rect 19516 46582 19572 46620
rect 19404 45444 19460 46284
rect 19404 45378 19460 45388
rect 19180 45276 19348 45332
rect 19180 45108 19236 45118
rect 19068 45106 19236 45108
rect 19068 45054 19182 45106
rect 19234 45054 19236 45106
rect 19068 45052 19236 45054
rect 18396 39060 18452 39070
rect 18396 38966 18452 39004
rect 18284 38434 18340 38444
rect 18396 38610 18452 38622
rect 18396 38558 18398 38610
rect 18450 38558 18452 38610
rect 18396 38162 18452 38558
rect 18396 38110 18398 38162
rect 18450 38110 18452 38162
rect 18396 38098 18452 38110
rect 18284 37492 18340 37502
rect 18284 37398 18340 37436
rect 18508 36596 18564 39340
rect 18620 38836 18676 38846
rect 18620 38722 18676 38780
rect 18620 38670 18622 38722
rect 18674 38670 18676 38722
rect 18620 38658 18676 38670
rect 18732 37492 18788 43932
rect 19068 43652 19124 45052
rect 19180 45042 19236 45052
rect 19292 44884 19348 45276
rect 19068 43586 19124 43596
rect 19180 44828 19348 44884
rect 19068 43204 19124 43214
rect 19068 42642 19124 43148
rect 19068 42590 19070 42642
rect 19122 42590 19124 42642
rect 19068 42578 19124 42590
rect 19180 42420 19236 44828
rect 19068 42364 19236 42420
rect 19292 43762 19348 43774
rect 19292 43710 19294 43762
rect 19346 43710 19348 43762
rect 18956 42196 19012 42206
rect 18732 37426 18788 37436
rect 18844 42194 19012 42196
rect 18844 42142 18958 42194
rect 19010 42142 19012 42194
rect 18844 42140 19012 42142
rect 18508 36502 18564 36540
rect 18620 37380 18676 37390
rect 18620 35700 18676 37324
rect 18620 35634 18676 35644
rect 18732 35588 18788 35598
rect 18732 35494 18788 35532
rect 18396 35476 18452 35486
rect 18620 35476 18676 35486
rect 18396 35382 18452 35420
rect 18508 35474 18676 35476
rect 18508 35422 18622 35474
rect 18674 35422 18676 35474
rect 18508 35420 18676 35422
rect 18172 34962 18228 34972
rect 18284 35364 18340 35374
rect 17388 34514 17444 34524
rect 17500 34916 17556 34926
rect 17836 34916 17892 34926
rect 17388 34132 17444 34142
rect 17276 34130 17444 34132
rect 17276 34078 17390 34130
rect 17442 34078 17444 34130
rect 17276 34076 17444 34078
rect 17276 32788 17332 34076
rect 17388 34066 17444 34076
rect 17388 33572 17444 33582
rect 17388 33458 17444 33516
rect 17388 33406 17390 33458
rect 17442 33406 17444 33458
rect 17388 33394 17444 33406
rect 17500 33124 17556 34860
rect 17724 34914 17892 34916
rect 17724 34862 17838 34914
rect 17890 34862 17892 34914
rect 17724 34860 17892 34862
rect 17724 34354 17780 34860
rect 17836 34850 17892 34860
rect 17724 34302 17726 34354
rect 17778 34302 17780 34354
rect 17724 34290 17780 34302
rect 18060 34802 18116 34814
rect 18060 34750 18062 34802
rect 18114 34750 18116 34802
rect 18060 34356 18116 34750
rect 18172 34804 18228 34814
rect 18172 34710 18228 34748
rect 18060 34290 18116 34300
rect 17612 34130 17668 34142
rect 17612 34078 17614 34130
rect 17666 34078 17668 34130
rect 17612 33908 17668 34078
rect 17612 33842 17668 33852
rect 17836 34130 17892 34142
rect 17836 34078 17838 34130
rect 17890 34078 17892 34130
rect 17836 33572 17892 34078
rect 17948 34130 18004 34142
rect 17948 34078 17950 34130
rect 18002 34078 18004 34130
rect 17948 34020 18004 34078
rect 17948 33954 18004 33964
rect 17892 33516 18004 33572
rect 17836 33506 17892 33516
rect 17276 32722 17332 32732
rect 17388 33068 17556 33124
rect 17612 33460 17668 33470
rect 17388 29652 17444 33068
rect 17500 32900 17556 32910
rect 17500 32786 17556 32844
rect 17500 32734 17502 32786
rect 17554 32734 17556 32786
rect 17500 32722 17556 32734
rect 17612 32340 17668 33404
rect 17836 33346 17892 33358
rect 17836 33294 17838 33346
rect 17890 33294 17892 33346
rect 17836 32900 17892 33294
rect 17836 32834 17892 32844
rect 17836 32564 17892 32574
rect 17948 32564 18004 33516
rect 17836 32562 18004 32564
rect 17836 32510 17838 32562
rect 17890 32510 18004 32562
rect 17836 32508 18004 32510
rect 17836 32498 17892 32508
rect 17612 31890 17668 32284
rect 18060 32340 18116 32350
rect 18060 32246 18116 32284
rect 17612 31838 17614 31890
rect 17666 31838 17668 31890
rect 17612 31826 17668 31838
rect 18060 30772 18116 30782
rect 17500 29652 17556 29662
rect 17444 29650 17668 29652
rect 17444 29598 17502 29650
rect 17554 29598 17668 29650
rect 17444 29596 17668 29598
rect 17388 29558 17444 29596
rect 17500 29586 17556 29596
rect 17612 28084 17668 29596
rect 17948 28532 18004 28542
rect 17612 27990 17668 28028
rect 17836 28196 17892 28206
rect 17836 28082 17892 28140
rect 17836 28030 17838 28082
rect 17890 28030 17892 28082
rect 17724 27972 17780 27982
rect 17724 27878 17780 27916
rect 17388 27860 17444 27870
rect 17388 27766 17444 27804
rect 17500 27412 17556 27422
rect 17556 27356 17780 27412
rect 17500 27346 17556 27356
rect 17052 27132 17220 27188
rect 17724 27186 17780 27356
rect 17724 27134 17726 27186
rect 17778 27134 17780 27186
rect 16940 27076 16996 27114
rect 16716 26786 16772 26796
rect 16828 27020 16940 27076
rect 16604 26450 16660 26460
rect 16828 26514 16884 27020
rect 16940 27010 16996 27020
rect 17052 26908 17108 27132
rect 17724 27122 17780 27134
rect 16828 26462 16830 26514
rect 16882 26462 16884 26514
rect 16492 26236 16772 26292
rect 16380 26178 16548 26180
rect 16380 26126 16382 26178
rect 16434 26126 16548 26178
rect 16380 26124 16548 26126
rect 16380 26114 16436 26124
rect 15484 25396 15540 26012
rect 16156 26068 16212 26078
rect 16156 25974 16212 26012
rect 15484 25330 15540 25340
rect 15484 23940 15540 23950
rect 16268 23940 16324 23950
rect 15484 22372 15540 23884
rect 15596 23938 16324 23940
rect 15596 23886 16270 23938
rect 16322 23886 16324 23938
rect 15596 23884 16324 23886
rect 15596 22482 15652 23884
rect 16268 23874 16324 23884
rect 16380 23826 16436 23838
rect 16380 23774 16382 23826
rect 16434 23774 16436 23826
rect 15596 22430 15598 22482
rect 15650 22430 15652 22482
rect 15596 22418 15652 22430
rect 15820 23716 15876 23726
rect 15484 22306 15540 22316
rect 15484 22146 15540 22158
rect 15484 22094 15486 22146
rect 15538 22094 15540 22146
rect 15484 21252 15540 22094
rect 15708 22148 15764 22158
rect 15708 22054 15764 22092
rect 15820 21812 15876 23660
rect 16268 23604 16324 23614
rect 16268 23044 16324 23548
rect 15932 23042 16324 23044
rect 15932 22990 16270 23042
rect 16322 22990 16324 23042
rect 15932 22988 16324 22990
rect 15932 22370 15988 22988
rect 16268 22978 16324 22988
rect 16380 22708 16436 23774
rect 16492 23044 16548 26124
rect 16716 23716 16772 26236
rect 16716 23650 16772 23660
rect 16716 23380 16772 23390
rect 16828 23380 16884 26462
rect 16940 26852 17108 26908
rect 17164 26964 17220 26974
rect 16940 24050 16996 26852
rect 17052 26068 17108 26078
rect 17052 25618 17108 26012
rect 17052 25566 17054 25618
rect 17106 25566 17108 25618
rect 17052 25554 17108 25566
rect 16940 23998 16942 24050
rect 16994 23998 16996 24050
rect 16940 23986 16996 23998
rect 17164 23548 17220 26908
rect 17836 26908 17892 28030
rect 17948 28082 18004 28476
rect 17948 28030 17950 28082
rect 18002 28030 18004 28082
rect 17948 28018 18004 28030
rect 17836 26852 18004 26908
rect 16716 23378 16884 23380
rect 16716 23326 16718 23378
rect 16770 23326 16884 23378
rect 16716 23324 16884 23326
rect 17052 23492 17220 23548
rect 17276 26740 17332 26750
rect 16716 23268 16772 23324
rect 16716 23202 16772 23212
rect 16828 23044 16884 23054
rect 16492 22988 16772 23044
rect 15932 22318 15934 22370
rect 15986 22318 15988 22370
rect 15932 22306 15988 22318
rect 16044 22652 16436 22708
rect 15932 21812 15988 21822
rect 15820 21810 15988 21812
rect 15820 21758 15934 21810
rect 15986 21758 15988 21810
rect 15820 21756 15988 21758
rect 15708 21588 15764 21598
rect 15484 21186 15540 21196
rect 15596 21586 15764 21588
rect 15596 21534 15710 21586
rect 15762 21534 15764 21586
rect 15596 21532 15764 21534
rect 15372 18274 15428 18284
rect 13692 17668 13748 17678
rect 13356 17612 13524 17668
rect 13580 17666 13748 17668
rect 13580 17614 13694 17666
rect 13746 17614 13748 17666
rect 13580 17612 13748 17614
rect 13356 17556 13412 17612
rect 13356 17490 13412 17500
rect 13468 17444 13524 17454
rect 13468 17350 13524 17388
rect 13468 16324 13524 16334
rect 13580 16324 13636 17612
rect 13692 17602 13748 17612
rect 14476 17556 14532 17566
rect 14476 17554 14868 17556
rect 14476 17502 14478 17554
rect 14530 17502 14868 17554
rect 14476 17500 14868 17502
rect 14476 17490 14532 17500
rect 14140 17444 14196 17454
rect 13468 16322 13636 16324
rect 13468 16270 13470 16322
rect 13522 16270 13636 16322
rect 13468 16268 13636 16270
rect 13916 17442 14196 17444
rect 13916 17390 14142 17442
rect 14194 17390 14196 17442
rect 13916 17388 14196 17390
rect 13468 16258 13524 16268
rect 13804 16212 13860 16222
rect 13804 16118 13860 16156
rect 13916 15426 13972 17388
rect 14140 17378 14196 17388
rect 14812 17220 14868 17500
rect 14924 17442 14980 17454
rect 14924 17390 14926 17442
rect 14978 17390 14980 17442
rect 14924 17332 14980 17390
rect 14924 17276 15204 17332
rect 14812 17164 15092 17220
rect 15036 17106 15092 17164
rect 15036 17054 15038 17106
rect 15090 17054 15092 17106
rect 15036 17042 15092 17054
rect 14700 16884 14756 16894
rect 14700 16770 14756 16828
rect 14700 16718 14702 16770
rect 14754 16718 14756 16770
rect 14700 16706 14756 16718
rect 15148 16660 15204 17276
rect 15596 16884 15652 21532
rect 15708 21522 15764 21532
rect 15932 21028 15988 21756
rect 16044 21810 16100 22652
rect 16380 22482 16436 22494
rect 16380 22430 16382 22482
rect 16434 22430 16436 22482
rect 16044 21758 16046 21810
rect 16098 21758 16100 21810
rect 16044 21746 16100 21758
rect 16156 22372 16212 22382
rect 16380 22372 16436 22430
rect 16716 22372 16772 22988
rect 16884 22988 16996 23044
rect 16828 22978 16884 22988
rect 16212 22316 16436 22372
rect 16604 22316 16772 22372
rect 16156 21810 16212 22316
rect 16156 21758 16158 21810
rect 16210 21758 16212 21810
rect 16156 21746 16212 21758
rect 16380 21812 16436 21822
rect 16380 21586 16436 21756
rect 16380 21534 16382 21586
rect 16434 21534 16436 21586
rect 16380 21522 16436 21534
rect 15596 16790 15652 16828
rect 15820 20972 16436 21028
rect 15372 16660 15428 16670
rect 15148 16658 15428 16660
rect 15148 16606 15374 16658
rect 15426 16606 15428 16658
rect 15148 16604 15428 16606
rect 14700 16548 14756 16558
rect 14028 16100 14084 16110
rect 14476 16100 14532 16110
rect 14028 16098 14308 16100
rect 14028 16046 14030 16098
rect 14082 16046 14308 16098
rect 14028 16044 14308 16046
rect 14028 16034 14084 16044
rect 13916 15374 13918 15426
rect 13970 15374 13972 15426
rect 13916 15362 13972 15374
rect 14252 15988 14308 16044
rect 14476 16006 14532 16044
rect 13244 15092 13412 15148
rect 13356 12402 13412 15092
rect 14140 14308 14196 14318
rect 13804 14306 14196 14308
rect 13804 14254 14142 14306
rect 14194 14254 14196 14306
rect 13804 14252 14196 14254
rect 13804 12962 13860 14252
rect 14140 14242 14196 14252
rect 13804 12910 13806 12962
rect 13858 12910 13860 12962
rect 13804 12898 13860 12910
rect 13356 12350 13358 12402
rect 13410 12350 13412 12402
rect 13356 12292 13412 12350
rect 13356 12226 13412 12236
rect 13468 12738 13524 12750
rect 13468 12686 13470 12738
rect 13522 12686 13524 12738
rect 12684 12178 12964 12180
rect 12684 12126 12686 12178
rect 12738 12126 12964 12178
rect 12684 12124 12964 12126
rect 12684 12114 12740 12124
rect 12908 11508 12964 12124
rect 13468 11844 13524 12686
rect 13804 12404 13860 12414
rect 13804 12310 13860 12348
rect 12908 11414 12964 11452
rect 13020 11788 13524 11844
rect 11844 10780 12068 10836
rect 11788 10742 11844 10780
rect 11564 10386 11620 10398
rect 11564 10334 11566 10386
rect 11618 10334 11620 10386
rect 11564 9940 11620 10334
rect 11564 9846 11620 9884
rect 12012 10050 12068 10780
rect 12124 10610 12180 11116
rect 12124 10558 12126 10610
rect 12178 10558 12180 10610
rect 12124 10546 12180 10558
rect 12348 11340 12516 11396
rect 12012 9998 12014 10050
rect 12066 9998 12068 10050
rect 12012 9938 12068 9998
rect 12012 9886 12014 9938
rect 12066 9886 12068 9938
rect 12012 9874 12068 9886
rect 11116 9774 11118 9826
rect 11170 9774 11172 9826
rect 11116 9762 11172 9774
rect 11340 9772 11508 9828
rect 10892 9602 10948 9614
rect 10892 9550 10894 9602
rect 10946 9550 10948 9602
rect 10780 9268 10836 9278
rect 10332 7074 10388 7084
rect 10668 7700 10724 7710
rect 10444 6916 10500 6926
rect 9660 5854 9662 5906
rect 9714 5854 9716 5906
rect 9660 5842 9716 5854
rect 10108 6076 10276 6132
rect 10332 6860 10444 6916
rect 10108 5796 10164 6076
rect 10332 6020 10388 6860
rect 10444 6850 10500 6860
rect 10444 6692 10500 6702
rect 10444 6598 10500 6636
rect 10668 6580 10724 7644
rect 10780 6916 10836 9212
rect 10780 6822 10836 6860
rect 10892 6804 10948 9550
rect 11116 7700 11172 7710
rect 11116 7474 11172 7644
rect 11116 7422 11118 7474
rect 11170 7422 11172 7474
rect 11116 7410 11172 7422
rect 11004 6804 11060 6814
rect 10948 6802 11060 6804
rect 10948 6750 11006 6802
rect 11058 6750 11060 6802
rect 10948 6748 11060 6750
rect 10892 6710 10948 6748
rect 11004 6738 11060 6748
rect 10668 6514 10724 6524
rect 10332 5964 10500 6020
rect 10332 5796 10388 5806
rect 10108 5794 10388 5796
rect 10108 5742 10334 5794
rect 10386 5742 10388 5794
rect 10108 5740 10388 5742
rect 10332 5730 10388 5740
rect 9324 5572 9380 5582
rect 9324 5234 9380 5516
rect 9324 5182 9326 5234
rect 9378 5182 9380 5234
rect 9324 5170 9380 5182
rect 10108 5236 10164 5246
rect 10444 5236 10500 5964
rect 10108 5234 10500 5236
rect 10108 5182 10110 5234
rect 10162 5182 10500 5234
rect 10108 5180 10500 5182
rect 10108 5170 10164 5180
rect 8988 4900 9044 4910
rect 8988 4898 9156 4900
rect 8988 4846 8990 4898
rect 9042 4846 9156 4898
rect 8988 4844 9156 4846
rect 8988 4834 9044 4844
rect 8988 4564 9044 4574
rect 8540 4562 9044 4564
rect 8540 4510 8990 4562
rect 9042 4510 9044 4562
rect 8540 4508 9044 4510
rect 8540 4338 8596 4508
rect 8988 4498 9044 4508
rect 8540 4286 8542 4338
rect 8594 4286 8596 4338
rect 8540 4274 8596 4286
rect 8316 3490 8372 3500
rect 8540 3554 8596 3566
rect 8540 3502 8542 3554
rect 8594 3502 8596 3554
rect 8540 3388 8596 3502
rect 6412 2830 6414 2882
rect 6466 2830 6468 2882
rect 6412 2818 6468 2830
rect 7084 3164 7588 3220
rect 7980 3332 8596 3388
rect 8764 3556 8820 3566
rect 6188 1822 6190 1874
rect 6242 1822 6244 1874
rect 6188 1810 6244 1822
rect 7084 1874 7140 3164
rect 7644 2658 7700 2670
rect 7644 2606 7646 2658
rect 7698 2606 7700 2658
rect 7644 1876 7700 2606
rect 7084 1822 7086 1874
rect 7138 1822 7140 1874
rect 7084 1810 7140 1822
rect 7420 1874 7700 1876
rect 7420 1822 7646 1874
rect 7698 1822 7700 1874
rect 7420 1820 7700 1822
rect 6748 1764 6804 1774
rect 6524 1708 6748 1764
rect 6524 400 6580 1708
rect 6748 1670 6804 1708
rect 7420 400 7476 1820
rect 7644 1810 7700 1820
rect 7980 1874 8036 3332
rect 8540 2658 8596 2670
rect 8540 2606 8542 2658
rect 8594 2606 8596 2658
rect 8540 1986 8596 2606
rect 8540 1934 8542 1986
rect 8594 1934 8596 1986
rect 8540 1876 8596 1934
rect 7980 1822 7982 1874
rect 8034 1822 8036 1874
rect 7980 1810 8036 1822
rect 8316 1820 8596 1876
rect 8764 1874 8820 3500
rect 9100 3444 9156 4844
rect 9772 4564 9828 4574
rect 9772 4470 9828 4508
rect 10780 4564 10836 4574
rect 10836 4508 10948 4564
rect 10780 4498 10836 4508
rect 10220 4450 10276 4462
rect 10220 4398 10222 4450
rect 10274 4398 10276 4450
rect 10108 4340 10164 4350
rect 10108 4246 10164 4284
rect 10108 3556 10164 3566
rect 9100 3378 9156 3388
rect 9884 3554 10164 3556
rect 9884 3502 10110 3554
rect 10162 3502 10164 3554
rect 9884 3500 10164 3502
rect 8764 1822 8766 1874
rect 8818 1822 8820 1874
rect 8316 400 8372 1820
rect 8764 1810 8820 1822
rect 9100 2658 9156 2670
rect 9100 2606 9102 2658
rect 9154 2606 9156 2658
rect 9100 1876 9156 2606
rect 9772 2660 9828 2670
rect 9772 2566 9828 2604
rect 9436 1876 9492 1886
rect 9100 1874 9492 1876
rect 9100 1822 9438 1874
rect 9490 1822 9492 1874
rect 9100 1820 9492 1822
rect 9212 400 9268 1820
rect 9436 1810 9492 1820
rect 9772 1876 9828 1886
rect 9884 1876 9940 3500
rect 10108 3490 10164 3500
rect 10220 3388 10276 4398
rect 10892 4450 10948 4508
rect 11340 4562 11396 9772
rect 11900 7364 11956 7374
rect 11900 7362 12292 7364
rect 11900 7310 11902 7362
rect 11954 7310 12292 7362
rect 11900 7308 12292 7310
rect 11900 7298 11956 7308
rect 11452 6916 11508 6926
rect 11452 6802 11508 6860
rect 12124 6916 12180 6926
rect 12124 6822 12180 6860
rect 11452 6750 11454 6802
rect 11506 6750 11508 6802
rect 11452 6738 11508 6750
rect 11788 6468 11844 6478
rect 11788 6466 12180 6468
rect 11788 6414 11790 6466
rect 11842 6414 12180 6466
rect 11788 6412 12180 6414
rect 11788 6402 11844 6412
rect 12124 5122 12180 6412
rect 12124 5070 12126 5122
rect 12178 5070 12180 5122
rect 12124 5058 12180 5070
rect 11900 4900 11956 4910
rect 12236 4900 12292 7308
rect 12348 6692 12404 11340
rect 12460 11172 12516 11182
rect 12460 11078 12516 11116
rect 12908 10724 12964 10734
rect 13020 10724 13076 11788
rect 14252 11508 14308 15932
rect 14588 15204 14644 15214
rect 14476 14530 14532 14542
rect 14476 14478 14478 14530
rect 14530 14478 14532 14530
rect 14476 14308 14532 14478
rect 14140 11452 14308 11508
rect 14364 12180 14420 12190
rect 12908 10722 13076 10724
rect 12908 10670 12910 10722
rect 12962 10670 13076 10722
rect 12908 10668 13076 10670
rect 13356 11172 13412 11182
rect 12908 10658 12964 10668
rect 13356 10052 13412 11116
rect 13356 9996 13524 10052
rect 13468 9826 13524 9996
rect 13468 9774 13470 9826
rect 13522 9774 13524 9826
rect 13468 7700 13524 9774
rect 13468 6692 13524 7644
rect 14028 7364 14084 7374
rect 14140 7364 14196 11452
rect 14252 11284 14308 11294
rect 14364 11284 14420 12124
rect 14476 11618 14532 14252
rect 14476 11566 14478 11618
rect 14530 11566 14532 11618
rect 14476 11554 14532 11566
rect 14252 11282 14420 11284
rect 14252 11230 14254 11282
rect 14306 11230 14420 11282
rect 14252 11228 14420 11230
rect 14252 11218 14308 11228
rect 14476 11172 14532 11182
rect 14364 11116 14476 11172
rect 14252 9940 14308 9950
rect 14364 9940 14420 11116
rect 14476 11106 14532 11116
rect 14252 9938 14420 9940
rect 14252 9886 14254 9938
rect 14306 9886 14420 9938
rect 14252 9884 14420 9886
rect 14252 9874 14308 9884
rect 14476 7700 14532 7710
rect 14476 7606 14532 7644
rect 14028 7362 14196 7364
rect 14028 7310 14030 7362
rect 14082 7310 14196 7362
rect 14028 7308 14196 7310
rect 14028 7298 14084 7308
rect 13692 6916 13748 6926
rect 13692 6802 13748 6860
rect 14364 6916 14420 6926
rect 14364 6822 14420 6860
rect 13692 6750 13694 6802
rect 13746 6750 13748 6802
rect 13692 6738 13748 6750
rect 14588 6802 14644 15148
rect 14700 14642 14756 16492
rect 15148 16100 15204 16604
rect 15372 16594 15428 16604
rect 15148 16034 15204 16044
rect 14924 15874 14980 15886
rect 14924 15822 14926 15874
rect 14978 15822 14980 15874
rect 14924 15316 14980 15822
rect 15820 15652 15876 20972
rect 16380 20914 16436 20972
rect 16380 20862 16382 20914
rect 16434 20862 16436 20914
rect 16380 20850 16436 20862
rect 16604 20692 16660 22316
rect 16828 22148 16884 22158
rect 16716 21812 16772 21822
rect 16716 20916 16772 21756
rect 16828 21810 16884 22092
rect 16828 21758 16830 21810
rect 16882 21758 16884 21810
rect 16828 21746 16884 21758
rect 16828 20916 16884 20926
rect 16716 20914 16884 20916
rect 16716 20862 16830 20914
rect 16882 20862 16884 20914
rect 16716 20860 16884 20862
rect 16044 20636 16660 20692
rect 15932 16212 15988 16222
rect 16044 16212 16100 20636
rect 16828 19460 16884 20860
rect 16716 19404 16884 19460
rect 16380 19348 16436 19358
rect 16156 19346 16436 19348
rect 16156 19294 16382 19346
rect 16434 19294 16436 19346
rect 16156 19292 16436 19294
rect 16156 16882 16212 19292
rect 16380 19282 16436 19292
rect 16268 17108 16324 17118
rect 16268 17014 16324 17052
rect 16716 16996 16772 19404
rect 16828 19236 16884 19246
rect 16828 19142 16884 19180
rect 16828 18452 16884 18462
rect 16940 18452 16996 22988
rect 17052 19236 17108 23492
rect 17276 19572 17332 26684
rect 17388 26516 17444 26526
rect 17388 26422 17444 26460
rect 17948 26290 18004 26852
rect 17948 26238 17950 26290
rect 18002 26238 18004 26290
rect 17948 26226 18004 26238
rect 17724 26068 17780 26078
rect 18060 26068 18116 30716
rect 18284 29428 18340 35308
rect 18396 34132 18452 34142
rect 18396 32786 18452 34076
rect 18396 32734 18398 32786
rect 18450 32734 18452 32786
rect 18396 32722 18452 32734
rect 17780 26012 18116 26068
rect 18172 29372 18340 29428
rect 18396 30212 18452 30222
rect 17724 25974 17780 26012
rect 18172 23492 18228 29372
rect 18396 29314 18452 30156
rect 18508 29764 18564 35420
rect 18620 35410 18676 35420
rect 18620 34914 18676 34926
rect 18844 34916 18900 42140
rect 18956 42130 19012 42140
rect 18956 38724 19012 38762
rect 18956 38658 19012 38668
rect 19068 38500 19124 42364
rect 19180 41972 19236 41982
rect 19180 41076 19236 41916
rect 19180 41010 19236 41020
rect 19180 40852 19236 40862
rect 19180 40402 19236 40796
rect 19180 40350 19182 40402
rect 19234 40350 19236 40402
rect 19180 39060 19236 40350
rect 19180 38994 19236 39004
rect 19180 38836 19236 38874
rect 19180 38770 19236 38780
rect 19292 38668 19348 43710
rect 19516 43538 19572 43550
rect 19516 43486 19518 43538
rect 19570 43486 19572 43538
rect 19516 42196 19572 43486
rect 19516 42130 19572 42140
rect 19516 41972 19572 41982
rect 19516 41878 19572 41916
rect 19516 41076 19572 41086
rect 19516 39842 19572 41020
rect 19516 39790 19518 39842
rect 19570 39790 19572 39842
rect 19516 39778 19572 39790
rect 18956 38444 19124 38500
rect 19180 38612 19348 38668
rect 19516 39508 19572 39518
rect 19516 38836 19572 39452
rect 19516 38722 19572 38780
rect 19516 38670 19518 38722
rect 19570 38670 19572 38722
rect 19516 38658 19572 38670
rect 18956 35028 19012 38444
rect 19180 35308 19236 38612
rect 19404 38500 19460 38510
rect 19292 35588 19348 35598
rect 19292 35474 19348 35532
rect 19292 35422 19294 35474
rect 19346 35422 19348 35474
rect 19292 35410 19348 35422
rect 19180 35252 19348 35308
rect 18956 34962 19012 34972
rect 18620 34862 18622 34914
rect 18674 34862 18676 34914
rect 18620 34580 18676 34862
rect 18620 34514 18676 34524
rect 18732 34860 18900 34916
rect 18620 34242 18676 34254
rect 18620 34190 18622 34242
rect 18674 34190 18676 34242
rect 18620 33458 18676 34190
rect 18620 33406 18622 33458
rect 18674 33406 18676 33458
rect 18620 33394 18676 33406
rect 18732 30100 18788 34860
rect 18844 34692 18900 34702
rect 18844 34598 18900 34636
rect 19180 34690 19236 34702
rect 19180 34638 19182 34690
rect 19234 34638 19236 34690
rect 19180 34580 19236 34638
rect 18956 34356 19012 34366
rect 18844 34132 18900 34142
rect 18844 34038 18900 34076
rect 18844 30324 18900 30334
rect 18844 30230 18900 30268
rect 18732 30044 18900 30100
rect 18508 29698 18564 29708
rect 18396 29262 18398 29314
rect 18450 29262 18452 29314
rect 18396 28756 18452 29262
rect 18396 28690 18452 28700
rect 18732 29652 18788 29662
rect 18620 28644 18676 28654
rect 18508 28084 18564 28094
rect 18396 28028 18508 28084
rect 18284 23826 18340 23838
rect 18284 23774 18286 23826
rect 18338 23774 18340 23826
rect 18284 23604 18340 23774
rect 18284 23538 18340 23548
rect 18172 23426 18228 23436
rect 17388 23268 17444 23278
rect 17388 22372 17444 23212
rect 17948 23268 18004 23278
rect 17948 23154 18004 23212
rect 17948 23102 17950 23154
rect 18002 23102 18004 23154
rect 17948 23090 18004 23102
rect 17612 23044 17668 23054
rect 17612 22950 17668 22988
rect 18172 23044 18228 23054
rect 18172 22950 18228 22988
rect 17388 21586 17444 22316
rect 18396 21700 18452 28028
rect 18508 27990 18564 28028
rect 18620 27860 18676 28588
rect 18508 23938 18564 23950
rect 18508 23886 18510 23938
rect 18562 23886 18564 23938
rect 18508 23380 18564 23886
rect 18508 23314 18564 23324
rect 18508 22930 18564 22942
rect 18508 22878 18510 22930
rect 18562 22878 18564 22930
rect 18508 22596 18564 22878
rect 18508 22530 18564 22540
rect 18508 22260 18564 22270
rect 18508 22166 18564 22204
rect 17388 21534 17390 21586
rect 17442 21534 17444 21586
rect 17388 21476 17444 21534
rect 17388 21410 17444 21420
rect 17500 21644 18452 21700
rect 17052 19170 17108 19180
rect 17164 19516 17332 19572
rect 17388 20804 17444 20814
rect 17164 19234 17220 19516
rect 17276 19348 17332 19358
rect 17276 19254 17332 19292
rect 17164 19182 17166 19234
rect 17218 19182 17220 19234
rect 17164 19170 17220 19182
rect 17276 19124 17332 19134
rect 16828 18450 16996 18452
rect 16828 18398 16830 18450
rect 16882 18398 16996 18450
rect 16828 18396 16996 18398
rect 16828 18386 16884 18396
rect 16940 18228 16996 18396
rect 16940 18162 16996 18172
rect 17164 19010 17220 19022
rect 17164 18958 17166 19010
rect 17218 18958 17220 19010
rect 16940 18004 16996 18014
rect 16156 16830 16158 16882
rect 16210 16830 16212 16882
rect 16156 16548 16212 16830
rect 16492 16882 16548 16894
rect 16492 16830 16494 16882
rect 16546 16830 16548 16882
rect 16380 16772 16436 16782
rect 16380 16678 16436 16716
rect 16156 16482 16212 16492
rect 15932 16210 16100 16212
rect 15932 16158 15934 16210
rect 15986 16158 16100 16210
rect 15932 16156 16100 16158
rect 15932 16146 15988 16156
rect 16492 15764 16548 16830
rect 16716 16882 16772 16940
rect 16716 16830 16718 16882
rect 16770 16830 16772 16882
rect 16716 16818 16772 16830
rect 16828 17948 16940 18004
rect 15820 15586 15876 15596
rect 16044 15708 16548 15764
rect 14924 15250 14980 15260
rect 16044 15204 16100 15708
rect 16044 15138 16100 15148
rect 16492 15540 16548 15550
rect 16492 15316 16548 15484
rect 14700 14590 14702 14642
rect 14754 14590 14756 14642
rect 14700 14578 14756 14590
rect 15148 14308 15204 14318
rect 15148 13636 15204 14252
rect 15148 13524 15204 13580
rect 15036 13468 15204 13524
rect 15036 12402 15092 13468
rect 16156 13076 16212 13086
rect 15036 12350 15038 12402
rect 15090 12350 15092 12402
rect 15036 12338 15092 12350
rect 15484 12404 15540 12414
rect 15932 12404 15988 12414
rect 15484 12310 15540 12348
rect 15820 12348 15932 12404
rect 14812 12180 14868 12190
rect 14700 12124 14812 12180
rect 14700 11284 14756 12124
rect 14812 12114 14868 12124
rect 14812 11508 14868 11518
rect 14812 11506 15428 11508
rect 14812 11454 14814 11506
rect 14866 11454 15428 11506
rect 14812 11452 15428 11454
rect 14812 11442 14868 11452
rect 15372 11394 15428 11452
rect 15372 11342 15374 11394
rect 15426 11342 15428 11394
rect 15372 11330 15428 11342
rect 15820 11394 15876 12348
rect 15932 12338 15988 12348
rect 16156 12402 16212 13020
rect 16156 12350 16158 12402
rect 16210 12350 16212 12402
rect 16156 12338 16212 12350
rect 16492 12404 16548 15260
rect 16492 12338 16548 12348
rect 16604 12516 16660 12526
rect 15932 12180 15988 12190
rect 15932 12086 15988 12124
rect 16268 12180 16324 12190
rect 16268 12086 16324 12124
rect 16380 12178 16436 12190
rect 16380 12126 16382 12178
rect 16434 12126 16436 12178
rect 15820 11342 15822 11394
rect 15874 11342 15876 11394
rect 15708 11284 15764 11294
rect 14700 11228 15092 11284
rect 15036 10498 15092 11228
rect 15148 11172 15204 11182
rect 15148 11078 15204 11116
rect 15036 10446 15038 10498
rect 15090 10446 15092 10498
rect 15036 10434 15092 10446
rect 15708 9266 15764 11228
rect 15820 10836 15876 11342
rect 15820 10770 15876 10780
rect 16156 10836 16212 10846
rect 16156 10742 16212 10780
rect 15820 10610 15876 10622
rect 15820 10558 15822 10610
rect 15874 10558 15876 10610
rect 15820 10500 15876 10558
rect 15820 10434 15876 10444
rect 16380 10164 16436 12126
rect 16604 12178 16660 12460
rect 16604 12126 16606 12178
rect 16658 12126 16660 12178
rect 16604 12114 16660 12126
rect 16604 11284 16660 11294
rect 16604 11190 16660 11228
rect 16604 10836 16660 10846
rect 16660 10780 16772 10836
rect 16604 10770 16660 10780
rect 16380 10108 16548 10164
rect 16380 9940 16436 9950
rect 16380 9846 16436 9884
rect 15708 9214 15710 9266
rect 15762 9214 15764 9266
rect 15708 9202 15764 9214
rect 15484 9042 15540 9054
rect 15484 8990 15486 9042
rect 15538 8990 15540 9042
rect 15484 8932 15540 8990
rect 16268 8932 16324 8942
rect 15484 8930 16324 8932
rect 15484 8878 16270 8930
rect 16322 8878 16324 8930
rect 15484 8876 16324 8878
rect 16268 8866 16324 8876
rect 15932 8036 15988 8046
rect 15932 7924 15988 7980
rect 15708 7868 15988 7924
rect 15708 7252 15764 7868
rect 16492 7700 16548 10108
rect 16716 9940 16772 10780
rect 16828 10500 16884 17948
rect 16940 17938 16996 17948
rect 16940 17108 16996 17118
rect 16940 13076 16996 17052
rect 17052 13076 17108 13086
rect 16940 13020 17052 13076
rect 17052 12982 17108 13020
rect 17164 12404 17220 18958
rect 17276 15538 17332 19068
rect 17388 18004 17444 20748
rect 17388 17938 17444 17948
rect 17500 17108 17556 21644
rect 17724 21476 17780 21486
rect 17724 20914 17780 21420
rect 17724 20862 17726 20914
rect 17778 20862 17780 20914
rect 17724 20850 17780 20862
rect 18172 21474 18228 21486
rect 18172 21422 18174 21474
rect 18226 21422 18228 21474
rect 18172 20242 18228 21422
rect 18620 21028 18676 27804
rect 18284 20972 18676 21028
rect 18732 21028 18788 29596
rect 18844 23940 18900 30044
rect 18844 23874 18900 23884
rect 18844 23716 18900 23726
rect 18844 23622 18900 23660
rect 18732 20972 18900 21028
rect 18284 20914 18340 20972
rect 18284 20862 18286 20914
rect 18338 20862 18340 20914
rect 18284 20804 18340 20862
rect 18284 20738 18340 20748
rect 18172 20190 18174 20242
rect 18226 20190 18228 20242
rect 18172 20178 18228 20190
rect 17836 20020 17892 20030
rect 17724 20018 17892 20020
rect 17724 19966 17838 20018
rect 17890 19966 17892 20018
rect 17724 19964 17892 19966
rect 17724 18674 17780 19964
rect 17836 19954 17892 19964
rect 17724 18622 17726 18674
rect 17778 18622 17780 18674
rect 17724 18610 17780 18622
rect 18284 18338 18340 18350
rect 18284 18286 18286 18338
rect 18338 18286 18340 18338
rect 18060 18228 18116 18238
rect 18060 18134 18116 18172
rect 17500 17014 17556 17052
rect 17836 17778 17892 17790
rect 17836 17726 17838 17778
rect 17890 17726 17892 17778
rect 17612 16996 17668 17006
rect 17276 15486 17278 15538
rect 17330 15486 17332 15538
rect 17276 15474 17332 15486
rect 17388 16772 17444 16782
rect 17388 15316 17444 16716
rect 17500 15316 17556 15326
rect 17388 15314 17556 15316
rect 17388 15262 17502 15314
rect 17554 15262 17556 15314
rect 17388 15260 17556 15262
rect 17500 15250 17556 15260
rect 17612 15148 17668 16940
rect 17836 16324 17892 17726
rect 17948 16996 18004 17006
rect 17948 16902 18004 16940
rect 18284 16548 18340 18286
rect 18284 16482 18340 16492
rect 18732 16772 18788 16782
rect 17836 16258 17892 16268
rect 18732 16098 18788 16716
rect 18732 16046 18734 16098
rect 18786 16046 18788 16098
rect 18060 15988 18116 15998
rect 17388 15092 17668 15148
rect 17724 15986 18116 15988
rect 17724 15934 18062 15986
rect 18114 15934 18116 15986
rect 17724 15932 18116 15934
rect 17388 13076 17444 15092
rect 17500 14532 17556 14542
rect 17500 14530 17668 14532
rect 17500 14478 17502 14530
rect 17554 14478 17668 14530
rect 17500 14476 17668 14478
rect 17500 14466 17556 14476
rect 17612 13970 17668 14476
rect 17724 14418 17780 15932
rect 18060 15922 18116 15932
rect 18732 15540 18788 16046
rect 18732 15474 18788 15484
rect 17836 15428 17892 15438
rect 17836 15334 17892 15372
rect 18172 15426 18228 15438
rect 18172 15374 18174 15426
rect 18226 15374 18228 15426
rect 18172 15316 18228 15374
rect 18172 15250 18228 15260
rect 18284 15204 18340 15242
rect 18844 15148 18900 20972
rect 18956 18452 19012 34300
rect 19180 32228 19236 34524
rect 19292 34356 19348 35252
rect 19292 34290 19348 34300
rect 19180 32162 19236 32172
rect 19292 34130 19348 34142
rect 19292 34078 19294 34130
rect 19346 34078 19348 34130
rect 19068 30882 19124 30894
rect 19068 30830 19070 30882
rect 19122 30830 19124 30882
rect 19068 29876 19124 30830
rect 19180 30324 19236 30334
rect 19292 30324 19348 34078
rect 19404 30660 19460 38444
rect 19516 37492 19572 37502
rect 19516 37398 19572 37436
rect 19628 36484 19684 51660
rect 20188 51604 20244 52110
rect 20300 52052 20356 53228
rect 20524 53060 20580 58492
rect 20748 58482 20804 58492
rect 20636 57652 20692 57662
rect 20636 55410 20692 57596
rect 20636 55358 20638 55410
rect 20690 55358 20692 55410
rect 20636 53732 20692 55358
rect 20860 55412 20916 55422
rect 20748 54402 20804 54414
rect 20748 54350 20750 54402
rect 20802 54350 20804 54402
rect 20748 53956 20804 54350
rect 20748 53890 20804 53900
rect 20692 53676 20804 53732
rect 20636 53666 20692 53676
rect 20300 51958 20356 51996
rect 20412 52722 20468 52734
rect 20412 52670 20414 52722
rect 20466 52670 20468 52722
rect 19964 51548 20244 51604
rect 19964 51378 20020 51548
rect 19964 51326 19966 51378
rect 20018 51326 20020 51378
rect 19964 51314 20020 51326
rect 20412 51378 20468 52670
rect 20524 52050 20580 53004
rect 20636 53506 20692 53518
rect 20636 53454 20638 53506
rect 20690 53454 20692 53506
rect 20636 52948 20692 53454
rect 20636 52854 20692 52892
rect 20748 52836 20804 53676
rect 20860 53506 20916 55356
rect 20860 53454 20862 53506
rect 20914 53454 20916 53506
rect 20860 53442 20916 53454
rect 20748 52770 20804 52780
rect 20860 52164 20916 52174
rect 20860 52070 20916 52108
rect 20524 51998 20526 52050
rect 20578 51998 20580 52050
rect 20524 51986 20580 51998
rect 20412 51326 20414 51378
rect 20466 51326 20468 51378
rect 20412 51314 20468 51326
rect 20524 51492 20580 51502
rect 20076 50484 20132 50494
rect 20076 50372 20468 50428
rect 19836 50204 20100 50214
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 19836 50138 20100 50148
rect 20412 50148 20468 50372
rect 20412 50082 20468 50092
rect 20524 50034 20580 51436
rect 20636 51380 20692 51390
rect 20860 51380 20916 51390
rect 20636 51378 20916 51380
rect 20636 51326 20638 51378
rect 20690 51326 20862 51378
rect 20914 51326 20916 51378
rect 20636 51324 20916 51326
rect 20636 51314 20692 51324
rect 20860 51314 20916 51324
rect 20524 49982 20526 50034
rect 20578 49982 20580 50034
rect 20524 49970 20580 49982
rect 20636 50596 20692 50606
rect 20300 49924 20356 49934
rect 20300 49922 20468 49924
rect 20300 49870 20302 49922
rect 20354 49870 20468 49922
rect 20300 49868 20468 49870
rect 20300 49858 20356 49868
rect 20188 49812 20244 49822
rect 20188 49718 20244 49756
rect 19852 49698 19908 49710
rect 19852 49646 19854 49698
rect 19906 49646 19908 49698
rect 19852 49586 19908 49646
rect 19852 49534 19854 49586
rect 19906 49534 19908 49586
rect 19852 49522 19908 49534
rect 20188 48914 20244 48926
rect 20188 48862 20190 48914
rect 20242 48862 20244 48914
rect 19836 48636 20100 48646
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 19836 48570 20100 48580
rect 20188 48468 20244 48862
rect 20076 48412 20244 48468
rect 20076 47460 20132 48412
rect 20076 47404 20244 47460
rect 20076 47236 20132 47274
rect 20076 47170 20132 47180
rect 19836 47068 20100 47078
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 19836 47002 20100 47012
rect 19964 46788 20020 46798
rect 20188 46788 20244 47404
rect 20020 46732 20244 46788
rect 19964 46694 20020 46732
rect 19852 45780 19908 45790
rect 19852 45686 19908 45724
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 20300 44436 20356 44446
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 19852 43538 19908 43550
rect 19852 43486 19854 43538
rect 19906 43486 19908 43538
rect 19852 43428 19908 43486
rect 19852 43362 19908 43372
rect 20300 43204 20356 44380
rect 20412 43876 20468 49868
rect 20524 49588 20580 49598
rect 20524 48244 20580 49532
rect 20636 48804 20692 50540
rect 20748 50596 20804 50606
rect 20748 50594 20916 50596
rect 20748 50542 20750 50594
rect 20802 50542 20916 50594
rect 20748 50540 20916 50542
rect 20748 50530 20804 50540
rect 20860 50036 20916 50540
rect 20860 49970 20916 49980
rect 20748 49924 20804 49934
rect 20748 49028 20804 49868
rect 20748 49026 20916 49028
rect 20748 48974 20750 49026
rect 20802 48974 20916 49026
rect 20748 48972 20916 48974
rect 20748 48962 20804 48972
rect 20636 48748 20804 48804
rect 20524 47068 20580 48188
rect 20748 47234 20804 48748
rect 20748 47182 20750 47234
rect 20802 47182 20804 47234
rect 20524 47012 20692 47068
rect 20524 45892 20580 45902
rect 20524 45798 20580 45836
rect 20412 43810 20468 43820
rect 20524 45106 20580 45118
rect 20524 45054 20526 45106
rect 20578 45054 20580 45106
rect 20188 43148 20356 43204
rect 20412 43652 20468 43662
rect 20524 43652 20580 45054
rect 20412 43650 20580 43652
rect 20412 43598 20414 43650
rect 20466 43598 20580 43650
rect 20412 43596 20580 43598
rect 20636 44436 20692 47012
rect 20748 44884 20804 47182
rect 20860 47124 20916 48972
rect 20860 46564 20916 47068
rect 20860 46498 20916 46508
rect 20748 44818 20804 44828
rect 20748 44436 20804 44446
rect 20636 44434 20804 44436
rect 20636 44382 20750 44434
rect 20802 44382 20804 44434
rect 20636 44380 20804 44382
rect 20412 43204 20468 43596
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 20076 42084 20132 42094
rect 20076 41074 20132 42028
rect 20076 41022 20078 41074
rect 20130 41022 20132 41074
rect 20076 40964 20132 41022
rect 20076 40898 20132 40908
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 19964 39842 20020 39854
rect 19964 39790 19966 39842
rect 20018 39790 20020 39842
rect 19964 39730 20020 39790
rect 19964 39678 19966 39730
rect 20018 39678 20020 39730
rect 19964 39666 20020 39678
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 19964 37154 20020 37166
rect 19964 37102 19966 37154
rect 20018 37102 20020 37154
rect 19964 37044 20020 37102
rect 19964 36978 20020 36988
rect 19628 36418 19684 36428
rect 19628 36260 19684 36270
rect 19628 35812 19684 36204
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19964 35924 20020 35934
rect 19740 35812 19796 35822
rect 19628 35810 19796 35812
rect 19628 35758 19742 35810
rect 19794 35758 19796 35810
rect 19628 35756 19796 35758
rect 19740 35746 19796 35756
rect 19964 35810 20020 35868
rect 19964 35758 19966 35810
rect 20018 35758 20020 35810
rect 19964 35746 20020 35758
rect 19516 35698 19572 35710
rect 19516 35646 19518 35698
rect 19570 35646 19572 35698
rect 19516 34356 19572 35646
rect 20076 35698 20132 35710
rect 20076 35646 20078 35698
rect 20130 35646 20132 35698
rect 20076 35588 20132 35646
rect 20076 35522 20132 35532
rect 19628 35364 19684 35374
rect 19628 35026 19684 35308
rect 19628 34974 19630 35026
rect 19682 34974 19684 35026
rect 19628 34804 19684 34974
rect 19628 34738 19684 34748
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19628 34356 19684 34366
rect 19516 34354 19684 34356
rect 19516 34302 19630 34354
rect 19682 34302 19684 34354
rect 19516 34300 19684 34302
rect 19628 34290 19684 34300
rect 19516 34130 19572 34142
rect 19516 34078 19518 34130
rect 19570 34078 19572 34130
rect 19516 33908 19572 34078
rect 19516 31108 19572 33852
rect 19740 34130 19796 34142
rect 19740 34078 19742 34130
rect 19794 34078 19796 34130
rect 19740 33572 19796 34078
rect 19852 34130 19908 34142
rect 19852 34078 19854 34130
rect 19906 34078 19908 34130
rect 19852 34020 19908 34078
rect 19852 33954 19908 33964
rect 19740 33506 19796 33516
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19628 32228 19684 32238
rect 19628 31220 19684 32172
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19628 31164 19796 31220
rect 19516 31042 19572 31052
rect 19516 30884 19572 30894
rect 19516 30882 19684 30884
rect 19516 30830 19518 30882
rect 19570 30830 19684 30882
rect 19516 30828 19684 30830
rect 19516 30818 19572 30828
rect 19404 30604 19572 30660
rect 19404 30436 19460 30446
rect 19404 30342 19460 30380
rect 19236 30268 19348 30324
rect 19180 30230 19236 30268
rect 19516 30212 19572 30604
rect 19628 30436 19684 30828
rect 19628 30370 19684 30380
rect 19740 30212 19796 31164
rect 19964 31108 20020 31118
rect 19964 31106 20132 31108
rect 19964 31054 19966 31106
rect 20018 31054 20132 31106
rect 19964 31052 20132 31054
rect 19964 31042 20020 31052
rect 19852 30996 19908 31006
rect 19852 30902 19908 30940
rect 19964 30884 20020 30894
rect 19964 30770 20020 30828
rect 19964 30718 19966 30770
rect 20018 30718 20020 30770
rect 19964 30706 20020 30718
rect 20076 30548 20132 31052
rect 19068 29428 19124 29820
rect 19068 28868 19124 29372
rect 19404 30156 19572 30212
rect 19628 30156 19796 30212
rect 19964 30492 20132 30548
rect 19964 30212 20020 30492
rect 19180 28868 19236 28878
rect 19068 28866 19236 28868
rect 19068 28814 19182 28866
rect 19234 28814 19236 28866
rect 19068 28812 19236 28814
rect 19180 28802 19236 28812
rect 19068 25396 19124 25406
rect 19068 23380 19124 25340
rect 19404 24164 19460 30156
rect 19628 26908 19684 30156
rect 19964 30146 20020 30156
rect 20076 30098 20132 30110
rect 20076 30046 20078 30098
rect 20130 30046 20132 30098
rect 19740 29988 19796 29998
rect 20076 29988 20132 30046
rect 19740 29986 20132 29988
rect 19740 29934 19742 29986
rect 19794 29934 20132 29986
rect 19740 29932 20132 29934
rect 19740 29922 19796 29932
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 20188 29764 20244 43148
rect 20412 43138 20468 43148
rect 20636 42980 20692 44380
rect 20748 44370 20804 44380
rect 20300 42924 20692 42980
rect 20300 42754 20356 42924
rect 20748 42868 20804 42878
rect 20748 42774 20804 42812
rect 20300 42702 20302 42754
rect 20354 42702 20356 42754
rect 20300 41972 20356 42702
rect 20636 42420 20692 42430
rect 20636 42084 20692 42364
rect 20300 39730 20356 41916
rect 20524 42082 20692 42084
rect 20524 42030 20638 42082
rect 20690 42030 20692 42082
rect 20524 42028 20692 42030
rect 20412 40516 20468 40526
rect 20524 40516 20580 42028
rect 20636 42018 20692 42028
rect 20748 41972 20804 41982
rect 20468 40460 20580 40516
rect 20636 41636 20692 41646
rect 20412 40422 20468 40460
rect 20300 39678 20302 39730
rect 20354 39678 20356 39730
rect 20300 38724 20356 39678
rect 20636 39732 20692 41580
rect 20748 41186 20804 41916
rect 20748 41134 20750 41186
rect 20802 41134 20804 41186
rect 20748 41122 20804 41134
rect 20860 40964 20916 40974
rect 20860 40514 20916 40908
rect 20860 40462 20862 40514
rect 20914 40462 20916 40514
rect 20860 40450 20916 40462
rect 20860 39732 20916 39742
rect 20636 39730 20916 39732
rect 20636 39678 20862 39730
rect 20914 39678 20916 39730
rect 20636 39676 20916 39678
rect 20860 39666 20916 39676
rect 20300 38658 20356 38668
rect 20412 39060 20468 39070
rect 20300 37268 20356 37278
rect 20300 29988 20356 37212
rect 20412 37156 20468 39004
rect 20524 38162 20580 38174
rect 20524 38110 20526 38162
rect 20578 38110 20580 38162
rect 20524 37940 20580 38110
rect 20524 37874 20580 37884
rect 20748 38052 20804 38062
rect 20748 37490 20804 37996
rect 20748 37438 20750 37490
rect 20802 37438 20804 37490
rect 20748 37426 20804 37438
rect 20524 37156 20580 37166
rect 20412 37154 20692 37156
rect 20412 37102 20526 37154
rect 20578 37102 20692 37154
rect 20412 37100 20692 37102
rect 20524 37090 20580 37100
rect 20524 36708 20580 36718
rect 20524 35922 20580 36652
rect 20524 35870 20526 35922
rect 20578 35870 20580 35922
rect 20524 35858 20580 35870
rect 20300 29922 20356 29932
rect 20412 29988 20468 29998
rect 20412 29986 20580 29988
rect 20412 29934 20414 29986
rect 20466 29934 20580 29986
rect 20412 29932 20580 29934
rect 20412 29922 20468 29932
rect 20188 29708 20468 29764
rect 20300 29540 20356 29550
rect 20300 28866 20356 29484
rect 20300 28814 20302 28866
rect 20354 28814 20356 28866
rect 20300 28802 20356 28814
rect 20188 28532 20244 28542
rect 20188 28438 20244 28476
rect 20300 28418 20356 28430
rect 20300 28366 20302 28418
rect 20354 28366 20356 28418
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 20300 28084 20356 28366
rect 19852 28028 20356 28084
rect 19852 27186 19908 28028
rect 20076 27860 20132 27870
rect 20076 27766 20132 27804
rect 19852 27134 19854 27186
rect 19906 27134 19908 27186
rect 19852 27122 19908 27134
rect 20300 27076 20356 27086
rect 20300 26982 20356 27020
rect 19068 23286 19124 23324
rect 19292 24108 19460 24164
rect 19516 26852 19684 26908
rect 19180 22372 19236 22382
rect 19180 22278 19236 22316
rect 19292 21028 19348 24108
rect 19516 24052 19572 26852
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19628 25284 19684 25294
rect 19628 24162 19684 25228
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 19628 24110 19630 24162
rect 19682 24110 19684 24162
rect 19628 24098 19684 24110
rect 20412 24052 20468 29708
rect 20524 29538 20580 29932
rect 20524 29486 20526 29538
rect 20578 29486 20580 29538
rect 20524 29474 20580 29486
rect 20524 28532 20580 28542
rect 20524 28082 20580 28476
rect 20524 28030 20526 28082
rect 20578 28030 20580 28082
rect 20524 28018 20580 28030
rect 20636 26908 20692 37100
rect 20860 35924 20916 35934
rect 20972 35924 21028 59054
rect 21308 59108 21364 59724
rect 21532 59444 21588 59454
rect 21532 59330 21588 59388
rect 21532 59278 21534 59330
rect 21586 59278 21588 59330
rect 21532 59266 21588 59278
rect 21308 59052 21588 59108
rect 21420 58436 21476 58446
rect 21420 58342 21476 58380
rect 21420 55076 21476 55086
rect 21420 54982 21476 55020
rect 21420 54626 21476 54638
rect 21420 54574 21422 54626
rect 21474 54574 21476 54626
rect 21196 54516 21252 54526
rect 21196 54514 21364 54516
rect 21196 54462 21198 54514
rect 21250 54462 21364 54514
rect 21196 54460 21364 54462
rect 21196 54450 21252 54460
rect 21308 53954 21364 54460
rect 21308 53902 21310 53954
rect 21362 53902 21364 53954
rect 21308 53890 21364 53902
rect 21308 52948 21364 52958
rect 21196 52892 21308 52948
rect 21084 52164 21140 52174
rect 21084 49700 21140 52108
rect 21084 49634 21140 49644
rect 21084 48354 21140 48366
rect 21084 48302 21086 48354
rect 21138 48302 21140 48354
rect 21084 46788 21140 48302
rect 21084 45780 21140 46732
rect 21084 45714 21140 45724
rect 21196 48242 21252 52892
rect 21308 52854 21364 52892
rect 21420 52276 21476 54574
rect 21532 54516 21588 59052
rect 21756 58772 21812 60060
rect 21868 60004 21924 60396
rect 21980 60004 22036 60014
rect 21868 60002 22036 60004
rect 21868 59950 21982 60002
rect 22034 59950 22036 60002
rect 21868 59948 22036 59950
rect 21980 59938 22036 59948
rect 21756 58716 22148 58772
rect 22092 58546 22148 58716
rect 22092 58494 22094 58546
rect 22146 58494 22148 58546
rect 22092 58482 22148 58494
rect 21868 57650 21924 57662
rect 21868 57598 21870 57650
rect 21922 57598 21924 57650
rect 21868 57540 21924 57598
rect 21868 55076 21924 57484
rect 22092 57092 22148 57102
rect 22092 56978 22148 57036
rect 22092 56926 22094 56978
rect 22146 56926 22148 56978
rect 22092 56914 22148 56926
rect 22092 55412 22148 55422
rect 22092 55188 22148 55356
rect 22092 55122 22148 55132
rect 21868 55010 21924 55020
rect 22204 54852 22260 62972
rect 22876 62468 22932 63084
rect 22988 62580 23044 63870
rect 23100 63700 23156 65660
rect 23212 65492 23268 65502
rect 23436 65492 23492 66894
rect 23212 65398 23268 65436
rect 23324 65490 23492 65492
rect 23324 65438 23438 65490
rect 23490 65438 23492 65490
rect 23324 65436 23492 65438
rect 23324 64932 23380 65436
rect 23436 65426 23492 65436
rect 23772 66946 23940 66948
rect 23772 66894 23886 66946
rect 23938 66894 23940 66946
rect 23772 66892 23940 66894
rect 23772 65268 23828 66892
rect 23884 66882 23940 66892
rect 23996 66834 24052 66846
rect 23996 66782 23998 66834
rect 24050 66782 24052 66834
rect 23996 66724 24052 66782
rect 23212 64876 23380 64932
rect 23436 65212 23828 65268
rect 23884 66668 24052 66724
rect 23884 65490 23940 66668
rect 23884 65438 23886 65490
rect 23938 65438 23940 65490
rect 23212 64372 23268 64876
rect 23212 64146 23268 64316
rect 23212 64094 23214 64146
rect 23266 64094 23268 64146
rect 23212 63812 23268 64094
rect 23324 64708 23380 64718
rect 23436 64708 23492 65212
rect 23324 64706 23492 64708
rect 23324 64654 23326 64706
rect 23378 64654 23492 64706
rect 23324 64652 23492 64654
rect 23548 64708 23604 64718
rect 23548 64706 23716 64708
rect 23548 64654 23550 64706
rect 23602 64654 23716 64706
rect 23548 64652 23716 64654
rect 23324 64036 23380 64652
rect 23548 64642 23604 64652
rect 23324 63970 23380 63980
rect 23548 63924 23604 63934
rect 23548 63830 23604 63868
rect 23660 63812 23716 64652
rect 23884 64596 23940 65438
rect 23996 65492 24052 65502
rect 23996 65398 24052 65436
rect 24108 65268 24164 67902
rect 24332 66946 24388 66958
rect 24332 66894 24334 66946
rect 24386 66894 24388 66946
rect 24332 66834 24388 66894
rect 24332 66782 24334 66834
rect 24386 66782 24388 66834
rect 24332 66770 24388 66782
rect 24220 65380 24276 65390
rect 24220 65286 24276 65324
rect 24108 65202 24164 65212
rect 24108 64708 24164 64718
rect 24108 64614 24164 64652
rect 24332 64706 24388 64718
rect 24332 64654 24334 64706
rect 24386 64654 24388 64706
rect 23884 64530 23940 64540
rect 23772 64372 23828 64382
rect 23772 63922 23828 64316
rect 24332 64372 24388 64654
rect 24332 64306 24388 64316
rect 23772 63870 23774 63922
rect 23826 63870 23828 63922
rect 23772 63858 23828 63870
rect 23884 63924 23940 63934
rect 23212 63756 23492 63812
rect 23100 63644 23268 63700
rect 23100 63138 23156 63150
rect 23100 63086 23102 63138
rect 23154 63086 23156 63138
rect 23100 63028 23156 63086
rect 23100 62962 23156 62972
rect 23100 62580 23156 62590
rect 22988 62524 23100 62580
rect 23100 62486 23156 62524
rect 22876 62412 23044 62468
rect 22988 62354 23044 62412
rect 22988 62302 22990 62354
rect 23042 62302 23044 62354
rect 22316 62244 22372 62254
rect 22316 57874 22372 62188
rect 22652 61348 22708 61358
rect 22540 61012 22596 61022
rect 22316 57822 22318 57874
rect 22370 57822 22372 57874
rect 22316 57652 22372 57822
rect 22316 57586 22372 57596
rect 22428 60676 22484 60686
rect 22428 60114 22484 60620
rect 22428 60062 22430 60114
rect 22482 60062 22484 60114
rect 21868 54796 22260 54852
rect 21868 54738 21924 54796
rect 21868 54686 21870 54738
rect 21922 54686 21924 54738
rect 21868 54674 21924 54686
rect 21532 54450 21588 54460
rect 21644 53956 21700 53966
rect 21644 53862 21700 53900
rect 21868 53620 21924 53630
rect 21532 53060 21588 53070
rect 21868 53060 21924 53564
rect 21980 53508 22036 54796
rect 22428 54628 22484 60062
rect 22540 55412 22596 60956
rect 22652 58828 22708 61292
rect 22988 61348 23044 62302
rect 23212 62244 23268 63644
rect 22988 61282 23044 61292
rect 23100 62020 23156 62030
rect 23100 61458 23156 61964
rect 23100 61406 23102 61458
rect 23154 61406 23156 61458
rect 23100 61012 23156 61406
rect 23100 60946 23156 60956
rect 23212 61010 23268 62188
rect 23212 60958 23214 61010
rect 23266 60958 23268 61010
rect 23212 60946 23268 60958
rect 22764 60788 22820 60798
rect 22764 60694 22820 60732
rect 23212 59780 23268 59790
rect 22764 59778 23268 59780
rect 22764 59726 23214 59778
rect 23266 59726 23268 59778
rect 22764 59724 23268 59726
rect 22764 59218 22820 59724
rect 23212 59714 23268 59724
rect 22764 59166 22766 59218
rect 22818 59166 22820 59218
rect 22764 59154 22820 59166
rect 23212 59108 23268 59118
rect 23436 59108 23492 63756
rect 23660 62188 23716 63756
rect 23268 59052 23492 59108
rect 23548 62132 23716 62188
rect 23884 62188 23940 63868
rect 24220 63924 24276 63934
rect 24220 62188 24276 63868
rect 24332 63922 24388 63934
rect 24332 63870 24334 63922
rect 24386 63870 24388 63922
rect 24332 63812 24388 63870
rect 24332 63746 24388 63756
rect 24332 63028 24388 63038
rect 24444 63028 24500 69244
rect 24780 66946 24836 66958
rect 24780 66894 24782 66946
rect 24834 66894 24836 66946
rect 24780 66834 24836 66894
rect 24780 66782 24782 66834
rect 24834 66782 24836 66834
rect 24780 66770 24836 66782
rect 24780 66612 24836 66622
rect 25228 66612 25284 70364
rect 25340 70326 25396 70364
rect 25676 70084 25732 70532
rect 25788 70308 25844 70814
rect 25900 70532 25956 71596
rect 26012 71586 26068 71596
rect 26796 70978 26852 72380
rect 26796 70926 26798 70978
rect 26850 70926 26852 70978
rect 26796 70914 26852 70926
rect 26460 70756 26516 70766
rect 25900 70466 25956 70476
rect 26236 70754 26516 70756
rect 26236 70702 26462 70754
rect 26514 70702 26516 70754
rect 26236 70700 26516 70702
rect 26236 70418 26292 70700
rect 26460 70644 26516 70700
rect 26460 70578 26516 70588
rect 27020 70532 27076 73892
rect 27244 73554 27300 73892
rect 27244 73502 27246 73554
rect 27298 73502 27300 73554
rect 27244 73490 27300 73502
rect 27580 73556 27636 74846
rect 27804 74338 27860 75292
rect 27804 74286 27806 74338
rect 27858 74286 27860 74338
rect 27804 74274 27860 74286
rect 27580 73490 27636 73500
rect 27804 74116 27860 74126
rect 27804 73108 27860 74060
rect 28028 73948 28084 77308
rect 28140 77298 28196 77308
rect 28364 77140 28420 77150
rect 28476 77140 28532 77756
rect 29260 77252 29316 77262
rect 29260 77158 29316 77196
rect 28364 77138 28532 77140
rect 28364 77086 28366 77138
rect 28418 77086 28532 77138
rect 28364 77084 28532 77086
rect 28364 76804 28420 77084
rect 28588 77028 28644 77038
rect 28364 76738 28420 76748
rect 28476 76972 28588 77028
rect 28364 76580 28420 76590
rect 28476 76580 28532 76972
rect 28588 76962 28644 76972
rect 29372 76580 29428 77980
rect 29484 77970 29540 77980
rect 29708 78034 29764 78046
rect 29708 77982 29710 78034
rect 29762 77982 29764 78034
rect 29708 77252 29764 77982
rect 29708 77186 29764 77196
rect 29708 77028 29764 77038
rect 29708 76934 29764 76972
rect 28364 76578 28532 76580
rect 28364 76526 28366 76578
rect 28418 76526 28532 76578
rect 28364 76524 28532 76526
rect 28812 76524 29428 76580
rect 28364 76514 28420 76524
rect 28252 76244 28308 76254
rect 28252 76150 28308 76188
rect 28700 75908 28756 75918
rect 28364 75572 28420 75582
rect 27804 73042 27860 73052
rect 27916 73892 28084 73948
rect 28140 74114 28196 74126
rect 28140 74062 28142 74114
rect 28194 74062 28196 74114
rect 28140 73948 28196 74062
rect 28364 74116 28420 75516
rect 28476 74898 28532 74910
rect 28476 74846 28478 74898
rect 28530 74846 28532 74898
rect 28476 74788 28532 74846
rect 28476 74722 28532 74732
rect 28364 74022 28420 74060
rect 28140 73892 28308 73948
rect 27804 72548 27860 72558
rect 27804 71762 27860 72492
rect 27804 71710 27806 71762
rect 27858 71710 27860 71762
rect 27356 70978 27412 70990
rect 27356 70926 27358 70978
rect 27410 70926 27412 70978
rect 26572 70476 27076 70532
rect 27132 70644 27188 70654
rect 26236 70366 26238 70418
rect 26290 70366 26292 70418
rect 26236 70354 26292 70366
rect 26460 70420 26516 70430
rect 26572 70420 26628 70476
rect 27132 70420 27188 70588
rect 26460 70418 26628 70420
rect 26460 70366 26462 70418
rect 26514 70366 26628 70418
rect 26460 70364 26628 70366
rect 26684 70364 27188 70420
rect 26460 70354 26516 70364
rect 25788 70242 25844 70252
rect 26684 70306 26740 70364
rect 26684 70254 26686 70306
rect 26738 70254 26740 70306
rect 26684 70242 26740 70254
rect 26124 70194 26180 70206
rect 26124 70142 26126 70194
rect 26178 70142 26180 70194
rect 25900 70084 25956 70094
rect 25676 70082 25956 70084
rect 25676 70030 25902 70082
rect 25954 70030 25956 70082
rect 25676 70028 25956 70030
rect 25900 70018 25956 70028
rect 26124 69412 26180 70142
rect 26796 70196 26852 70206
rect 27244 70196 27300 70206
rect 26796 70194 27300 70196
rect 26796 70142 26798 70194
rect 26850 70142 27246 70194
rect 27298 70142 27300 70194
rect 26796 70140 27300 70142
rect 26796 70130 26852 70140
rect 27244 70130 27300 70140
rect 26796 69972 26852 69982
rect 26796 69634 26852 69916
rect 27356 69972 27412 70926
rect 27692 70866 27748 70878
rect 27692 70814 27694 70866
rect 27746 70814 27748 70866
rect 27692 70756 27748 70814
rect 27468 70532 27524 70542
rect 27468 70418 27524 70476
rect 27468 70366 27470 70418
rect 27522 70366 27524 70418
rect 27468 70354 27524 70366
rect 27356 69906 27412 69916
rect 27580 70194 27636 70206
rect 27580 70142 27582 70194
rect 27634 70142 27636 70194
rect 26796 69582 26798 69634
rect 26850 69582 26852 69634
rect 26796 69570 26852 69582
rect 26124 69346 26180 69356
rect 26684 69412 26740 69422
rect 26684 69318 26740 69356
rect 27356 69410 27412 69422
rect 27356 69358 27358 69410
rect 27410 69358 27412 69410
rect 27356 69300 27412 69358
rect 27468 69300 27524 69310
rect 27356 69244 27468 69300
rect 27468 69234 27524 69244
rect 27580 68180 27636 70142
rect 27692 69410 27748 70700
rect 27804 70420 27860 71710
rect 27916 70754 27972 73892
rect 28140 73668 28196 73678
rect 28028 73108 28084 73118
rect 28028 70980 28084 73052
rect 28140 72436 28196 73612
rect 28252 73220 28308 73892
rect 28700 73554 28756 75852
rect 28700 73502 28702 73554
rect 28754 73502 28756 73554
rect 28700 73490 28756 73502
rect 28364 73332 28420 73342
rect 28364 73238 28420 73276
rect 28252 72770 28308 73164
rect 28252 72718 28254 72770
rect 28306 72718 28308 72770
rect 28252 72706 28308 72718
rect 28252 72436 28308 72446
rect 28196 72434 28308 72436
rect 28196 72382 28254 72434
rect 28306 72382 28308 72434
rect 28196 72380 28308 72382
rect 28140 72342 28196 72380
rect 28252 72370 28308 72380
rect 28364 72434 28420 72446
rect 28364 72382 28366 72434
rect 28418 72382 28420 72434
rect 28028 70866 28084 70924
rect 28028 70814 28030 70866
rect 28082 70814 28084 70866
rect 28028 70802 28084 70814
rect 28140 71652 28196 71662
rect 27916 70702 27918 70754
rect 27970 70702 27972 70754
rect 27916 70690 27972 70702
rect 28140 70644 28196 71596
rect 27804 70354 27860 70364
rect 28028 70588 28196 70644
rect 28252 70980 28308 70990
rect 27916 70194 27972 70206
rect 27916 70142 27918 70194
rect 27970 70142 27972 70194
rect 27916 69524 27972 70142
rect 27916 69458 27972 69468
rect 27692 69358 27694 69410
rect 27746 69358 27748 69410
rect 27692 69346 27748 69358
rect 27916 69300 27972 69310
rect 27916 69206 27972 69244
rect 27692 68180 27748 68190
rect 27580 68124 27692 68180
rect 27692 68114 27748 68124
rect 27020 67844 27076 67854
rect 27468 67844 27524 67854
rect 27020 67842 27524 67844
rect 27020 67790 27022 67842
rect 27074 67790 27470 67842
rect 27522 67790 27524 67842
rect 27020 67788 27524 67790
rect 26236 67732 26292 67742
rect 24836 66556 25284 66612
rect 25564 67730 26292 67732
rect 25564 67678 26238 67730
rect 26290 67678 26292 67730
rect 25564 67676 26292 67678
rect 24668 65380 24724 65390
rect 24556 65324 24668 65380
rect 24556 63922 24612 65324
rect 24668 65286 24724 65324
rect 24668 64596 24724 64606
rect 24668 64036 24724 64540
rect 24668 63970 24724 63980
rect 24556 63870 24558 63922
rect 24610 63870 24612 63922
rect 24556 63476 24612 63870
rect 24556 63420 24724 63476
rect 24556 63140 24612 63150
rect 24556 63046 24612 63084
rect 24388 62972 24500 63028
rect 24332 62962 24388 62972
rect 23884 62132 24052 62188
rect 24220 62132 24612 62188
rect 23212 59014 23268 59052
rect 22652 58772 22820 58828
rect 22764 57540 22820 58772
rect 23212 57652 23268 57662
rect 23212 57558 23268 57596
rect 22764 57446 22820 57484
rect 23548 57092 23604 62132
rect 23884 61348 23940 61358
rect 23884 61254 23940 61292
rect 23660 61012 23716 61022
rect 23660 60918 23716 60956
rect 23660 60002 23716 60014
rect 23660 59950 23662 60002
rect 23714 59950 23716 60002
rect 23660 59108 23716 59950
rect 23884 60004 23940 60014
rect 23884 59910 23940 59948
rect 23996 59220 24052 62132
rect 24444 61684 24500 61694
rect 24108 61682 24500 61684
rect 24108 61630 24446 61682
rect 24498 61630 24500 61682
rect 24108 61628 24500 61630
rect 24108 59892 24164 61628
rect 24444 61618 24500 61628
rect 24220 60788 24276 60798
rect 24220 60114 24276 60732
rect 24556 60228 24612 62132
rect 24668 60788 24724 63420
rect 24668 60722 24724 60732
rect 24668 60228 24724 60238
rect 24556 60226 24724 60228
rect 24556 60174 24670 60226
rect 24722 60174 24724 60226
rect 24556 60172 24724 60174
rect 24220 60062 24222 60114
rect 24274 60062 24276 60114
rect 24220 60050 24276 60062
rect 24668 60114 24724 60172
rect 24668 60062 24670 60114
rect 24722 60062 24724 60114
rect 24668 60004 24724 60062
rect 24668 59938 24724 59948
rect 24108 59890 24388 59892
rect 24108 59838 24110 59890
rect 24162 59838 24388 59890
rect 24108 59836 24388 59838
rect 24108 59826 24164 59836
rect 24332 59444 24388 59836
rect 24332 59388 24724 59444
rect 24444 59220 24500 59230
rect 23996 59218 24500 59220
rect 23996 59166 24446 59218
rect 24498 59166 24500 59218
rect 23996 59164 24500 59166
rect 23660 59042 23716 59052
rect 23772 59108 23828 59118
rect 23996 59108 24052 59164
rect 24444 59154 24500 59164
rect 24668 59218 24724 59388
rect 24668 59166 24670 59218
rect 24722 59166 24724 59218
rect 24668 59154 24724 59166
rect 23772 59106 24052 59108
rect 23772 59054 23774 59106
rect 23826 59054 24052 59106
rect 23772 59052 24052 59054
rect 23548 57026 23604 57036
rect 23772 56532 23828 59052
rect 24108 58994 24164 59006
rect 24108 58942 24110 58994
rect 24162 58942 24164 58994
rect 24108 57764 24164 58942
rect 24220 58548 24276 58558
rect 24220 58546 24388 58548
rect 24220 58494 24222 58546
rect 24274 58494 24388 58546
rect 24220 58492 24388 58494
rect 24220 58482 24276 58492
rect 24220 57764 24276 57774
rect 24108 57762 24276 57764
rect 24108 57710 24222 57762
rect 24274 57710 24276 57762
rect 24108 57708 24276 57710
rect 24220 57698 24276 57708
rect 24220 56756 24276 56766
rect 23548 56476 23828 56532
rect 23884 56754 24276 56756
rect 23884 56702 24222 56754
rect 24274 56702 24276 56754
rect 23884 56700 24276 56702
rect 23324 55412 23380 55422
rect 22596 55356 22820 55412
rect 22540 55318 22596 55356
rect 22204 54572 22484 54628
rect 21980 53442 22036 53452
rect 22092 53506 22148 53518
rect 22092 53454 22094 53506
rect 22146 53454 22148 53506
rect 21532 53058 21924 53060
rect 21532 53006 21534 53058
rect 21586 53006 21924 53058
rect 21532 53004 21924 53006
rect 22092 53058 22148 53454
rect 22092 53006 22094 53058
rect 22146 53006 22148 53058
rect 21532 52994 21588 53004
rect 22092 52994 22148 53006
rect 21980 52946 22036 52958
rect 21980 52894 21982 52946
rect 22034 52894 22036 52946
rect 21644 52836 21700 52846
rect 21420 52210 21476 52220
rect 21532 52724 21588 52734
rect 21308 52164 21364 52174
rect 21308 52070 21364 52108
rect 21532 52052 21588 52668
rect 21420 51996 21588 52052
rect 21420 50482 21476 51996
rect 21532 51490 21588 51502
rect 21532 51438 21534 51490
rect 21586 51438 21588 51490
rect 21532 50932 21588 51438
rect 21532 50866 21588 50876
rect 21420 50430 21422 50482
rect 21474 50430 21476 50482
rect 21420 50418 21476 50430
rect 21420 49364 21476 49374
rect 21420 49250 21476 49308
rect 21420 49198 21422 49250
rect 21474 49198 21476 49250
rect 21420 49186 21476 49198
rect 21644 48804 21700 52780
rect 21756 52052 21812 52062
rect 21756 50596 21812 51996
rect 21980 50708 22036 52894
rect 22092 52276 22148 52286
rect 22092 52182 22148 52220
rect 22204 51940 22260 54572
rect 22428 54402 22484 54414
rect 22428 54350 22430 54402
rect 22482 54350 22484 54402
rect 22428 53620 22484 54350
rect 22764 53844 22820 55356
rect 23324 55298 23380 55356
rect 23324 55246 23326 55298
rect 23378 55246 23380 55298
rect 23324 55234 23380 55246
rect 22876 54402 22932 54414
rect 22876 54350 22878 54402
rect 22930 54350 22932 54402
rect 22876 54292 22932 54350
rect 23436 54404 23492 54414
rect 23436 54310 23492 54348
rect 23100 54292 23156 54302
rect 22876 54236 23100 54292
rect 22876 53844 22932 53854
rect 22764 53842 22932 53844
rect 22764 53790 22878 53842
rect 22930 53790 22932 53842
rect 22764 53788 22932 53790
rect 22428 53618 22596 53620
rect 22428 53566 22430 53618
rect 22482 53566 22596 53618
rect 22428 53564 22596 53566
rect 22428 53554 22484 53564
rect 22316 53508 22372 53518
rect 22316 52388 22372 53452
rect 22316 52322 22372 52332
rect 22428 53170 22484 53182
rect 22428 53118 22430 53170
rect 22482 53118 22484 53170
rect 22204 50820 22260 51884
rect 22428 51380 22484 53118
rect 22428 51314 22484 51324
rect 22540 50932 22596 53564
rect 22540 50866 22596 50876
rect 22652 53058 22708 53070
rect 22652 53006 22654 53058
rect 22706 53006 22708 53058
rect 22204 50754 22260 50764
rect 21980 50642 22036 50652
rect 21756 50502 21812 50540
rect 22652 50428 22708 53006
rect 22764 52948 22820 53788
rect 22876 53778 22932 53788
rect 22764 52882 22820 52892
rect 22988 51380 23044 51390
rect 22988 51286 23044 51324
rect 22428 50370 22484 50382
rect 22428 50318 22430 50370
rect 22482 50318 22484 50370
rect 22316 49810 22372 49822
rect 22316 49758 22318 49810
rect 22370 49758 22372 49810
rect 22316 49028 22372 49758
rect 21644 48738 21700 48748
rect 22092 48914 22148 48926
rect 22092 48862 22094 48914
rect 22146 48862 22148 48914
rect 21980 48580 22036 48590
rect 21196 48190 21198 48242
rect 21250 48190 21252 48242
rect 21196 44660 21252 48190
rect 21868 48244 21924 48254
rect 21868 48150 21924 48188
rect 21644 48018 21700 48030
rect 21644 47966 21646 48018
rect 21698 47966 21700 48018
rect 21532 47124 21588 47134
rect 21532 46674 21588 47068
rect 21532 46622 21534 46674
rect 21586 46622 21588 46674
rect 21532 46610 21588 46622
rect 21532 45890 21588 45902
rect 21532 45838 21534 45890
rect 21586 45838 21588 45890
rect 21532 45108 21588 45838
rect 21308 44884 21364 44894
rect 21308 44790 21364 44828
rect 21196 44594 21252 44604
rect 21532 44548 21588 45052
rect 21532 44482 21588 44492
rect 21644 45220 21700 47966
rect 21868 47458 21924 47470
rect 21868 47406 21870 47458
rect 21922 47406 21924 47458
rect 21308 44324 21364 44334
rect 21308 44230 21364 44268
rect 21532 44210 21588 44222
rect 21532 44158 21534 44210
rect 21586 44158 21588 44210
rect 21532 44100 21588 44158
rect 21084 44044 21588 44100
rect 21084 37268 21140 44044
rect 21196 43876 21252 43886
rect 21252 43820 21476 43876
rect 21196 43810 21252 43820
rect 21308 42868 21364 42878
rect 21308 42754 21364 42812
rect 21308 42702 21310 42754
rect 21362 42702 21364 42754
rect 21308 42690 21364 42702
rect 21420 41298 21476 43820
rect 21644 43540 21700 45164
rect 21644 42868 21700 43484
rect 21532 42812 21700 42868
rect 21756 46676 21812 46686
rect 21756 46002 21812 46620
rect 21756 45950 21758 46002
rect 21810 45950 21812 46002
rect 21532 42810 21588 42812
rect 21532 42758 21534 42810
rect 21586 42758 21588 42810
rect 21532 42746 21588 42758
rect 21756 42754 21812 45950
rect 21868 44436 21924 47406
rect 21980 46674 22036 48524
rect 21980 46622 21982 46674
rect 22034 46622 22036 46674
rect 21980 45892 22036 46622
rect 22092 48244 22148 48862
rect 22316 48580 22372 48972
rect 22316 48514 22372 48524
rect 22092 46676 22148 48188
rect 22204 48130 22260 48142
rect 22204 48078 22206 48130
rect 22258 48078 22260 48130
rect 22204 47124 22260 48078
rect 22204 47058 22260 47068
rect 22092 46610 22148 46620
rect 21980 45826 22036 45836
rect 22316 46562 22372 46574
rect 22316 46510 22318 46562
rect 22370 46510 22372 46562
rect 22092 45780 22148 45790
rect 21868 44370 21924 44380
rect 21980 45332 22036 45342
rect 21980 43538 22036 45276
rect 21980 43486 21982 43538
rect 22034 43486 22036 43538
rect 21868 43316 21924 43326
rect 21868 43222 21924 43260
rect 21756 42702 21758 42754
rect 21810 42702 21812 42754
rect 21756 42690 21812 42702
rect 21868 42196 21924 42206
rect 21532 42084 21588 42094
rect 21588 42028 21700 42084
rect 21532 42018 21588 42028
rect 21644 41970 21700 42028
rect 21644 41918 21646 41970
rect 21698 41918 21700 41970
rect 21644 41748 21700 41918
rect 21868 41970 21924 42140
rect 21868 41918 21870 41970
rect 21922 41918 21924 41970
rect 21868 41860 21924 41918
rect 21980 41972 22036 43486
rect 22092 43540 22148 45724
rect 22204 45332 22260 45342
rect 22204 44210 22260 45276
rect 22204 44158 22206 44210
rect 22258 44158 22260 44210
rect 22204 44146 22260 44158
rect 22204 43540 22260 43550
rect 22092 43484 22204 43540
rect 22204 43474 22260 43484
rect 22092 42532 22148 42542
rect 22092 42530 22260 42532
rect 22092 42478 22094 42530
rect 22146 42478 22260 42530
rect 22092 42476 22260 42478
rect 22092 42466 22148 42476
rect 22092 41972 22148 41982
rect 21980 41970 22148 41972
rect 21980 41918 22094 41970
rect 22146 41918 22148 41970
rect 21980 41916 22148 41918
rect 21868 41804 22036 41860
rect 21644 41682 21700 41692
rect 21420 41246 21422 41298
rect 21474 41246 21476 41298
rect 21420 41234 21476 41246
rect 21532 41300 21588 41310
rect 21980 41300 22036 41804
rect 22092 41524 22148 41916
rect 22092 41458 22148 41468
rect 21980 41244 22148 41300
rect 21308 41188 21364 41198
rect 21308 41094 21364 41132
rect 21532 41186 21588 41244
rect 21532 41134 21534 41186
rect 21586 41134 21588 41186
rect 21532 41122 21588 41134
rect 21868 41188 21924 41198
rect 21756 40962 21812 40974
rect 21756 40910 21758 40962
rect 21810 40910 21812 40962
rect 21196 40514 21252 40526
rect 21196 40462 21198 40514
rect 21250 40462 21252 40514
rect 21196 39620 21252 40462
rect 21756 40404 21812 40910
rect 21756 40338 21812 40348
rect 21196 39564 21588 39620
rect 21532 38948 21588 39564
rect 21868 39618 21924 41132
rect 21868 39566 21870 39618
rect 21922 39566 21924 39618
rect 21868 39554 21924 39566
rect 21980 41074 22036 41086
rect 21980 41022 21982 41074
rect 22034 41022 22036 41074
rect 21644 39508 21700 39518
rect 21644 39414 21700 39452
rect 21644 38948 21700 38958
rect 21532 38946 21700 38948
rect 21532 38894 21646 38946
rect 21698 38894 21700 38946
rect 21532 38892 21700 38894
rect 21644 38882 21700 38892
rect 21644 38724 21700 38734
rect 21644 38612 21812 38668
rect 21644 37940 21700 37950
rect 21644 37380 21700 37884
rect 21756 37604 21812 38612
rect 21868 37940 21924 37950
rect 21868 37846 21924 37884
rect 21756 37548 21924 37604
rect 21868 37490 21924 37548
rect 21868 37438 21870 37490
rect 21922 37438 21924 37490
rect 21868 37426 21924 37438
rect 21756 37380 21812 37390
rect 21644 37324 21756 37380
rect 21756 37314 21812 37324
rect 21084 37202 21140 37212
rect 21308 37154 21364 37166
rect 21308 37102 21310 37154
rect 21362 37102 21364 37154
rect 20916 35868 21028 35924
rect 21084 37044 21140 37054
rect 20860 35830 20916 35868
rect 20972 34020 21028 34030
rect 21084 34020 21140 36988
rect 21308 36260 21364 37102
rect 21532 36260 21588 36270
rect 21308 36204 21532 36260
rect 21532 36166 21588 36204
rect 20972 34018 21140 34020
rect 20972 33966 20974 34018
rect 21026 33966 21140 34018
rect 20972 33964 21140 33966
rect 20748 33572 20804 33582
rect 20748 33458 20804 33516
rect 20748 33406 20750 33458
rect 20802 33406 20804 33458
rect 20748 33394 20804 33406
rect 20972 33348 21028 33964
rect 21868 33572 21924 33582
rect 21868 33458 21924 33516
rect 21868 33406 21870 33458
rect 21922 33406 21924 33458
rect 21868 33394 21924 33406
rect 21644 33348 21700 33358
rect 20972 33346 21700 33348
rect 20972 33294 21646 33346
rect 21698 33294 21700 33346
rect 20972 33292 21700 33294
rect 21308 33124 21364 33134
rect 21196 33122 21364 33124
rect 21196 33070 21310 33122
rect 21362 33070 21364 33122
rect 21196 33068 21364 33070
rect 21196 32562 21252 33068
rect 21308 33058 21364 33068
rect 21196 32510 21198 32562
rect 21250 32510 21252 32562
rect 21196 32498 21252 32510
rect 21420 32674 21476 32686
rect 21420 32622 21422 32674
rect 21474 32622 21476 32674
rect 21308 31890 21364 31902
rect 21308 31838 21310 31890
rect 21362 31838 21364 31890
rect 21308 31780 21364 31838
rect 21420 31892 21476 32622
rect 21420 31826 21476 31836
rect 21308 31714 21364 31724
rect 21196 29428 21252 29438
rect 21196 29334 21252 29372
rect 21644 29204 21700 33292
rect 21980 31780 22036 41022
rect 22092 40740 22148 41244
rect 22092 40626 22148 40684
rect 22092 40574 22094 40626
rect 22146 40574 22148 40626
rect 22092 40562 22148 40574
rect 22204 40068 22260 42476
rect 22316 41188 22372 46510
rect 22428 41972 22484 50318
rect 22540 50372 22708 50428
rect 23100 50428 23156 54236
rect 23548 54292 23604 56476
rect 23884 56306 23940 56700
rect 24220 56690 24276 56700
rect 23884 56254 23886 56306
rect 23938 56254 23940 56306
rect 23884 56242 23940 56254
rect 23660 56084 23716 56094
rect 23660 56082 23940 56084
rect 23660 56030 23662 56082
rect 23714 56030 23940 56082
rect 23660 56028 23940 56030
rect 23660 56018 23716 56028
rect 23884 54738 23940 56028
rect 24220 55410 24276 55422
rect 24220 55358 24222 55410
rect 24274 55358 24276 55410
rect 24220 55076 24276 55358
rect 24220 55010 24276 55020
rect 23884 54686 23886 54738
rect 23938 54686 23940 54738
rect 23884 54674 23940 54686
rect 23548 54226 23604 54236
rect 24220 54292 24276 54302
rect 24220 54198 24276 54236
rect 23436 53508 23492 53518
rect 23436 53414 23492 53452
rect 23660 53172 23716 53182
rect 23436 52834 23492 52846
rect 23436 52782 23438 52834
rect 23490 52782 23492 52834
rect 23436 52500 23492 52782
rect 23436 52434 23492 52444
rect 23436 51940 23492 51950
rect 23436 50706 23492 51884
rect 23548 51492 23604 51502
rect 23548 51398 23604 51436
rect 23436 50654 23438 50706
rect 23490 50654 23492 50706
rect 23436 50484 23492 50654
rect 23100 50372 23268 50428
rect 23436 50418 23492 50428
rect 22540 47012 22596 50372
rect 23100 50148 23156 50158
rect 22988 49700 23044 49710
rect 22652 49026 22708 49038
rect 22876 49028 22932 49038
rect 22652 48974 22654 49026
rect 22706 48974 22708 49026
rect 22652 48804 22708 48974
rect 22652 48738 22708 48748
rect 22764 49026 22932 49028
rect 22764 48974 22878 49026
rect 22930 48974 22932 49026
rect 22764 48972 22932 48974
rect 22764 48692 22820 48972
rect 22876 48962 22932 48972
rect 22988 48692 23044 49644
rect 23100 48916 23156 50092
rect 23100 48822 23156 48860
rect 22764 48626 22820 48636
rect 22876 48636 23044 48692
rect 22652 48244 22708 48254
rect 22652 48150 22708 48188
rect 22540 46956 22708 47012
rect 22540 44436 22596 44446
rect 22540 44342 22596 44380
rect 22652 43652 22708 46956
rect 22876 45892 22932 48636
rect 22988 48468 23044 48478
rect 22988 48354 23044 48412
rect 22988 48302 22990 48354
rect 23042 48302 23044 48354
rect 22988 48290 23044 48302
rect 22876 45826 22932 45836
rect 23100 48130 23156 48142
rect 23100 48078 23102 48130
rect 23154 48078 23156 48130
rect 22764 45780 22820 45790
rect 22764 45686 22820 45724
rect 22876 45556 22932 45566
rect 22652 43586 22708 43596
rect 22764 45500 22876 45556
rect 22540 43540 22596 43550
rect 22540 43428 22596 43484
rect 22540 43372 22708 43428
rect 22540 43092 22596 43102
rect 22540 42642 22596 43036
rect 22540 42590 22542 42642
rect 22594 42590 22596 42642
rect 22540 42578 22596 42590
rect 22428 41906 22484 41916
rect 22316 41122 22372 41132
rect 22428 41746 22484 41758
rect 22428 41694 22430 41746
rect 22482 41694 22484 41746
rect 22316 40964 22372 40974
rect 22316 40870 22372 40908
rect 22428 40852 22484 41694
rect 22652 41636 22708 43372
rect 22652 41570 22708 41580
rect 22428 40786 22484 40796
rect 22652 41412 22708 41422
rect 22652 40516 22708 41356
rect 22652 40450 22708 40460
rect 22540 40292 22596 40302
rect 22540 40198 22596 40236
rect 22204 40002 22260 40012
rect 22764 39842 22820 45500
rect 22876 45490 22932 45500
rect 23100 45332 23156 48078
rect 23212 45444 23268 50372
rect 23324 49924 23380 49934
rect 23324 49830 23380 49868
rect 23548 49924 23604 49934
rect 23212 45378 23268 45388
rect 23324 46788 23380 46798
rect 23100 45266 23156 45276
rect 23212 45220 23268 45230
rect 23324 45220 23380 46732
rect 23548 46004 23604 49868
rect 23660 48692 23716 53116
rect 23884 52834 23940 52846
rect 23884 52782 23886 52834
rect 23938 52782 23940 52834
rect 23884 52724 23940 52782
rect 23884 52658 23940 52668
rect 23660 48626 23716 48636
rect 23772 52612 23828 52622
rect 23660 48356 23716 48366
rect 23660 48130 23716 48300
rect 23660 48078 23662 48130
rect 23714 48078 23716 48130
rect 23660 47348 23716 48078
rect 23660 47282 23716 47292
rect 23660 46788 23716 46826
rect 23660 46722 23716 46732
rect 23212 45218 23380 45220
rect 23212 45166 23214 45218
rect 23266 45166 23380 45218
rect 23212 45164 23380 45166
rect 23212 45154 23268 45164
rect 22876 44324 22932 44334
rect 22876 41860 22932 44268
rect 23212 43764 23268 43774
rect 23212 43538 23268 43708
rect 23212 43486 23214 43538
rect 23266 43486 23268 43538
rect 23212 43092 23268 43486
rect 23212 43026 23268 43036
rect 23324 42082 23380 45164
rect 23436 45948 23604 46004
rect 23660 46004 23716 46014
rect 23436 45108 23492 45948
rect 23436 44324 23492 45052
rect 23548 45778 23604 45790
rect 23548 45726 23550 45778
rect 23602 45726 23604 45778
rect 23548 44548 23604 45726
rect 23660 45778 23716 45948
rect 23660 45726 23662 45778
rect 23714 45726 23716 45778
rect 23660 45714 23716 45726
rect 23772 45444 23828 52556
rect 24220 52274 24276 52286
rect 24220 52222 24222 52274
rect 24274 52222 24276 52274
rect 23996 52164 24052 52174
rect 23996 50596 24052 52108
rect 23996 50530 24052 50540
rect 24220 50428 24276 52222
rect 23996 50372 24276 50428
rect 23884 48244 23940 48254
rect 23884 48150 23940 48188
rect 23884 45780 23940 45790
rect 23884 45686 23940 45724
rect 23772 45388 23940 45444
rect 23772 45220 23828 45230
rect 23660 45108 23716 45118
rect 23660 45014 23716 45052
rect 23772 45106 23828 45164
rect 23772 45054 23774 45106
rect 23826 45054 23828 45106
rect 23772 45042 23828 45054
rect 23548 44482 23604 44492
rect 23436 44268 23716 44324
rect 23660 44210 23716 44268
rect 23660 44158 23662 44210
rect 23714 44158 23716 44210
rect 23660 44146 23716 44158
rect 23772 43876 23828 43886
rect 23884 43876 23940 45388
rect 23828 43820 23940 43876
rect 23324 42030 23326 42082
rect 23378 42030 23380 42082
rect 23324 41972 23380 42030
rect 23100 41916 23380 41972
rect 23436 43650 23492 43662
rect 23436 43598 23438 43650
rect 23490 43598 23492 43650
rect 23436 43540 23492 43598
rect 23660 43652 23716 43662
rect 23660 43558 23716 43596
rect 23772 43650 23828 43820
rect 23996 43764 24052 50372
rect 24220 49812 24276 49822
rect 24108 48916 24164 48926
rect 24108 46676 24164 48860
rect 24220 48466 24276 49756
rect 24220 48414 24222 48466
rect 24274 48414 24276 48466
rect 24220 48402 24276 48414
rect 24220 47012 24276 47022
rect 24220 46898 24276 46956
rect 24220 46846 24222 46898
rect 24274 46846 24276 46898
rect 24220 46834 24276 46846
rect 24108 46610 24164 46620
rect 24108 45890 24164 45902
rect 24108 45838 24110 45890
rect 24162 45838 24164 45890
rect 24108 44436 24164 45838
rect 24220 45778 24276 45790
rect 24220 45726 24222 45778
rect 24274 45726 24276 45778
rect 24220 45556 24276 45726
rect 24220 45490 24276 45500
rect 24220 44884 24276 44894
rect 24220 44790 24276 44828
rect 24108 44370 24164 44380
rect 24332 43764 24388 58492
rect 24668 58436 24724 58446
rect 24668 58342 24724 58380
rect 24556 57762 24612 57774
rect 24556 57710 24558 57762
rect 24610 57710 24612 57762
rect 24556 56980 24612 57710
rect 24556 56914 24612 56924
rect 24668 56868 24724 56878
rect 24556 55188 24612 55198
rect 24556 55094 24612 55132
rect 24444 54404 24500 54414
rect 24444 45892 24500 54348
rect 24668 54180 24724 56812
rect 24556 54124 24724 54180
rect 24556 51602 24612 54124
rect 24668 52164 24724 52174
rect 24668 52070 24724 52108
rect 24556 51550 24558 51602
rect 24610 51550 24612 51602
rect 24556 51538 24612 51550
rect 24668 50482 24724 50494
rect 24444 45826 24500 45836
rect 24556 50428 24612 50438
rect 24556 49810 24612 50372
rect 24556 49758 24558 49810
rect 24610 49758 24612 49810
rect 24556 45780 24612 49758
rect 24668 50430 24670 50482
rect 24722 50430 24724 50482
rect 24668 49364 24724 50430
rect 24668 49298 24724 49308
rect 24668 48580 24724 48590
rect 24668 48466 24724 48524
rect 24668 48414 24670 48466
rect 24722 48414 24724 48466
rect 24668 48402 24724 48414
rect 24780 47570 24836 66556
rect 24892 66386 24948 66398
rect 24892 66334 24894 66386
rect 24946 66334 24948 66386
rect 24892 65492 24948 66334
rect 25228 66164 25284 66174
rect 25228 66162 25508 66164
rect 25228 66110 25230 66162
rect 25282 66110 25508 66162
rect 25228 66108 25508 66110
rect 25228 66098 25284 66108
rect 25452 65828 25508 66108
rect 25564 66162 25620 67676
rect 26236 67666 26292 67676
rect 26012 66724 26068 66734
rect 26012 66388 26068 66668
rect 26012 66294 26068 66332
rect 27020 66388 27076 67788
rect 27468 67778 27524 67788
rect 25564 66110 25566 66162
rect 25618 66110 25620 66162
rect 25564 66098 25620 66110
rect 26348 66164 26404 66174
rect 25452 65772 25844 65828
rect 25788 65714 25844 65772
rect 25788 65662 25790 65714
rect 25842 65662 25844 65714
rect 25788 65650 25844 65662
rect 24892 65426 24948 65436
rect 25228 65492 25284 65502
rect 25228 65398 25284 65436
rect 25116 65380 25172 65390
rect 24892 65268 24948 65278
rect 24892 64706 24948 65212
rect 25116 64820 25172 65324
rect 25564 65380 25620 65390
rect 25340 65268 25396 65278
rect 25340 64820 25396 65212
rect 25452 65268 25508 65278
rect 25564 65268 25620 65324
rect 26236 65380 26292 65390
rect 26236 65286 26292 65324
rect 25452 65266 25620 65268
rect 25452 65214 25454 65266
rect 25506 65214 25620 65266
rect 25452 65212 25620 65214
rect 25452 65202 25508 65212
rect 25452 64820 25508 64830
rect 25116 64818 25284 64820
rect 25116 64766 25118 64818
rect 25170 64766 25284 64818
rect 25116 64764 25284 64766
rect 25340 64818 25508 64820
rect 25340 64766 25454 64818
rect 25506 64766 25508 64818
rect 25340 64764 25508 64766
rect 25116 64754 25172 64764
rect 24892 64654 24894 64706
rect 24946 64654 24948 64706
rect 24892 64642 24948 64654
rect 25228 64148 25284 64764
rect 25452 64754 25508 64764
rect 25564 64708 25620 65212
rect 26348 64930 26404 66108
rect 26684 65380 26740 65390
rect 26684 65286 26740 65324
rect 26348 64878 26350 64930
rect 26402 64878 26404 64930
rect 26348 64866 26404 64878
rect 25676 64708 25732 64718
rect 25564 64706 25732 64708
rect 25564 64654 25678 64706
rect 25730 64654 25732 64706
rect 25564 64652 25732 64654
rect 25340 64148 25396 64158
rect 25228 64146 25396 64148
rect 25228 64094 25342 64146
rect 25394 64094 25396 64146
rect 25228 64092 25396 64094
rect 25340 64082 25396 64092
rect 25564 64148 25620 64652
rect 25676 64642 25732 64652
rect 26460 64594 26516 64606
rect 26460 64542 26462 64594
rect 26514 64542 26516 64594
rect 26012 64484 26068 64494
rect 25564 64082 25620 64092
rect 25676 64482 26068 64484
rect 25676 64430 26014 64482
rect 26066 64430 26068 64482
rect 25676 64428 26068 64430
rect 25228 63026 25284 63038
rect 25228 62974 25230 63026
rect 25282 62974 25284 63026
rect 25228 61012 25284 62974
rect 25676 62354 25732 64428
rect 26012 64418 26068 64428
rect 26236 64372 26292 64382
rect 26236 64146 26292 64316
rect 26236 64094 26238 64146
rect 26290 64094 26292 64146
rect 26236 64082 26292 64094
rect 25788 63922 25844 63934
rect 25788 63870 25790 63922
rect 25842 63870 25844 63922
rect 25788 63028 25844 63870
rect 26460 63812 26516 64542
rect 26908 64484 26964 64494
rect 26908 64390 26964 64428
rect 26460 63746 26516 63756
rect 26684 63810 26740 63822
rect 26684 63758 26686 63810
rect 26738 63758 26740 63810
rect 25788 62962 25844 62972
rect 26684 63700 26740 63758
rect 26684 62580 26740 63644
rect 27020 63140 27076 66332
rect 28028 64818 28084 70588
rect 28140 70420 28196 70430
rect 28140 70326 28196 70364
rect 28252 70306 28308 70924
rect 28252 70254 28254 70306
rect 28306 70254 28308 70306
rect 28140 70196 28196 70206
rect 28140 68852 28196 70140
rect 28252 69300 28308 70254
rect 28364 70084 28420 72382
rect 28812 70196 28868 76524
rect 29596 76468 29652 76478
rect 29596 76374 29652 76412
rect 29148 76354 29204 76366
rect 29148 76302 29150 76354
rect 29202 76302 29204 76354
rect 29036 76242 29092 76254
rect 29036 76190 29038 76242
rect 29090 76190 29092 76242
rect 29036 75010 29092 76190
rect 29148 76020 29204 76302
rect 29148 75954 29204 75964
rect 29708 76244 29764 76254
rect 29260 75796 29316 75806
rect 29260 75702 29316 75740
rect 29036 74958 29038 75010
rect 29090 74958 29092 75010
rect 29036 74946 29092 74958
rect 29148 74898 29204 74910
rect 29148 74846 29150 74898
rect 29202 74846 29204 74898
rect 29036 73890 29092 73902
rect 29036 73838 29038 73890
rect 29090 73838 29092 73890
rect 29036 73332 29092 73838
rect 29036 73238 29092 73276
rect 28924 71204 28980 71214
rect 28924 70306 28980 71148
rect 29148 70420 29204 74846
rect 29596 74900 29652 74910
rect 29260 74788 29316 74798
rect 29260 74694 29316 74732
rect 29260 74116 29316 74126
rect 29260 74002 29316 74060
rect 29260 73950 29262 74002
rect 29314 73950 29316 74002
rect 29260 73668 29316 73950
rect 29260 73602 29316 73612
rect 29372 74002 29428 74014
rect 29372 73950 29374 74002
rect 29426 73950 29428 74002
rect 29260 73218 29316 73230
rect 29260 73166 29262 73218
rect 29314 73166 29316 73218
rect 29260 73108 29316 73166
rect 29260 73042 29316 73052
rect 29372 72546 29428 73950
rect 29372 72494 29374 72546
rect 29426 72494 29428 72546
rect 29260 72434 29316 72446
rect 29260 72382 29262 72434
rect 29314 72382 29316 72434
rect 29260 71204 29316 72382
rect 29372 71540 29428 72494
rect 29596 73330 29652 74844
rect 29708 74338 29764 76188
rect 29820 76020 29876 82348
rect 29932 81956 29988 81966
rect 29932 81954 30100 81956
rect 29932 81902 29934 81954
rect 29986 81902 30100 81954
rect 29932 81900 30100 81902
rect 29932 81890 29988 81900
rect 29932 80948 29988 80958
rect 29932 80854 29988 80892
rect 30044 80612 30100 81900
rect 30268 81172 30324 82572
rect 30380 82292 30436 84814
rect 30604 84644 30660 84654
rect 30604 84530 30660 84588
rect 30604 84478 30606 84530
rect 30658 84478 30660 84530
rect 30604 84466 30660 84478
rect 30492 83636 30548 83646
rect 30492 83542 30548 83580
rect 30604 83188 30660 83198
rect 30604 82964 30660 83132
rect 30380 81396 30436 82236
rect 30380 81330 30436 81340
rect 30492 82962 30660 82964
rect 30492 82910 30606 82962
rect 30658 82910 30660 82962
rect 30492 82908 30660 82910
rect 30268 81116 30436 81172
rect 29932 80556 30100 80612
rect 30268 80946 30324 80958
rect 30268 80894 30270 80946
rect 30322 80894 30324 80946
rect 29932 77924 29988 80556
rect 30044 80386 30100 80398
rect 30044 80334 30046 80386
rect 30098 80334 30100 80386
rect 30044 78820 30100 80334
rect 30268 79492 30324 80894
rect 30268 79426 30324 79436
rect 30380 79268 30436 81116
rect 30492 81060 30548 82908
rect 30604 82898 30660 82908
rect 30604 81954 30660 81966
rect 30604 81902 30606 81954
rect 30658 81902 30660 81954
rect 30604 81172 30660 81902
rect 30716 81956 30772 85708
rect 31052 85652 31444 85708
rect 31500 86098 31556 86110
rect 31500 86046 31502 86098
rect 31554 86046 31556 86098
rect 31500 85708 31556 86046
rect 31612 85986 31668 86268
rect 31612 85934 31614 85986
rect 31666 85934 31668 85986
rect 31612 85922 31668 85934
rect 31500 85652 31668 85708
rect 30828 85204 30884 85214
rect 30828 85110 30884 85148
rect 31052 84644 31108 84654
rect 31052 84530 31108 84588
rect 31052 84478 31054 84530
rect 31106 84478 31108 84530
rect 31052 84466 31108 84478
rect 30940 83300 30996 83310
rect 30940 83206 30996 83244
rect 31164 82626 31220 85652
rect 31276 85092 31332 85102
rect 31276 84998 31332 85036
rect 31612 85090 31668 85652
rect 31724 85202 31780 86494
rect 31836 85874 31892 85886
rect 31836 85822 31838 85874
rect 31890 85822 31892 85874
rect 31836 85764 31892 85822
rect 31836 85698 31892 85708
rect 31724 85150 31726 85202
rect 31778 85150 31780 85202
rect 31724 85138 31780 85150
rect 31948 85316 32004 87164
rect 31612 85038 31614 85090
rect 31666 85038 31668 85090
rect 31612 85026 31668 85038
rect 31836 85092 31892 85102
rect 31948 85092 32004 85260
rect 31836 85090 32004 85092
rect 31836 85038 31838 85090
rect 31890 85038 32004 85090
rect 31836 85036 32004 85038
rect 32060 85092 32116 87388
rect 32508 87330 32564 87950
rect 35084 88004 35140 90636
rect 35196 90188 35460 90198
rect 35252 90132 35300 90188
rect 35356 90132 35404 90188
rect 35196 90122 35460 90132
rect 37884 89010 37940 92206
rect 38220 92146 38276 92158
rect 38220 92094 38222 92146
rect 38274 92094 38276 92146
rect 38220 92036 38276 92094
rect 38220 91476 38276 91980
rect 38220 91410 38276 91420
rect 37884 88958 37886 89010
rect 37938 88958 37940 89010
rect 37884 88946 37940 88958
rect 36540 88898 36596 88910
rect 36540 88846 36542 88898
rect 36594 88846 36596 88898
rect 35196 88620 35460 88630
rect 35252 88564 35300 88620
rect 35356 88564 35404 88620
rect 35196 88554 35460 88564
rect 35644 88116 35700 88126
rect 35644 88114 35812 88116
rect 35644 88062 35646 88114
rect 35698 88062 35812 88114
rect 35644 88060 35812 88062
rect 35644 88050 35700 88060
rect 35084 87910 35140 87948
rect 35308 88004 35364 88014
rect 35532 88004 35588 88014
rect 35308 88002 35476 88004
rect 35308 87950 35310 88002
rect 35362 87950 35476 88002
rect 35308 87948 35476 87950
rect 35308 87938 35364 87948
rect 35420 87556 35476 87948
rect 35532 87910 35588 87948
rect 35644 87556 35700 87566
rect 35420 87554 35700 87556
rect 35420 87502 35646 87554
rect 35698 87502 35700 87554
rect 35420 87500 35700 87502
rect 35644 87490 35700 87500
rect 32956 87444 33012 87454
rect 32956 87350 33012 87388
rect 33404 87442 33460 87454
rect 33404 87390 33406 87442
rect 33458 87390 33460 87442
rect 32508 87278 32510 87330
rect 32562 87278 32564 87330
rect 32508 86658 32564 87278
rect 32844 86772 32900 86782
rect 32844 86770 33012 86772
rect 32844 86718 32846 86770
rect 32898 86718 33012 86770
rect 32844 86716 33012 86718
rect 32844 86706 32900 86716
rect 32508 86606 32510 86658
rect 32562 86606 32564 86658
rect 32508 85764 32564 86606
rect 32508 85670 32564 85708
rect 32844 86100 32900 86110
rect 32508 85316 32564 85326
rect 32508 85222 32564 85260
rect 32844 85314 32900 86044
rect 32956 85764 33012 86716
rect 33404 85876 33460 87390
rect 33628 87442 33684 87454
rect 33628 87390 33630 87442
rect 33682 87390 33684 87442
rect 33516 87332 33572 87342
rect 33516 87238 33572 87276
rect 33628 86100 33684 87390
rect 33628 86034 33684 86044
rect 34524 87444 34580 87454
rect 34860 87444 34916 87454
rect 34524 87442 34916 87444
rect 34524 87390 34526 87442
rect 34578 87390 34862 87442
rect 34914 87390 34916 87442
rect 34524 87388 34916 87390
rect 33628 85876 33684 85886
rect 33404 85874 33684 85876
rect 33404 85822 33630 85874
rect 33682 85822 33684 85874
rect 33404 85820 33684 85822
rect 33068 85764 33124 85774
rect 32956 85762 33124 85764
rect 32956 85710 33070 85762
rect 33122 85710 33124 85762
rect 32956 85708 33124 85710
rect 32844 85262 32846 85314
rect 32898 85262 32900 85314
rect 32844 85250 32900 85262
rect 31836 85026 31892 85036
rect 32060 84978 32116 85036
rect 32060 84926 32062 84978
rect 32114 84926 32116 84978
rect 32060 84914 32116 84926
rect 31500 84868 31556 84878
rect 31388 83412 31444 83422
rect 31388 83318 31444 83356
rect 31164 82574 31166 82626
rect 31218 82574 31220 82626
rect 31164 82292 31220 82574
rect 31388 82516 31444 82526
rect 31500 82516 31556 84812
rect 32732 84868 32788 84878
rect 33068 84868 33124 85708
rect 33292 85650 33348 85662
rect 33292 85598 33294 85650
rect 33346 85598 33348 85650
rect 33292 85316 33348 85598
rect 33292 85250 33348 85260
rect 33628 85092 33684 85820
rect 33628 85026 33684 85036
rect 33852 85540 33908 85550
rect 32788 84812 33124 84868
rect 32732 84774 32788 84812
rect 33852 84194 33908 85484
rect 34524 85540 34580 87388
rect 34860 87378 34916 87388
rect 34972 87332 35028 87342
rect 34972 86770 35028 87276
rect 35196 87052 35460 87062
rect 35252 86996 35300 87052
rect 35356 86996 35404 87052
rect 35196 86986 35460 86996
rect 34972 86718 34974 86770
rect 35026 86718 35028 86770
rect 34972 86706 35028 86718
rect 35644 86660 35700 86670
rect 35532 86658 35700 86660
rect 35532 86606 35646 86658
rect 35698 86606 35700 86658
rect 35532 86604 35700 86606
rect 34972 85876 35028 85886
rect 34860 85874 35028 85876
rect 34860 85822 34974 85874
rect 35026 85822 35028 85874
rect 34860 85820 35028 85822
rect 34860 85708 34916 85820
rect 34972 85810 35028 85820
rect 34524 85474 34580 85484
rect 34748 85652 34916 85708
rect 35084 85762 35140 85774
rect 35084 85710 35086 85762
rect 35138 85710 35140 85762
rect 34748 85204 34804 85652
rect 34412 85092 34468 85102
rect 34412 84998 34468 85036
rect 33964 84866 34020 84878
rect 33964 84814 33966 84866
rect 34018 84814 34020 84866
rect 33964 84756 34020 84814
rect 34524 84866 34580 84878
rect 34748 84868 34804 85148
rect 35084 85092 35140 85710
rect 35196 85484 35460 85494
rect 35252 85428 35300 85484
rect 35356 85428 35404 85484
rect 35196 85418 35460 85428
rect 35084 85026 35140 85036
rect 34524 84814 34526 84866
rect 34578 84814 34580 84866
rect 34020 84700 34244 84756
rect 33964 84690 34020 84700
rect 34188 84530 34244 84700
rect 34188 84478 34190 84530
rect 34242 84478 34244 84530
rect 34188 84466 34244 84478
rect 33852 84142 33854 84194
rect 33906 84142 33908 84194
rect 31948 84084 32004 84094
rect 31612 82628 31668 82638
rect 31612 82534 31668 82572
rect 31388 82514 31556 82516
rect 31388 82462 31390 82514
rect 31442 82462 31556 82514
rect 31388 82460 31556 82462
rect 31388 82450 31444 82460
rect 31164 82236 31444 82292
rect 31164 81956 31220 81966
rect 30716 81954 31220 81956
rect 30716 81902 31166 81954
rect 31218 81902 31220 81954
rect 30716 81900 31220 81902
rect 30716 81842 30772 81900
rect 31164 81890 31220 81900
rect 30716 81790 30718 81842
rect 30770 81790 30772 81842
rect 30716 81778 30772 81790
rect 31276 81732 31332 81742
rect 31276 81638 31332 81676
rect 31388 81508 31444 82236
rect 30940 81452 31444 81508
rect 30716 81172 30772 81182
rect 30604 81170 30772 81172
rect 30604 81118 30718 81170
rect 30770 81118 30772 81170
rect 30604 81116 30772 81118
rect 30492 81004 30660 81060
rect 30492 79268 30548 79278
rect 30380 79212 30492 79268
rect 30492 79202 30548 79212
rect 30044 78754 30100 78764
rect 30492 78930 30548 78942
rect 30492 78878 30494 78930
rect 30546 78878 30548 78930
rect 30492 78820 30548 78878
rect 30492 78754 30548 78764
rect 30604 78932 30660 81004
rect 30604 78818 30660 78876
rect 30604 78766 30606 78818
rect 30658 78766 30660 78818
rect 30604 78754 30660 78766
rect 30716 80386 30772 81116
rect 30716 80334 30718 80386
rect 30770 80334 30772 80386
rect 30716 79716 30772 80334
rect 30828 80276 30884 80286
rect 30940 80276 30996 81452
rect 31052 81284 31108 81294
rect 31500 81284 31556 82460
rect 31836 82516 31892 82526
rect 31948 82516 32004 84028
rect 33180 82628 33236 82638
rect 31836 82514 32004 82516
rect 31836 82462 31838 82514
rect 31890 82462 32004 82514
rect 31836 82460 32004 82462
rect 31836 82450 31892 82460
rect 31612 81396 31668 81406
rect 31612 81302 31668 81340
rect 31052 81282 31556 81284
rect 31052 81230 31054 81282
rect 31106 81230 31556 81282
rect 31052 81228 31556 81230
rect 31052 81218 31108 81228
rect 30828 80274 30996 80276
rect 30828 80222 30830 80274
rect 30882 80222 30996 80274
rect 30828 80220 30996 80222
rect 30828 80210 30884 80220
rect 31500 79716 31556 79726
rect 30716 79714 31556 79716
rect 30716 79662 31502 79714
rect 31554 79662 31556 79714
rect 30716 79660 31556 79662
rect 30156 78596 30212 78606
rect 30156 78258 30212 78540
rect 30492 78596 30548 78634
rect 30492 78530 30548 78540
rect 30716 78372 30772 79660
rect 31500 79650 31556 79660
rect 31948 79714 32004 82460
rect 32284 82514 32340 82526
rect 32284 82462 32286 82514
rect 32338 82462 32340 82514
rect 32172 81844 32228 81854
rect 32284 81844 32340 82462
rect 32956 81956 33012 81966
rect 32956 81862 33012 81900
rect 32172 81842 32340 81844
rect 32172 81790 32174 81842
rect 32226 81790 32340 81842
rect 32172 81788 32340 81790
rect 32172 81778 32228 81788
rect 33180 81732 33236 82572
rect 33852 82404 33908 84142
rect 34524 84084 34580 84814
rect 34524 84018 34580 84028
rect 34636 84866 34804 84868
rect 34636 84814 34750 84866
rect 34802 84814 34804 84866
rect 34636 84812 34804 84814
rect 34636 83860 34692 84812
rect 34748 84802 34804 84812
rect 34972 84978 35028 84990
rect 34972 84926 34974 84978
rect 35026 84926 35028 84978
rect 34972 84868 35028 84926
rect 35308 84978 35364 84990
rect 35308 84926 35310 84978
rect 35362 84926 35364 84978
rect 34972 84802 35028 84812
rect 35084 84866 35140 84878
rect 35084 84814 35086 84866
rect 35138 84814 35140 84866
rect 34524 83804 34692 83860
rect 34748 84532 34804 84542
rect 34076 83300 34132 83310
rect 34412 83300 34468 83310
rect 34076 83298 34468 83300
rect 34076 83246 34078 83298
rect 34130 83246 34414 83298
rect 34466 83246 34468 83298
rect 34076 83244 34468 83246
rect 34076 83234 34132 83244
rect 33852 82338 33908 82348
rect 31948 79662 31950 79714
rect 32002 79662 32004 79714
rect 31948 79650 32004 79662
rect 32956 81676 33236 81732
rect 34188 81956 34244 81966
rect 34188 81730 34244 81900
rect 34188 81678 34190 81730
rect 34242 81678 34244 81730
rect 30940 79380 30996 79390
rect 30940 79286 30996 79324
rect 31276 79380 31332 79390
rect 31276 79378 31668 79380
rect 31276 79326 31278 79378
rect 31330 79326 31668 79378
rect 31276 79324 31668 79326
rect 31276 79314 31332 79324
rect 31276 78988 31556 79044
rect 31052 78820 31108 78830
rect 31276 78820 31332 78988
rect 31500 78930 31556 78988
rect 31500 78878 31502 78930
rect 31554 78878 31556 78930
rect 31500 78866 31556 78878
rect 31052 78818 31332 78820
rect 31052 78766 31054 78818
rect 31106 78766 31332 78818
rect 31052 78764 31332 78766
rect 31388 78818 31444 78830
rect 31388 78766 31390 78818
rect 31442 78766 31444 78818
rect 31052 78754 31108 78764
rect 31388 78708 31444 78766
rect 31500 78708 31556 78718
rect 31388 78652 31500 78708
rect 31500 78642 31556 78652
rect 30828 78596 30884 78606
rect 30828 78594 31108 78596
rect 30828 78542 30830 78594
rect 30882 78542 31108 78594
rect 30828 78540 31108 78542
rect 30828 78530 30884 78540
rect 30156 78206 30158 78258
rect 30210 78206 30212 78258
rect 30156 78194 30212 78206
rect 30604 78316 30772 78372
rect 30268 78034 30324 78046
rect 30268 77982 30270 78034
rect 30322 77982 30324 78034
rect 30156 77924 30212 77934
rect 29932 77922 30212 77924
rect 29932 77870 30158 77922
rect 30210 77870 30212 77922
rect 29932 77868 30212 77870
rect 30156 77858 30212 77868
rect 30268 77700 30324 77982
rect 30268 77026 30324 77644
rect 30268 76974 30270 77026
rect 30322 76974 30324 77026
rect 30268 76916 30324 76974
rect 30380 78036 30436 78046
rect 30380 77028 30436 77980
rect 30380 76962 30436 76972
rect 30492 78034 30548 78046
rect 30492 77982 30494 78034
rect 30546 77982 30548 78034
rect 30156 76860 30324 76916
rect 30156 76804 30212 76860
rect 30492 76804 30548 77982
rect 30604 77812 30660 78316
rect 30716 78036 30772 78046
rect 30716 78034 30996 78036
rect 30716 77982 30718 78034
rect 30770 77982 30996 78034
rect 30716 77980 30996 77982
rect 30716 77970 30772 77980
rect 30828 77812 30884 77822
rect 30604 77756 30772 77812
rect 30156 76738 30212 76748
rect 30268 76748 30548 76804
rect 30604 77026 30660 77038
rect 30604 76974 30606 77026
rect 30658 76974 30660 77026
rect 29932 76244 29988 76254
rect 29932 76242 30100 76244
rect 29932 76190 29934 76242
rect 29986 76190 30100 76242
rect 29932 76188 30100 76190
rect 29932 76178 29988 76188
rect 29820 75964 29988 76020
rect 29708 74286 29710 74338
rect 29762 74286 29764 74338
rect 29708 74274 29764 74286
rect 29820 75572 29876 75582
rect 29820 74228 29876 75516
rect 29820 74134 29876 74172
rect 29820 73444 29876 73454
rect 29820 73350 29876 73388
rect 29596 73278 29598 73330
rect 29650 73278 29652 73330
rect 29596 71876 29652 73278
rect 29708 73218 29764 73230
rect 29708 73166 29710 73218
rect 29762 73166 29764 73218
rect 29708 71988 29764 73166
rect 29820 72660 29876 72670
rect 29820 72566 29876 72604
rect 29708 71932 29876 71988
rect 29596 71820 29764 71876
rect 29372 71474 29428 71484
rect 29260 71148 29652 71204
rect 29372 70980 29428 70990
rect 29428 70924 29540 70980
rect 29372 70886 29428 70924
rect 29148 70354 29204 70364
rect 28924 70254 28926 70306
rect 28978 70254 28980 70306
rect 28924 70242 28980 70254
rect 28588 70140 28868 70196
rect 29148 70194 29204 70206
rect 29148 70142 29150 70194
rect 29202 70142 29204 70194
rect 28476 70084 28532 70094
rect 28364 70082 28532 70084
rect 28364 70030 28478 70082
rect 28530 70030 28532 70082
rect 28364 70028 28532 70030
rect 28476 69972 28532 70028
rect 28476 69906 28532 69916
rect 28364 69636 28420 69646
rect 28364 69522 28420 69580
rect 28364 69470 28366 69522
rect 28418 69470 28420 69522
rect 28364 69458 28420 69470
rect 28588 69524 28644 70140
rect 28700 69970 28756 69982
rect 28700 69918 28702 69970
rect 28754 69918 28756 69970
rect 28700 69636 28756 69918
rect 29148 69748 29204 70142
rect 29484 70082 29540 70924
rect 29484 70030 29486 70082
rect 29538 70030 29540 70082
rect 29484 70018 29540 70030
rect 29260 69748 29316 69758
rect 29148 69692 29260 69748
rect 29260 69682 29316 69692
rect 29596 69636 29652 71148
rect 29708 70196 29764 71820
rect 29820 70644 29876 71932
rect 29932 71874 29988 75964
rect 30044 75794 30100 76188
rect 30044 75742 30046 75794
rect 30098 75742 30100 75794
rect 30044 75730 30100 75742
rect 30156 75796 30212 75806
rect 30156 75682 30212 75740
rect 30156 75630 30158 75682
rect 30210 75630 30212 75682
rect 30156 75618 30212 75630
rect 30044 75460 30100 75470
rect 30044 75366 30100 75404
rect 29932 71822 29934 71874
rect 29986 71822 29988 71874
rect 29932 71810 29988 71822
rect 30156 74898 30212 74910
rect 30156 74846 30158 74898
rect 30210 74846 30212 74898
rect 30156 74338 30212 74846
rect 30268 74452 30324 76748
rect 30492 76580 30548 76590
rect 30492 76486 30548 76524
rect 30380 76466 30436 76478
rect 30380 76414 30382 76466
rect 30434 76414 30436 76466
rect 30380 76244 30436 76414
rect 30604 76244 30660 76974
rect 30380 76178 30436 76188
rect 30492 76188 30660 76244
rect 30716 76244 30772 77756
rect 30828 76244 30884 77756
rect 30940 77476 30996 77980
rect 31052 77588 31108 78540
rect 31388 78260 31444 78270
rect 31612 78260 31668 79324
rect 32396 78932 32452 78942
rect 32396 78838 32452 78876
rect 31836 78818 31892 78830
rect 31836 78766 31838 78818
rect 31890 78766 31892 78818
rect 31724 78706 31780 78718
rect 31724 78654 31726 78706
rect 31778 78654 31780 78706
rect 31724 78372 31780 78654
rect 31724 78306 31780 78316
rect 31836 78596 31892 78766
rect 31388 78258 31668 78260
rect 31388 78206 31390 78258
rect 31442 78206 31668 78258
rect 31388 78204 31668 78206
rect 31388 78194 31444 78204
rect 31164 78034 31220 78046
rect 31164 77982 31166 78034
rect 31218 77982 31220 78034
rect 31164 77588 31220 77982
rect 31276 78036 31332 78046
rect 31276 77942 31332 77980
rect 31500 78036 31556 78046
rect 31500 77942 31556 77980
rect 31724 78036 31780 78046
rect 31836 78036 31892 78540
rect 31724 78034 31892 78036
rect 31724 77982 31726 78034
rect 31778 77982 31892 78034
rect 31724 77980 31892 77982
rect 32060 78708 32116 78718
rect 31612 77588 31668 77598
rect 31164 77532 31444 77588
rect 31052 77522 31108 77532
rect 30940 77410 30996 77420
rect 31164 77364 31220 77374
rect 31220 77308 31332 77364
rect 31164 77298 31220 77308
rect 31276 77250 31332 77308
rect 31276 77198 31278 77250
rect 31330 77198 31332 77250
rect 31276 77186 31332 77198
rect 31164 77138 31220 77150
rect 31164 77086 31166 77138
rect 31218 77086 31220 77138
rect 31164 76916 31220 77086
rect 31164 76578 31220 76860
rect 31164 76526 31166 76578
rect 31218 76526 31220 76578
rect 31164 76514 31220 76526
rect 31276 77028 31332 77038
rect 30828 76188 31220 76244
rect 30380 75796 30436 75806
rect 30492 75796 30548 76188
rect 30716 76178 30772 76188
rect 30436 75740 30548 75796
rect 31052 76020 31108 76030
rect 31052 75794 31108 75964
rect 31052 75742 31054 75794
rect 31106 75742 31108 75794
rect 30380 75730 30436 75740
rect 31052 75730 31108 75742
rect 30604 75684 30660 75694
rect 30604 75590 30660 75628
rect 30940 75572 30996 75582
rect 30940 75478 30996 75516
rect 30380 75460 30436 75470
rect 31164 75460 31220 76188
rect 31276 75682 31332 76972
rect 31388 76690 31444 77532
rect 31500 77140 31556 77150
rect 31500 77046 31556 77084
rect 31388 76638 31390 76690
rect 31442 76638 31444 76690
rect 31388 76626 31444 76638
rect 31500 76580 31556 76590
rect 31612 76580 31668 77532
rect 31500 76578 31668 76580
rect 31500 76526 31502 76578
rect 31554 76526 31668 76578
rect 31500 76524 31668 76526
rect 31724 77138 31780 77980
rect 31724 77086 31726 77138
rect 31778 77086 31780 77138
rect 31724 76804 31780 77086
rect 31500 76514 31556 76524
rect 31724 76468 31780 76748
rect 32060 77476 32116 78652
rect 32732 78596 32788 78606
rect 32396 78372 32452 78382
rect 32172 78260 32228 78270
rect 32172 78166 32228 78204
rect 32060 77250 32116 77420
rect 32396 77364 32452 78316
rect 32396 77298 32452 77308
rect 32060 77198 32062 77250
rect 32114 77198 32116 77250
rect 32060 76916 32116 77198
rect 32172 77252 32228 77262
rect 32172 77158 32228 77196
rect 32508 77250 32564 77262
rect 32508 77198 32510 77250
rect 32562 77198 32564 77250
rect 32060 76692 32116 76860
rect 32396 77138 32452 77150
rect 32396 77086 32398 77138
rect 32450 77086 32452 77138
rect 32396 76916 32452 77086
rect 32396 76850 32452 76860
rect 32508 76804 32564 77198
rect 32508 76738 32564 76748
rect 31276 75630 31278 75682
rect 31330 75630 31332 75682
rect 31276 75618 31332 75630
rect 31612 76466 31780 76468
rect 31612 76414 31726 76466
rect 31778 76414 31780 76466
rect 31612 76412 31780 76414
rect 31500 75572 31556 75582
rect 31612 75572 31668 76412
rect 31724 76402 31780 76412
rect 31836 76636 32116 76692
rect 31836 75682 31892 76636
rect 32396 76580 32452 76590
rect 32620 76580 32676 76590
rect 32732 76580 32788 78540
rect 32844 78594 32900 78606
rect 32844 78542 32846 78594
rect 32898 78542 32900 78594
rect 32844 78036 32900 78542
rect 32844 77970 32900 77980
rect 32396 76578 32564 76580
rect 32396 76526 32398 76578
rect 32450 76526 32564 76578
rect 32396 76524 32564 76526
rect 32396 76514 32452 76524
rect 32284 76466 32340 76478
rect 32284 76414 32286 76466
rect 32338 76414 32340 76466
rect 32284 75796 32340 76414
rect 32508 75906 32564 76524
rect 32620 76578 32788 76580
rect 32620 76526 32622 76578
rect 32674 76526 32788 76578
rect 32620 76524 32788 76526
rect 32956 76580 33012 81676
rect 34188 80724 34244 81678
rect 34412 81732 34468 83244
rect 34524 82628 34580 83804
rect 34748 83634 34804 84476
rect 34972 84532 35028 84542
rect 35084 84532 35140 84814
rect 34972 84530 35140 84532
rect 34972 84478 34974 84530
rect 35026 84478 35140 84530
rect 34972 84476 35140 84478
rect 35308 84532 35364 84926
rect 35420 84866 35476 84878
rect 35420 84814 35422 84866
rect 35474 84814 35476 84866
rect 35420 84756 35476 84814
rect 35420 84690 35476 84700
rect 34972 84466 35028 84476
rect 35308 84466 35364 84476
rect 35308 84308 35364 84318
rect 35532 84308 35588 86604
rect 35644 86594 35700 86604
rect 35756 85762 35812 88060
rect 36204 88004 36260 88014
rect 36204 86772 36260 87948
rect 36204 86770 36372 86772
rect 36204 86718 36206 86770
rect 36258 86718 36372 86770
rect 36204 86716 36372 86718
rect 36204 86706 36260 86716
rect 36316 86100 36372 86716
rect 36316 86098 36484 86100
rect 36316 86046 36318 86098
rect 36370 86046 36484 86098
rect 36316 86044 36484 86046
rect 36316 86034 36372 86044
rect 36204 85876 36260 85886
rect 35756 85710 35758 85762
rect 35810 85710 35812 85762
rect 35756 85698 35812 85710
rect 35868 85874 36260 85876
rect 35868 85822 36206 85874
rect 36258 85822 36260 85874
rect 35868 85820 36260 85822
rect 35868 85428 35924 85820
rect 36204 85810 36260 85820
rect 35644 85372 35924 85428
rect 36316 85650 36372 85662
rect 36316 85598 36318 85650
rect 36370 85598 36372 85650
rect 35644 85090 35700 85372
rect 35980 85204 36036 85214
rect 35644 85038 35646 85090
rect 35698 85038 35700 85090
rect 35644 85026 35700 85038
rect 35868 85092 35924 85102
rect 35868 84998 35924 85036
rect 35980 84978 36036 85148
rect 35980 84926 35982 84978
rect 36034 84926 36036 84978
rect 35980 84914 36036 84926
rect 36204 84868 36260 84878
rect 36092 84866 36260 84868
rect 36092 84814 36206 84866
rect 36258 84814 36260 84866
rect 36092 84812 36260 84814
rect 36092 84420 36148 84812
rect 36204 84802 36260 84812
rect 34748 83582 34750 83634
rect 34802 83582 34804 83634
rect 34748 83570 34804 83582
rect 35084 84306 35588 84308
rect 35084 84254 35310 84306
rect 35362 84254 35588 84306
rect 35084 84252 35588 84254
rect 35980 84364 36148 84420
rect 34860 83524 34916 83534
rect 34860 83430 34916 83468
rect 34636 83300 34692 83310
rect 34636 83206 34692 83244
rect 34972 82740 35028 82750
rect 35084 82740 35140 84252
rect 35308 84242 35364 84252
rect 35644 83972 35700 83982
rect 35196 83916 35460 83926
rect 35252 83860 35300 83916
rect 35356 83860 35404 83916
rect 35196 83850 35460 83860
rect 35644 83522 35700 83916
rect 35644 83470 35646 83522
rect 35698 83470 35700 83522
rect 35644 83458 35700 83470
rect 35980 83524 36036 84364
rect 36092 84194 36148 84206
rect 36092 84142 36094 84194
rect 36146 84142 36148 84194
rect 36092 83748 36148 84142
rect 36092 83682 36148 83692
rect 35980 83430 36036 83468
rect 36204 83412 36260 83422
rect 36204 83318 36260 83356
rect 35756 82852 35812 82862
rect 36316 82852 36372 85598
rect 36428 84532 36484 86044
rect 36540 84644 36596 88846
rect 37772 87332 37828 87342
rect 37324 87330 37828 87332
rect 37324 87278 37774 87330
rect 37826 87278 37828 87330
rect 37324 87276 37828 87278
rect 36876 85764 36932 85774
rect 37324 85764 37380 87276
rect 37772 87266 37828 87276
rect 36876 85762 37380 85764
rect 36876 85710 36878 85762
rect 36930 85710 37326 85762
rect 37378 85710 37380 85762
rect 36876 85708 37380 85710
rect 36876 85204 36932 85708
rect 37324 85698 37380 85708
rect 37100 85204 37156 85214
rect 36932 85202 37156 85204
rect 36932 85150 37102 85202
rect 37154 85150 37156 85202
rect 36932 85148 37156 85150
rect 36876 85138 36932 85148
rect 37100 85138 37156 85148
rect 38332 84980 38388 99600
rect 38332 84914 38388 84924
rect 37660 84868 37716 84878
rect 37716 84812 37828 84868
rect 37660 84774 37716 84812
rect 36540 84578 36596 84588
rect 36428 84466 36484 84476
rect 37100 84532 37156 84542
rect 37156 84476 37268 84532
rect 37100 84466 37156 84476
rect 37212 84084 37268 84476
rect 37100 83748 37156 83758
rect 37100 83654 37156 83692
rect 36988 83412 37044 83422
rect 36988 83318 37044 83356
rect 37100 83412 37156 83422
rect 37212 83412 37268 84028
rect 37660 83972 37716 83982
rect 37660 83634 37716 83916
rect 37660 83582 37662 83634
rect 37714 83582 37716 83634
rect 37660 83570 37716 83582
rect 37100 83410 37268 83412
rect 37100 83358 37102 83410
rect 37154 83358 37268 83410
rect 37100 83356 37268 83358
rect 37100 83346 37156 83356
rect 37548 83300 37604 83310
rect 37548 83206 37604 83244
rect 35756 82850 36372 82852
rect 35756 82798 35758 82850
rect 35810 82798 36372 82850
rect 35756 82796 36372 82798
rect 35756 82786 35812 82796
rect 34972 82738 35140 82740
rect 34972 82686 34974 82738
rect 35026 82686 35140 82738
rect 34972 82684 35140 82686
rect 34524 82562 34580 82572
rect 34636 82628 34692 82638
rect 34972 82628 35028 82684
rect 34636 82626 35028 82628
rect 34636 82574 34638 82626
rect 34690 82574 35028 82626
rect 34636 82572 35028 82574
rect 37772 82628 37828 84812
rect 38220 84194 38276 84206
rect 38220 84142 38222 84194
rect 38274 84142 38276 84194
rect 38108 84084 38164 84094
rect 38108 83634 38164 84028
rect 38220 83972 38276 84142
rect 38220 83906 38276 83916
rect 38108 83582 38110 83634
rect 38162 83582 38164 83634
rect 38108 83570 38164 83582
rect 37884 82628 37940 82638
rect 37772 82626 37940 82628
rect 37772 82574 37886 82626
rect 37938 82574 37940 82626
rect 37772 82572 37940 82574
rect 34636 82404 34692 82572
rect 34636 82338 34692 82348
rect 35196 82348 35460 82358
rect 35252 82292 35300 82348
rect 35356 82292 35404 82348
rect 35196 82282 35460 82292
rect 35196 81956 35252 81966
rect 35196 81862 35252 81900
rect 36204 81956 36260 81966
rect 36204 81862 36260 81900
rect 37884 81956 37940 82572
rect 37884 81890 37940 81900
rect 34412 81666 34468 81676
rect 35308 81732 35364 81742
rect 35308 81638 35364 81676
rect 35196 80780 35460 80790
rect 35252 80724 35300 80780
rect 35356 80724 35404 80780
rect 35196 80714 35460 80724
rect 34188 80658 34244 80668
rect 33292 79492 33348 79502
rect 33292 79490 33572 79492
rect 33292 79438 33294 79490
rect 33346 79438 33572 79490
rect 33292 79436 33572 79438
rect 33292 79426 33348 79436
rect 33292 78932 33348 78942
rect 33516 78932 33572 79436
rect 35196 79212 35460 79222
rect 35252 79156 35300 79212
rect 35356 79156 35404 79212
rect 35196 79146 35460 79156
rect 33740 78932 33796 78942
rect 33516 78930 33796 78932
rect 33516 78878 33742 78930
rect 33794 78878 33796 78930
rect 33516 78876 33796 78878
rect 33292 78838 33348 78876
rect 33628 78260 33684 78876
rect 33740 78866 33796 78876
rect 34972 78706 35028 78718
rect 34972 78654 34974 78706
rect 35026 78654 35028 78706
rect 34636 78596 34692 78606
rect 33068 78258 33684 78260
rect 33068 78206 33630 78258
rect 33682 78206 33684 78258
rect 33068 78204 33684 78206
rect 33068 77476 33124 78204
rect 33628 78194 33684 78204
rect 34524 78594 34692 78596
rect 34524 78542 34638 78594
rect 34690 78542 34692 78594
rect 34524 78540 34692 78542
rect 34412 78036 34468 78046
rect 33180 77922 33236 77934
rect 33180 77870 33182 77922
rect 33234 77870 33236 77922
rect 33180 77700 33236 77870
rect 34076 77924 34132 77934
rect 34076 77830 34132 77868
rect 33180 77634 33236 77644
rect 34412 77810 34468 77980
rect 34412 77758 34414 77810
rect 34466 77758 34468 77810
rect 33068 77250 33124 77420
rect 33068 77198 33070 77250
rect 33122 77198 33124 77250
rect 33068 77186 33124 77198
rect 34412 77252 34468 77758
rect 34524 77588 34580 78540
rect 34636 78530 34692 78540
rect 34860 78596 34916 78606
rect 34860 78502 34916 78540
rect 34972 78260 35028 78654
rect 35644 78594 35700 78606
rect 35644 78542 35646 78594
rect 35698 78542 35700 78594
rect 35196 78260 35252 78270
rect 34972 78258 35252 78260
rect 34972 78206 35198 78258
rect 35250 78206 35252 78258
rect 34972 78204 35252 78206
rect 35196 78194 35252 78204
rect 35308 78260 35364 78270
rect 35308 78166 35364 78204
rect 34636 78148 34692 78158
rect 34636 78054 34692 78092
rect 35084 78036 35140 78074
rect 35084 77970 35140 77980
rect 35532 78036 35588 78046
rect 35532 77942 35588 77980
rect 34748 77812 34804 77822
rect 35084 77812 35140 77822
rect 34748 77810 35084 77812
rect 34748 77758 34750 77810
rect 34802 77758 35084 77810
rect 34748 77756 35084 77758
rect 34748 77746 34804 77756
rect 34524 77522 34580 77532
rect 33292 77140 33348 77150
rect 33292 77046 33348 77084
rect 33628 77138 33684 77150
rect 33628 77086 33630 77138
rect 33682 77086 33684 77138
rect 33516 77026 33572 77038
rect 33516 76974 33518 77026
rect 33570 76974 33572 77026
rect 33180 76916 33236 76926
rect 33236 76860 33460 76916
rect 33180 76850 33236 76860
rect 33404 76690 33460 76860
rect 33404 76638 33406 76690
rect 33458 76638 33460 76690
rect 33404 76626 33460 76638
rect 33516 76692 33572 76974
rect 33628 76916 33684 77086
rect 34188 77140 34244 77150
rect 34188 77046 34244 77084
rect 34300 77028 34356 77038
rect 34300 76934 34356 76972
rect 33628 76850 33684 76860
rect 33516 76636 33684 76692
rect 32620 76514 32676 76524
rect 32508 75854 32510 75906
rect 32562 75854 32564 75906
rect 32508 75842 32564 75854
rect 32284 75730 32340 75740
rect 32956 75794 33012 76524
rect 32956 75742 32958 75794
rect 33010 75742 33012 75794
rect 32956 75730 33012 75742
rect 33292 76466 33348 76478
rect 33292 76414 33294 76466
rect 33346 76414 33348 76466
rect 33292 75906 33348 76414
rect 33516 76468 33572 76478
rect 33516 76374 33572 76412
rect 33292 75854 33294 75906
rect 33346 75854 33348 75906
rect 31836 75630 31838 75682
rect 31890 75630 31892 75682
rect 31836 75572 31892 75630
rect 31948 75684 32004 75694
rect 31948 75590 32004 75628
rect 31500 75570 31668 75572
rect 31500 75518 31502 75570
rect 31554 75518 31668 75570
rect 31500 75516 31668 75518
rect 31500 75506 31556 75516
rect 31612 75460 31668 75516
rect 30380 75458 30884 75460
rect 30380 75406 30382 75458
rect 30434 75406 30884 75458
rect 30380 75404 30884 75406
rect 31164 75404 31332 75460
rect 30380 75394 30436 75404
rect 30492 75236 30548 75246
rect 30492 74898 30548 75180
rect 30492 74846 30494 74898
rect 30546 74846 30548 74898
rect 30492 74834 30548 74846
rect 30604 74900 30660 74910
rect 30604 74806 30660 74844
rect 30268 74396 30436 74452
rect 30156 74286 30158 74338
rect 30210 74286 30212 74338
rect 30156 73330 30212 74286
rect 30268 74228 30324 74238
rect 30268 74134 30324 74172
rect 30156 73278 30158 73330
rect 30210 73278 30212 73330
rect 29820 70578 29876 70588
rect 29932 71092 29988 71102
rect 29708 70130 29764 70140
rect 29708 69972 29764 69982
rect 29708 69970 29876 69972
rect 29708 69918 29710 69970
rect 29762 69918 29876 69970
rect 29708 69916 29876 69918
rect 29708 69906 29764 69916
rect 28700 69580 28980 69636
rect 28588 69468 28756 69524
rect 28308 69244 28532 69300
rect 28252 69234 28308 69244
rect 28252 68852 28308 68862
rect 28140 68850 28308 68852
rect 28140 68798 28254 68850
rect 28306 68798 28308 68850
rect 28140 68796 28308 68798
rect 28252 68786 28308 68796
rect 28476 68850 28532 69244
rect 28476 68798 28478 68850
rect 28530 68798 28532 68850
rect 28476 68516 28532 68798
rect 28476 68450 28532 68460
rect 28588 68626 28644 68638
rect 28588 68574 28590 68626
rect 28642 68574 28644 68626
rect 28588 67956 28644 68574
rect 28588 67890 28644 67900
rect 28700 66052 28756 69468
rect 28924 67396 28980 69580
rect 29372 69524 29428 69534
rect 29148 69412 29204 69422
rect 29148 69318 29204 69356
rect 29372 69186 29428 69468
rect 29596 69410 29652 69580
rect 29596 69358 29598 69410
rect 29650 69358 29652 69410
rect 29596 69346 29652 69358
rect 29372 69134 29374 69186
rect 29426 69134 29428 69186
rect 29372 69122 29428 69134
rect 29484 69298 29540 69310
rect 29484 69246 29486 69298
rect 29538 69246 29540 69298
rect 29484 69188 29540 69246
rect 29484 69132 29652 69188
rect 29036 68516 29092 68526
rect 29036 68422 29092 68460
rect 29260 68516 29316 68526
rect 29372 68516 29428 68526
rect 29484 68516 29540 68526
rect 29316 68514 29540 68516
rect 29316 68462 29374 68514
rect 29426 68462 29486 68514
rect 29538 68462 29540 68514
rect 29316 68460 29540 68462
rect 29596 68516 29652 69132
rect 29708 68516 29764 68526
rect 29596 68460 29708 68516
rect 29260 68450 29316 68460
rect 29372 68422 29428 68460
rect 29484 68450 29540 68460
rect 29708 68450 29764 68460
rect 29596 68292 29652 68302
rect 29596 67954 29652 68236
rect 29596 67902 29598 67954
rect 29650 67902 29652 67954
rect 28924 67340 29092 67396
rect 29036 67284 29092 67340
rect 29036 67228 29316 67284
rect 29260 67170 29316 67228
rect 29260 67118 29262 67170
rect 29314 67118 29316 67170
rect 29260 67106 29316 67118
rect 29596 67172 29652 67902
rect 29148 67060 29204 67070
rect 29148 66966 29204 67004
rect 29484 67058 29540 67070
rect 29484 67006 29486 67058
rect 29538 67006 29540 67058
rect 29484 66836 29540 67006
rect 29484 66770 29540 66780
rect 29596 66612 29652 67116
rect 29260 66556 29652 66612
rect 29708 68180 29764 68190
rect 29260 66498 29316 66556
rect 29260 66446 29262 66498
rect 29314 66446 29316 66498
rect 29260 66434 29316 66446
rect 29708 66386 29764 68124
rect 29820 67956 29876 69916
rect 29932 69748 29988 71036
rect 30156 71090 30212 73278
rect 30156 71038 30158 71090
rect 30210 71038 30212 71090
rect 30156 71026 30212 71038
rect 30268 71540 30324 71550
rect 30268 70868 30324 71484
rect 30268 70802 30324 70812
rect 30380 70644 30436 74396
rect 30716 74228 30772 74238
rect 30716 74134 30772 74172
rect 30492 73556 30548 73566
rect 30492 73462 30548 73500
rect 30604 73220 30660 73230
rect 30380 70578 30436 70588
rect 30492 73218 30660 73220
rect 30492 73166 30606 73218
rect 30658 73166 30660 73218
rect 30492 73164 30660 73166
rect 30380 70194 30436 70206
rect 30380 70142 30382 70194
rect 30434 70142 30436 70194
rect 30044 69972 30100 69982
rect 30044 69970 30324 69972
rect 30044 69918 30046 69970
rect 30098 69918 30324 69970
rect 30044 69916 30324 69918
rect 30044 69906 30100 69916
rect 29932 69692 30212 69748
rect 30044 68740 30100 68750
rect 29820 67890 29876 67900
rect 29932 68684 30044 68740
rect 29932 66500 29988 68684
rect 30044 68674 30100 68684
rect 30044 68516 30100 68526
rect 30156 68516 30212 69692
rect 30268 69410 30324 69916
rect 30268 69358 30270 69410
rect 30322 69358 30324 69410
rect 30268 69346 30324 69358
rect 30100 68460 30212 68516
rect 30380 68964 30436 70142
rect 30492 69524 30548 73164
rect 30604 73154 30660 73164
rect 30604 70980 30660 70990
rect 30604 70306 30660 70924
rect 30716 70868 30772 70878
rect 30828 70868 30884 75404
rect 31276 73948 31332 75404
rect 31500 74228 31556 74238
rect 31500 74004 31556 74172
rect 31276 73892 31444 73948
rect 31052 73444 31108 73454
rect 31052 73350 31108 73388
rect 31276 72548 31332 72558
rect 31276 72454 31332 72492
rect 31388 70980 31444 73892
rect 31500 73554 31556 73948
rect 31500 73502 31502 73554
rect 31554 73502 31556 73554
rect 31500 73490 31556 73502
rect 31276 70924 31444 70980
rect 31052 70868 31108 70906
rect 30828 70812 30996 70868
rect 30716 70588 30772 70812
rect 30716 70532 30884 70588
rect 30604 70254 30606 70306
rect 30658 70254 30660 70306
rect 30604 70242 30660 70254
rect 30828 70306 30884 70532
rect 30828 70254 30830 70306
rect 30882 70254 30884 70306
rect 30828 70242 30884 70254
rect 30492 69458 30548 69468
rect 30716 70196 30772 70206
rect 30380 68514 30436 68908
rect 30716 68852 30772 70140
rect 30940 70084 30996 70812
rect 31052 70802 31108 70812
rect 30380 68462 30382 68514
rect 30434 68462 30436 68514
rect 30044 68422 30100 68460
rect 30380 68402 30436 68462
rect 30380 68350 30382 68402
rect 30434 68350 30436 68402
rect 30380 68338 30436 68350
rect 30604 68796 30772 68852
rect 30828 70028 30996 70084
rect 31052 70644 31108 70654
rect 30380 67730 30436 67742
rect 30380 67678 30382 67730
rect 30434 67678 30436 67730
rect 30044 66948 30100 66958
rect 30100 66892 30324 66948
rect 30044 66854 30100 66892
rect 30044 66500 30100 66510
rect 29932 66498 30100 66500
rect 29932 66446 30046 66498
rect 30098 66446 30100 66498
rect 29932 66444 30100 66446
rect 30044 66434 30100 66444
rect 29708 66334 29710 66386
rect 29762 66334 29764 66386
rect 29708 66322 29764 66334
rect 29484 66274 29540 66286
rect 29484 66222 29486 66274
rect 29538 66222 29540 66274
rect 28812 66052 28868 66062
rect 28700 65996 28812 66052
rect 28812 65986 28868 65996
rect 28812 65492 28868 65502
rect 28700 65490 28868 65492
rect 28700 65438 28814 65490
rect 28866 65438 28868 65490
rect 28700 65436 28868 65438
rect 28588 65380 28644 65390
rect 28700 65380 28756 65436
rect 28812 65426 28868 65436
rect 28588 65378 28756 65380
rect 28588 65326 28590 65378
rect 28642 65326 28756 65378
rect 28588 65324 28756 65326
rect 28588 65314 28644 65324
rect 28588 64932 28644 64942
rect 28588 64838 28644 64876
rect 28028 64766 28030 64818
rect 28082 64766 28084 64818
rect 28028 64754 28084 64766
rect 28252 64708 28308 64718
rect 28140 64706 28308 64708
rect 28140 64654 28254 64706
rect 28306 64654 28308 64706
rect 28140 64652 28308 64654
rect 27804 64596 27860 64606
rect 27804 64502 27860 64540
rect 28140 64148 28196 64652
rect 28252 64642 28308 64652
rect 28700 64148 28756 65324
rect 29484 64932 29540 66222
rect 30268 66276 30324 66892
rect 30380 66498 30436 67678
rect 30604 67284 30660 68796
rect 30716 68628 30772 68638
rect 30716 67730 30772 68572
rect 30716 67678 30718 67730
rect 30770 67678 30772 67730
rect 30716 67666 30772 67678
rect 30604 67228 30772 67284
rect 30492 67172 30548 67182
rect 30492 67078 30548 67116
rect 30380 66446 30382 66498
rect 30434 66446 30436 66498
rect 30380 66434 30436 66446
rect 30716 66388 30772 67228
rect 30492 66332 30772 66388
rect 30380 66276 30436 66286
rect 30268 66274 30436 66276
rect 30268 66222 30382 66274
rect 30434 66222 30436 66274
rect 30268 66220 30436 66222
rect 30380 66210 30436 66220
rect 29820 66162 29876 66174
rect 29820 66110 29822 66162
rect 29874 66110 29876 66162
rect 29708 66052 29764 66062
rect 29484 64866 29540 64876
rect 29596 65492 29652 65502
rect 29596 64930 29652 65436
rect 29596 64878 29598 64930
rect 29650 64878 29652 64930
rect 29596 64866 29652 64878
rect 29260 64596 29316 64606
rect 29260 64502 29316 64540
rect 29484 64484 29540 64494
rect 28140 64082 28196 64092
rect 28476 64146 28756 64148
rect 28476 64094 28702 64146
rect 28754 64094 28756 64146
rect 28476 64092 28756 64094
rect 27132 64036 27188 64046
rect 27132 63942 27188 63980
rect 27804 64036 27860 64046
rect 27804 63924 27860 63980
rect 27692 63922 27860 63924
rect 27692 63870 27806 63922
rect 27858 63870 27860 63922
rect 27692 63868 27860 63870
rect 27356 63812 27412 63822
rect 27356 63250 27412 63756
rect 27356 63198 27358 63250
rect 27410 63198 27412 63250
rect 27356 63186 27412 63198
rect 27020 63074 27076 63084
rect 26684 62514 26740 62524
rect 25676 62302 25678 62354
rect 25730 62302 25732 62354
rect 25676 62290 25732 62302
rect 25900 62466 25956 62478
rect 25900 62414 25902 62466
rect 25954 62414 25956 62466
rect 25900 62188 25956 62414
rect 25900 62132 26628 62188
rect 26572 61682 26628 62132
rect 27580 61796 27636 61806
rect 26572 61630 26574 61682
rect 26626 61630 26628 61682
rect 26572 61618 26628 61630
rect 27356 61794 27636 61796
rect 27356 61742 27582 61794
rect 27634 61742 27636 61794
rect 27356 61740 27636 61742
rect 27356 61570 27412 61740
rect 27580 61730 27636 61740
rect 27356 61518 27358 61570
rect 27410 61518 27412 61570
rect 27356 61506 27412 61518
rect 25340 61012 25396 61022
rect 25228 61010 25396 61012
rect 25228 60958 25342 61010
rect 25394 60958 25396 61010
rect 25228 60956 25396 60958
rect 25340 60946 25396 60956
rect 27692 61012 27748 63868
rect 27804 63858 27860 63868
rect 28252 63812 28308 63822
rect 28476 63812 28532 64092
rect 28700 64082 28756 64092
rect 28812 64148 28868 64158
rect 28252 63810 28532 63812
rect 28252 63758 28254 63810
rect 28306 63758 28532 63810
rect 28252 63756 28532 63758
rect 28588 63924 28644 63934
rect 28812 63924 28868 64092
rect 29148 64148 29204 64158
rect 29148 64034 29204 64092
rect 29484 64148 29540 64428
rect 29484 64082 29540 64092
rect 29148 63982 29150 64034
rect 29202 63982 29204 64034
rect 29148 63970 29204 63982
rect 29260 64036 29316 64046
rect 29708 64036 29764 65996
rect 29820 64148 29876 66110
rect 30380 66052 30436 66062
rect 30268 65996 30380 66052
rect 30044 65490 30100 65502
rect 30044 65438 30046 65490
rect 30098 65438 30100 65490
rect 30044 64484 30100 65438
rect 30044 64390 30100 64428
rect 29820 64092 30212 64148
rect 29708 63980 29876 64036
rect 29260 63942 29316 63980
rect 28588 63922 28868 63924
rect 28588 63870 28590 63922
rect 28642 63870 28868 63922
rect 28588 63868 28868 63870
rect 28924 63924 28980 63934
rect 28252 63700 28308 63756
rect 28252 63634 28308 63644
rect 25564 60788 25620 60798
rect 25340 60786 25620 60788
rect 25340 60734 25566 60786
rect 25618 60734 25620 60786
rect 25340 60732 25620 60734
rect 25004 60226 25060 60238
rect 25004 60174 25006 60226
rect 25058 60174 25060 60226
rect 24892 58436 24948 58446
rect 24892 57092 24948 58380
rect 24892 56866 24948 57036
rect 24892 56814 24894 56866
rect 24946 56814 24948 56866
rect 24892 56308 24948 56814
rect 24892 56242 24948 56252
rect 25004 55076 25060 60174
rect 25340 60226 25396 60732
rect 25564 60722 25620 60732
rect 27468 60788 27524 60798
rect 27468 60694 27524 60732
rect 25340 60174 25342 60226
rect 25394 60174 25396 60226
rect 25340 60162 25396 60174
rect 25676 60004 25732 60014
rect 25676 59910 25732 59948
rect 26012 60004 26068 60014
rect 25900 59890 25956 59902
rect 25900 59838 25902 59890
rect 25954 59838 25956 59890
rect 25900 59556 25956 59838
rect 25452 59500 25956 59556
rect 25452 59442 25508 59500
rect 25452 59390 25454 59442
rect 25506 59390 25508 59442
rect 25452 59378 25508 59390
rect 25676 59220 25732 59230
rect 25676 57092 25732 59164
rect 25676 57036 25844 57092
rect 25340 56980 25396 56990
rect 25340 56978 25732 56980
rect 25340 56926 25342 56978
rect 25394 56926 25732 56978
rect 25340 56924 25732 56926
rect 25340 56914 25396 56924
rect 25340 56308 25396 56318
rect 25340 56214 25396 56252
rect 25676 55298 25732 56924
rect 25676 55246 25678 55298
rect 25730 55246 25732 55298
rect 25676 55234 25732 55246
rect 24892 49140 24948 49150
rect 24892 49046 24948 49084
rect 24780 47518 24782 47570
rect 24834 47518 24836 47570
rect 24780 47506 24836 47518
rect 25004 47012 25060 55020
rect 25564 55074 25620 55086
rect 25564 55022 25566 55074
rect 25618 55022 25620 55074
rect 25228 52834 25284 52846
rect 25228 52782 25230 52834
rect 25282 52782 25284 52834
rect 25116 52162 25172 52174
rect 25116 52110 25118 52162
rect 25170 52110 25172 52162
rect 25116 51940 25172 52110
rect 25116 51874 25172 51884
rect 25228 50428 25284 52782
rect 25340 52052 25396 52062
rect 25340 51602 25396 51996
rect 25340 51550 25342 51602
rect 25394 51550 25396 51602
rect 25340 51538 25396 51550
rect 25564 50428 25620 55022
rect 25788 51602 25844 57036
rect 25900 53396 25956 59500
rect 26012 53956 26068 59948
rect 26348 60004 26404 60014
rect 26348 59910 26404 59948
rect 27692 59892 27748 60956
rect 27692 59798 27748 59836
rect 27804 63140 27860 63150
rect 27804 61794 27860 63084
rect 27804 61742 27806 61794
rect 27858 61742 27860 61794
rect 27804 61682 27860 61742
rect 28476 63028 28532 63038
rect 28476 61796 28532 62972
rect 28588 62020 28644 63868
rect 28924 63830 28980 63868
rect 29484 63922 29540 63934
rect 29484 63870 29486 63922
rect 29538 63870 29540 63922
rect 29484 63700 29540 63870
rect 29484 63634 29540 63644
rect 29260 63028 29316 63038
rect 29260 62934 29316 62972
rect 29596 63028 29652 63038
rect 29596 62934 29652 62972
rect 29820 62804 29876 63980
rect 29932 63924 29988 63934
rect 29932 63830 29988 63868
rect 29708 62748 29876 62804
rect 29932 63138 29988 63150
rect 29932 63086 29934 63138
rect 29986 63086 29988 63138
rect 29484 62356 29540 62366
rect 29484 62262 29540 62300
rect 28588 61954 28644 61964
rect 29036 62242 29092 62254
rect 29036 62190 29038 62242
rect 29090 62190 29092 62242
rect 28476 61740 28644 61796
rect 27804 61630 27806 61682
rect 27858 61630 27860 61682
rect 27580 59218 27636 59230
rect 27580 59166 27582 59218
rect 27634 59166 27636 59218
rect 26012 53890 26068 53900
rect 26348 59108 26404 59118
rect 25900 53330 25956 53340
rect 25788 51550 25790 51602
rect 25842 51550 25844 51602
rect 25228 50372 25508 50428
rect 25564 50372 25732 50428
rect 25228 49812 25284 49822
rect 25228 49718 25284 49756
rect 25340 49364 25396 49374
rect 25228 48804 25284 48814
rect 25228 47124 25284 48748
rect 25340 48466 25396 49308
rect 25340 48414 25342 48466
rect 25394 48414 25396 48466
rect 25340 48402 25396 48414
rect 25452 48244 25508 50372
rect 25564 49922 25620 49934
rect 25564 49870 25566 49922
rect 25618 49870 25620 49922
rect 25564 49364 25620 49870
rect 25564 49298 25620 49308
rect 25676 48468 25732 50372
rect 25788 48692 25844 51550
rect 26124 51268 26180 51278
rect 26124 50708 26180 51212
rect 26124 49810 26180 50652
rect 26124 49758 26126 49810
rect 26178 49758 26180 49810
rect 26124 49746 26180 49758
rect 25900 49698 25956 49710
rect 25900 49646 25902 49698
rect 25954 49646 25956 49698
rect 25900 49140 25956 49646
rect 25900 49074 25956 49084
rect 25788 48626 25844 48636
rect 24780 46956 25060 47012
rect 25116 47068 25284 47124
rect 25340 48188 25508 48244
rect 25564 48412 25732 48468
rect 24668 46676 24724 46686
rect 24668 46582 24724 46620
rect 24556 45724 24724 45780
rect 23996 43708 24164 43764
rect 23772 43598 23774 43650
rect 23826 43598 23828 43650
rect 22988 41860 23044 41870
rect 22876 41858 23044 41860
rect 22876 41806 22990 41858
rect 23042 41806 23044 41858
rect 22876 41804 23044 41806
rect 22988 41794 23044 41804
rect 22988 41524 23044 41534
rect 22876 41300 22932 41310
rect 22876 41206 22932 41244
rect 22876 40964 22932 40974
rect 22876 40626 22932 40908
rect 22876 40574 22878 40626
rect 22930 40574 22932 40626
rect 22876 40562 22932 40574
rect 22988 40516 23044 41468
rect 22988 40450 23044 40460
rect 22764 39790 22766 39842
rect 22818 39790 22820 39842
rect 22764 39778 22820 39790
rect 22204 39730 22260 39742
rect 22204 39678 22206 39730
rect 22258 39678 22260 39730
rect 22204 39620 22260 39678
rect 22652 39620 22708 39630
rect 22204 39618 22708 39620
rect 22204 39566 22654 39618
rect 22706 39566 22708 39618
rect 22204 39564 22708 39566
rect 22652 39554 22708 39564
rect 22092 39394 22148 39406
rect 22092 39342 22094 39394
rect 22146 39342 22148 39394
rect 22092 39060 22148 39342
rect 22204 39396 22260 39406
rect 22764 39396 22820 39406
rect 22204 39302 22260 39340
rect 22428 39394 22820 39396
rect 22428 39342 22766 39394
rect 22818 39342 22820 39394
rect 22428 39340 22820 39342
rect 22092 38994 22148 39004
rect 22204 38836 22260 38846
rect 22260 38822 22372 38836
rect 22260 38780 22318 38822
rect 22204 38770 22260 38780
rect 22316 38770 22318 38780
rect 22370 38770 22372 38822
rect 22316 38758 22372 38770
rect 22428 38668 22484 39340
rect 22764 39330 22820 39340
rect 22988 39060 23044 39070
rect 23100 39060 23156 41916
rect 23324 41748 23380 41758
rect 23324 41298 23380 41692
rect 23324 41246 23326 41298
rect 23378 41246 23380 41298
rect 23324 41234 23380 41246
rect 23436 41748 23492 43484
rect 23772 42532 23828 43598
rect 23772 42466 23828 42476
rect 23996 43538 24052 43550
rect 23996 43486 23998 43538
rect 24050 43486 24052 43538
rect 23548 42308 23604 42318
rect 23548 41970 23604 42252
rect 23996 41972 24052 43486
rect 24108 43540 24164 43708
rect 24108 43474 24164 43484
rect 24220 43708 24388 43764
rect 24668 45108 24724 45724
rect 24780 45220 24836 46956
rect 25116 45556 25172 47068
rect 25228 46900 25284 46910
rect 25228 46786 25284 46844
rect 25228 46734 25230 46786
rect 25282 46734 25284 46786
rect 25228 46722 25284 46734
rect 25340 46788 25396 48188
rect 25564 47068 25620 48412
rect 25676 48244 25732 48254
rect 25676 48242 26068 48244
rect 25676 48190 25678 48242
rect 25730 48190 26068 48242
rect 25676 48188 26068 48190
rect 25676 48178 25732 48188
rect 26012 47348 26068 48188
rect 26124 48132 26180 48142
rect 26124 48038 26180 48076
rect 26012 47292 26292 47348
rect 25564 47012 26068 47068
rect 25340 46722 25396 46732
rect 25452 46674 25508 46686
rect 25452 46622 25454 46674
rect 25506 46622 25508 46674
rect 25452 46116 25508 46622
rect 25676 46674 25732 46686
rect 25676 46622 25678 46674
rect 25730 46622 25732 46674
rect 25564 46564 25620 46602
rect 25564 46498 25620 46508
rect 25452 46050 25508 46060
rect 25676 45892 25732 46622
rect 25676 45826 25732 45836
rect 25788 46674 25844 46686
rect 25788 46622 25790 46674
rect 25842 46622 25844 46674
rect 25788 46004 25844 46622
rect 26012 46564 26068 47012
rect 26236 46898 26292 47292
rect 26236 46846 26238 46898
rect 26290 46846 26292 46898
rect 26236 46834 26292 46846
rect 26012 46508 26292 46564
rect 26236 46340 26292 46508
rect 26236 46274 26292 46284
rect 25116 45500 25732 45556
rect 25340 45332 25396 45342
rect 24780 45154 24836 45164
rect 25228 45330 25396 45332
rect 25228 45278 25342 45330
rect 25394 45278 25396 45330
rect 25228 45276 25396 45278
rect 24668 44322 24724 45052
rect 24668 44270 24670 44322
rect 24722 44270 24724 44322
rect 24668 43764 24724 44270
rect 24892 44884 24948 44894
rect 24668 43762 24836 43764
rect 24668 43710 24670 43762
rect 24722 43710 24836 43762
rect 24668 43708 24836 43710
rect 24220 42980 24276 43708
rect 24668 43698 24724 43708
rect 23548 41918 23550 41970
rect 23602 41918 23604 41970
rect 23548 41906 23604 41918
rect 23772 41916 23996 41972
rect 23548 41748 23604 41758
rect 23436 41692 23548 41748
rect 22988 39058 23156 39060
rect 22988 39006 22990 39058
rect 23042 39006 23156 39058
rect 22988 39004 23156 39006
rect 23212 41188 23268 41198
rect 22988 38994 23044 39004
rect 22204 38612 22484 38668
rect 22764 38836 22820 38846
rect 22764 38668 22820 38780
rect 22652 38612 22708 38622
rect 22764 38612 22932 38668
rect 22204 38162 22260 38612
rect 22204 38110 22206 38162
rect 22258 38110 22260 38162
rect 22204 38098 22260 38110
rect 22316 38500 22372 38510
rect 22316 38050 22372 38444
rect 22316 37998 22318 38050
rect 22370 37998 22372 38050
rect 22092 37826 22148 37838
rect 22092 37774 22094 37826
rect 22146 37774 22148 37826
rect 22092 36260 22148 37774
rect 22316 36372 22372 37998
rect 22540 38388 22596 38398
rect 22428 37380 22484 37390
rect 22428 37286 22484 37324
rect 22428 36372 22484 36382
rect 22316 36316 22428 36372
rect 22428 36306 22484 36316
rect 22204 36260 22260 36298
rect 22092 36204 22204 36260
rect 22260 36204 22372 36260
rect 22204 36194 22260 36204
rect 22204 36036 22260 36046
rect 22204 35026 22260 35980
rect 22316 35364 22372 36204
rect 22316 35298 22372 35308
rect 22204 34974 22206 35026
rect 22258 34974 22260 35026
rect 22204 34962 22260 34974
rect 22428 33684 22484 33694
rect 22036 31724 22260 31780
rect 21980 31714 22036 31724
rect 22204 30210 22260 31724
rect 22204 30158 22206 30210
rect 22258 30158 22260 30210
rect 22204 30146 22260 30158
rect 22428 30210 22484 33628
rect 22428 30158 22430 30210
rect 22482 30158 22484 30210
rect 22428 29988 22484 30158
rect 22428 29922 22484 29932
rect 22428 29538 22484 29550
rect 22428 29486 22430 29538
rect 22482 29486 22484 29538
rect 21756 29428 21812 29438
rect 21756 29334 21812 29372
rect 21644 29148 21812 29204
rect 21644 28196 21700 28206
rect 21644 27860 21700 28140
rect 18956 18386 19012 18396
rect 19180 20972 19348 21028
rect 19404 23996 19572 24052
rect 20188 23996 20468 24052
rect 20524 26852 20692 26908
rect 21420 27858 21700 27860
rect 21420 27806 21646 27858
rect 21698 27806 21700 27858
rect 21420 27804 21700 27806
rect 19404 21028 19460 23996
rect 19628 23940 19684 23950
rect 19516 23884 19628 23940
rect 19516 23826 19572 23884
rect 19628 23874 19684 23884
rect 19516 23774 19518 23826
rect 19570 23774 19572 23826
rect 19516 23380 19572 23774
rect 19628 23714 19684 23726
rect 19628 23662 19630 23714
rect 19682 23662 19684 23714
rect 19628 23604 19684 23662
rect 19628 23538 19684 23548
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19964 23380 20020 23390
rect 19516 23378 20020 23380
rect 19516 23326 19966 23378
rect 20018 23326 20020 23378
rect 19516 23324 20020 23326
rect 19516 21812 19572 23324
rect 19964 23314 20020 23324
rect 19964 22596 20020 22606
rect 19964 22370 20020 22540
rect 19964 22318 19966 22370
rect 20018 22318 20020 22370
rect 19964 22306 20020 22318
rect 19628 22260 19684 22298
rect 19628 22194 19684 22204
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 19516 21746 19572 21756
rect 19404 20972 19572 21028
rect 19068 16772 19124 16782
rect 19068 16678 19124 16716
rect 19068 16548 19124 16558
rect 18956 15652 19012 15662
rect 18956 15538 19012 15596
rect 18956 15486 18958 15538
rect 19010 15486 19012 15538
rect 18956 15474 19012 15486
rect 18284 15138 18340 15148
rect 17724 14366 17726 14418
rect 17778 14366 17780 14418
rect 17724 14354 17780 14366
rect 18732 15092 18900 15148
rect 18956 15092 19012 15102
rect 17612 13918 17614 13970
rect 17666 13918 17668 13970
rect 17612 13906 17668 13918
rect 17948 13636 18004 13646
rect 17948 13542 18004 13580
rect 18172 13636 18228 13646
rect 18620 13636 18676 13646
rect 18172 13634 18452 13636
rect 18172 13582 18174 13634
rect 18226 13582 18452 13634
rect 18172 13580 18452 13582
rect 18172 13570 18228 13580
rect 17500 13076 17556 13086
rect 18284 13076 18340 13086
rect 17388 13074 17556 13076
rect 17388 13022 17502 13074
rect 17554 13022 17556 13074
rect 17388 13020 17556 13022
rect 17388 12516 17444 13020
rect 17500 13010 17556 13020
rect 18172 13020 18284 13076
rect 17276 12404 17332 12414
rect 17164 12402 17332 12404
rect 17164 12350 17278 12402
rect 17330 12350 17332 12402
rect 17164 12348 17332 12350
rect 17276 12338 17332 12348
rect 17388 11956 17444 12460
rect 17500 12180 17556 12190
rect 17500 12086 17556 12124
rect 17948 12178 18004 12190
rect 17948 12126 17950 12178
rect 18002 12126 18004 12178
rect 17836 11956 17892 11966
rect 17388 11890 17444 11900
rect 17724 11900 17836 11956
rect 17724 10836 17780 11900
rect 17836 11890 17892 11900
rect 17948 11844 18004 12126
rect 18060 12180 18116 12190
rect 18060 12086 18116 12124
rect 17948 11778 18004 11788
rect 17724 10770 17780 10780
rect 17836 11508 17892 11518
rect 17836 10834 17892 11452
rect 17836 10782 17838 10834
rect 17890 10782 17892 10834
rect 17836 10770 17892 10782
rect 18060 10612 18116 10622
rect 17948 10610 18116 10612
rect 17948 10558 18062 10610
rect 18114 10558 18116 10610
rect 17948 10556 18116 10558
rect 16828 10434 16884 10444
rect 17500 10500 17556 10510
rect 16828 9940 16884 9950
rect 16716 9938 16884 9940
rect 16716 9886 16830 9938
rect 16882 9886 16884 9938
rect 16716 9884 16884 9886
rect 16828 9874 16884 9884
rect 17164 9940 17220 9950
rect 17164 9828 17220 9884
rect 16940 9826 17220 9828
rect 16940 9774 17166 9826
rect 17218 9774 17220 9826
rect 16940 9772 17220 9774
rect 16828 9044 16884 9054
rect 16940 9044 16996 9772
rect 17164 9762 17220 9772
rect 17500 9828 17556 10444
rect 17948 10276 18004 10556
rect 18060 10546 18116 10556
rect 17612 10220 18004 10276
rect 17612 9938 17668 10220
rect 17612 9886 17614 9938
rect 17666 9886 17668 9938
rect 17612 9874 17668 9886
rect 17724 10052 17780 10062
rect 17500 9762 17556 9772
rect 17724 9828 17780 9996
rect 18172 9940 18228 13020
rect 18284 12982 18340 13020
rect 18396 12180 18452 13580
rect 18620 13188 18676 13580
rect 18620 13122 18676 13132
rect 18620 12180 18676 12190
rect 18396 12178 18676 12180
rect 18396 12126 18622 12178
rect 18674 12126 18676 12178
rect 18396 12124 18676 12126
rect 18732 12180 18788 15092
rect 18956 14642 19012 15036
rect 18956 14590 18958 14642
rect 19010 14590 19012 14642
rect 18956 14578 19012 14590
rect 18844 13076 18900 13086
rect 18844 12402 18900 13020
rect 18844 12350 18846 12402
rect 18898 12350 18900 12402
rect 18844 12338 18900 12350
rect 18956 12738 19012 12750
rect 18956 12686 18958 12738
rect 19010 12686 19012 12738
rect 18956 12404 19012 12686
rect 18956 12338 19012 12348
rect 19068 12292 19124 16492
rect 19180 15092 19236 20972
rect 19292 16098 19348 16110
rect 19292 16046 19294 16098
rect 19346 16046 19348 16098
rect 19292 15652 19348 16046
rect 19404 15988 19460 15998
rect 19404 15894 19460 15932
rect 19292 15586 19348 15596
rect 19292 15428 19348 15438
rect 19292 15334 19348 15372
rect 19404 15204 19460 15242
rect 19404 15138 19460 15148
rect 19180 12404 19236 15036
rect 19180 12338 19236 12348
rect 19516 12292 19572 20972
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 20076 18676 20132 18686
rect 19852 18564 19908 18574
rect 19628 18562 19908 18564
rect 19628 18510 19854 18562
rect 19906 18510 19908 18562
rect 19628 18508 19908 18510
rect 19628 16772 19684 18508
rect 19852 18498 19908 18508
rect 19964 18562 20020 18574
rect 19964 18510 19966 18562
rect 20018 18510 20020 18562
rect 19964 18452 20020 18510
rect 19964 18386 20020 18396
rect 19740 18340 19796 18350
rect 19740 18228 19796 18284
rect 19852 18228 19908 18238
rect 19740 18226 19908 18228
rect 19740 18174 19854 18226
rect 19906 18174 19908 18226
rect 19740 18172 19908 18174
rect 19852 18162 19908 18172
rect 19964 17780 20020 17790
rect 20076 17780 20132 18620
rect 19964 17778 20132 17780
rect 19964 17726 19966 17778
rect 20018 17726 20132 17778
rect 19964 17724 20132 17726
rect 19964 17714 20020 17724
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19740 16772 19796 16782
rect 19628 16770 19796 16772
rect 19628 16718 19742 16770
rect 19794 16718 19796 16770
rect 19628 16716 19796 16718
rect 19628 16324 19684 16334
rect 19628 15426 19684 16268
rect 19740 16212 19796 16716
rect 20188 16436 20244 23996
rect 20412 23826 20468 23838
rect 20412 23774 20414 23826
rect 20466 23774 20468 23826
rect 20412 23716 20468 23774
rect 20412 23650 20468 23660
rect 20300 23380 20356 23390
rect 20300 21474 20356 23324
rect 20524 23042 20580 26852
rect 21420 24722 21476 27804
rect 21644 27794 21700 27804
rect 21756 26908 21812 29148
rect 22316 27972 22372 27982
rect 22428 27972 22484 29486
rect 22316 27970 22484 27972
rect 22316 27918 22318 27970
rect 22370 27918 22484 27970
rect 22316 27916 22484 27918
rect 22316 27906 22372 27916
rect 21420 24670 21422 24722
rect 21474 24670 21476 24722
rect 21420 24658 21476 24670
rect 21644 26852 21812 26908
rect 22540 26908 22596 38332
rect 22652 37266 22708 38556
rect 22764 37826 22820 37838
rect 22764 37774 22766 37826
rect 22818 37774 22820 37826
rect 22764 37492 22820 37774
rect 22764 37426 22820 37436
rect 22652 37214 22654 37266
rect 22706 37214 22708 37266
rect 22652 36706 22708 37214
rect 22652 36654 22654 36706
rect 22706 36654 22708 36706
rect 22652 36642 22708 36654
rect 22764 36596 22820 36606
rect 22876 36596 22932 38612
rect 23100 38164 23156 38174
rect 23100 38070 23156 38108
rect 23100 37940 23156 37950
rect 22764 36594 22932 36596
rect 22764 36542 22766 36594
rect 22818 36542 22932 36594
rect 22764 36540 22932 36542
rect 22988 37042 23044 37054
rect 22988 36990 22990 37042
rect 23042 36990 23044 37042
rect 22764 36530 22820 36540
rect 22988 36484 23044 36990
rect 23100 36594 23156 37884
rect 23100 36542 23102 36594
rect 23154 36542 23156 36594
rect 23100 36530 23156 36542
rect 22988 36418 23044 36428
rect 22988 36260 23044 36270
rect 22988 34354 23044 36204
rect 22988 34302 22990 34354
rect 23042 34302 23044 34354
rect 22988 34132 23044 34302
rect 22764 34076 22988 34132
rect 22764 30212 22820 34076
rect 22988 34066 23044 34076
rect 23212 31220 23268 41132
rect 23436 41086 23492 41692
rect 23548 41682 23604 41692
rect 23772 41300 23828 41916
rect 23996 41878 24052 41916
rect 24108 42924 24276 42980
rect 24332 43538 24388 43550
rect 24332 43486 24334 43538
rect 24386 43486 24388 43538
rect 23884 41748 23940 41758
rect 23884 41746 24052 41748
rect 23884 41694 23886 41746
rect 23938 41694 24052 41746
rect 23884 41692 24052 41694
rect 23884 41682 23940 41692
rect 23324 41030 23492 41086
rect 23548 41244 23828 41300
rect 23884 41524 23940 41534
rect 23324 40068 23380 41030
rect 23436 40292 23492 40302
rect 23436 40198 23492 40236
rect 23324 40012 23492 40068
rect 23324 39394 23380 39406
rect 23324 39342 23326 39394
rect 23378 39342 23380 39394
rect 23324 38948 23380 39342
rect 23324 38854 23380 38892
rect 23436 38724 23492 40012
rect 23324 38668 23492 38724
rect 23324 37268 23380 38668
rect 23436 38388 23492 38398
rect 23436 37490 23492 38332
rect 23436 37438 23438 37490
rect 23490 37438 23492 37490
rect 23436 37426 23492 37438
rect 23324 37212 23492 37268
rect 23324 36706 23380 36718
rect 23324 36654 23326 36706
rect 23378 36654 23380 36706
rect 23324 35922 23380 36654
rect 23324 35870 23326 35922
rect 23378 35870 23380 35922
rect 23324 35858 23380 35870
rect 23324 34018 23380 34030
rect 23324 33966 23326 34018
rect 23378 33966 23380 34018
rect 23324 33684 23380 33966
rect 23324 33618 23380 33628
rect 23436 32116 23492 37212
rect 23548 36484 23604 41244
rect 23772 41076 23828 41086
rect 23772 40982 23828 41020
rect 23884 40740 23940 41468
rect 23884 40626 23940 40684
rect 23884 40574 23886 40626
rect 23938 40574 23940 40626
rect 23884 40562 23940 40574
rect 23660 40404 23716 40414
rect 23660 39732 23716 40348
rect 23772 40178 23828 40190
rect 23772 40126 23774 40178
rect 23826 40126 23828 40178
rect 23772 39842 23828 40126
rect 23996 39956 24052 41692
rect 24108 41300 24164 42924
rect 24108 41234 24164 41244
rect 24220 42754 24276 42766
rect 24220 42702 24222 42754
rect 24274 42702 24276 42754
rect 24220 41636 24276 42702
rect 24332 42308 24388 43486
rect 24332 42242 24388 42252
rect 24668 42644 24724 42654
rect 24332 42084 24388 42094
rect 24332 41860 24388 42028
rect 24444 41860 24500 41870
rect 24332 41858 24500 41860
rect 24332 41806 24446 41858
rect 24498 41806 24500 41858
rect 24332 41804 24500 41806
rect 24444 41794 24500 41804
rect 24108 41076 24164 41086
rect 24220 41076 24276 41580
rect 24444 41188 24500 41198
rect 24164 41020 24276 41076
rect 24332 41132 24444 41188
rect 24108 41010 24164 41020
rect 24220 40852 24276 40862
rect 24220 40628 24276 40796
rect 24220 40534 24276 40572
rect 24332 39956 24388 41132
rect 24444 41122 24500 41132
rect 24668 40628 24724 42588
rect 24780 41524 24836 43708
rect 24892 41748 24948 44828
rect 25004 44210 25060 44222
rect 25004 44158 25006 44210
rect 25058 44158 25060 44210
rect 25004 41972 25060 44158
rect 25228 42868 25284 45276
rect 25340 45266 25396 45276
rect 25564 45218 25620 45230
rect 25564 45166 25566 45218
rect 25618 45166 25620 45218
rect 25564 44212 25620 45166
rect 25564 43876 25620 44156
rect 25676 44212 25732 45500
rect 25788 44884 25844 45948
rect 26236 45890 26292 45902
rect 26236 45838 26238 45890
rect 26290 45838 26292 45890
rect 26012 45220 26068 45230
rect 26012 45126 26068 45164
rect 25788 44818 25844 44828
rect 25676 44210 25844 44212
rect 25676 44158 25678 44210
rect 25730 44158 25844 44210
rect 25676 44156 25844 44158
rect 25676 44146 25732 44156
rect 25564 43810 25620 43820
rect 25564 43428 25620 43438
rect 25564 43334 25620 43372
rect 25004 41906 25060 41916
rect 25116 42812 25284 42868
rect 24892 41692 25060 41748
rect 24780 41458 24836 41468
rect 24668 40534 24724 40572
rect 24780 41186 24836 41198
rect 24780 41134 24782 41186
rect 24834 41134 24836 41186
rect 24780 40178 24836 41134
rect 24780 40126 24782 40178
rect 24834 40126 24836 40178
rect 24780 40114 24836 40126
rect 23996 39890 24052 39900
rect 24220 39900 24388 39956
rect 24668 39956 24724 39966
rect 23772 39790 23774 39842
rect 23826 39790 23828 39842
rect 23772 39778 23828 39790
rect 24108 39844 24164 39854
rect 23660 39666 23716 39676
rect 24108 39620 24164 39788
rect 23884 39564 24164 39620
rect 23660 39506 23716 39518
rect 23660 39454 23662 39506
rect 23714 39454 23716 39506
rect 23660 38164 23716 39454
rect 23660 38098 23716 38108
rect 23884 37490 23940 39564
rect 24108 39396 24164 39406
rect 24108 39058 24164 39340
rect 24108 39006 24110 39058
rect 24162 39006 24164 39058
rect 24108 38994 24164 39006
rect 24220 39058 24276 39900
rect 24444 39732 24500 39742
rect 24444 39638 24500 39676
rect 24332 39508 24388 39518
rect 24332 39506 24500 39508
rect 24332 39454 24334 39506
rect 24386 39454 24500 39506
rect 24332 39452 24500 39454
rect 24332 39442 24388 39452
rect 24444 39396 24500 39452
rect 24444 39330 24500 39340
rect 24220 39006 24222 39058
rect 24274 39006 24276 39058
rect 24220 38994 24276 39006
rect 24444 39060 24500 39070
rect 24332 38948 24388 38958
rect 24444 38948 24500 39004
rect 24332 38946 24500 38948
rect 24332 38894 24334 38946
rect 24386 38894 24500 38946
rect 24332 38892 24500 38894
rect 23884 37438 23886 37490
rect 23938 37438 23940 37490
rect 23884 37426 23940 37438
rect 23996 38834 24052 38846
rect 23996 38782 23998 38834
rect 24050 38782 24052 38834
rect 23996 37492 24052 38782
rect 23996 37426 24052 37436
rect 24108 38164 24164 38174
rect 23996 36484 24052 36494
rect 23548 36428 23716 36484
rect 23548 36260 23604 36270
rect 23548 36166 23604 36204
rect 23548 34132 23604 34142
rect 23548 34038 23604 34076
rect 23548 33684 23604 33694
rect 23660 33684 23716 36428
rect 23996 36390 24052 36428
rect 23604 33628 23716 33684
rect 23772 35364 23828 35374
rect 23548 33618 23604 33628
rect 23772 33572 23828 35308
rect 24108 34580 24164 38108
rect 24332 37492 24388 38892
rect 24220 37490 24388 37492
rect 24220 37438 24334 37490
rect 24386 37438 24388 37490
rect 24220 37436 24388 37438
rect 24220 36036 24276 37436
rect 24332 37426 24388 37436
rect 24556 38836 24612 38846
rect 24668 38836 24724 39900
rect 24892 39508 24948 39518
rect 24892 39414 24948 39452
rect 25004 39284 25060 41692
rect 25116 41300 25172 42812
rect 25788 42644 25844 44156
rect 26236 43540 26292 45838
rect 26348 45220 26404 59052
rect 27356 59108 27412 59118
rect 27580 59108 27636 59166
rect 27356 59106 27636 59108
rect 27356 59054 27358 59106
rect 27410 59054 27636 59106
rect 27356 59052 27636 59054
rect 27132 57538 27188 57550
rect 27132 57486 27134 57538
rect 27186 57486 27188 57538
rect 27132 57428 27188 57486
rect 27356 57428 27412 59052
rect 27804 58658 27860 61630
rect 28476 61572 28532 61582
rect 28252 60900 28308 60910
rect 28252 60806 28308 60844
rect 28364 60898 28420 60910
rect 28364 60846 28366 60898
rect 28418 60846 28420 60898
rect 27916 60788 27972 60798
rect 27916 60694 27972 60732
rect 28364 60788 28420 60846
rect 28364 60722 28420 60732
rect 28364 60564 28420 60574
rect 28476 60564 28532 61516
rect 28364 60562 28532 60564
rect 28364 60510 28366 60562
rect 28418 60510 28532 60562
rect 28364 60508 28532 60510
rect 28588 61346 28644 61740
rect 29036 61684 29092 62190
rect 29260 62242 29316 62254
rect 29260 62190 29262 62242
rect 29314 62190 29316 62242
rect 29260 61908 29316 62190
rect 29260 61842 29316 61852
rect 29708 61794 29764 62748
rect 29820 62580 29876 62590
rect 29820 62486 29876 62524
rect 29708 61742 29710 61794
rect 29762 61742 29764 61794
rect 29708 61730 29764 61742
rect 29932 62020 29988 63086
rect 29372 61684 29428 61694
rect 29036 61682 29428 61684
rect 29036 61630 29374 61682
rect 29426 61630 29428 61682
rect 29036 61628 29428 61630
rect 29148 61460 29204 61470
rect 28588 61294 28590 61346
rect 28642 61294 28644 61346
rect 28588 60564 28644 61294
rect 29036 61404 29148 61460
rect 28812 60564 28868 60574
rect 28588 60562 28868 60564
rect 28588 60510 28814 60562
rect 28866 60510 28868 60562
rect 28588 60508 28868 60510
rect 28364 60498 28420 60508
rect 28252 59778 28308 59790
rect 28252 59726 28254 59778
rect 28306 59726 28308 59778
rect 27804 58606 27806 58658
rect 27858 58606 27860 58658
rect 27804 58594 27860 58606
rect 27916 59330 27972 59342
rect 27916 59278 27918 59330
rect 27970 59278 27972 59330
rect 27692 58324 27748 58334
rect 27692 58230 27748 58268
rect 27804 57762 27860 57774
rect 27804 57710 27806 57762
rect 27858 57710 27860 57762
rect 27804 57428 27860 57710
rect 27132 57372 27860 57428
rect 27916 57650 27972 59278
rect 28140 58658 28196 58670
rect 28140 58606 28142 58658
rect 28194 58606 28196 58658
rect 27916 57598 27918 57650
rect 27970 57598 27972 57650
rect 26684 57092 26740 57102
rect 26684 56082 26740 57036
rect 27132 56868 27188 57372
rect 27468 56980 27524 56990
rect 27468 56886 27524 56924
rect 26684 56030 26686 56082
rect 26738 56030 26740 56082
rect 26684 56018 26740 56030
rect 26908 56812 27188 56868
rect 26796 53956 26852 53966
rect 26796 53730 26852 53900
rect 26796 53678 26798 53730
rect 26850 53678 26852 53730
rect 26796 53666 26852 53678
rect 26796 53396 26852 53406
rect 26796 50706 26852 53340
rect 26796 50654 26798 50706
rect 26850 50654 26852 50706
rect 26796 49700 26852 50654
rect 26908 50036 26964 56812
rect 27468 55972 27524 55982
rect 27468 55970 27748 55972
rect 27468 55918 27470 55970
rect 27522 55918 27748 55970
rect 27468 55916 27748 55918
rect 27468 55906 27524 55916
rect 27692 55522 27748 55916
rect 27916 55860 27972 57598
rect 28028 58212 28084 58222
rect 28028 57652 28084 58156
rect 28028 57586 28084 57596
rect 28140 57092 28196 58606
rect 28252 58324 28308 59726
rect 28700 59780 28756 59790
rect 28700 59686 28756 59724
rect 28476 58658 28532 58670
rect 28812 58660 28868 60508
rect 28476 58606 28478 58658
rect 28530 58606 28532 58658
rect 28476 58546 28532 58606
rect 28476 58494 28478 58546
rect 28530 58494 28532 58546
rect 28476 58482 28532 58494
rect 28700 58604 28868 58660
rect 28252 58258 28308 58268
rect 28140 56866 28196 57036
rect 28140 56814 28142 56866
rect 28194 56814 28196 56866
rect 28140 56308 28196 56814
rect 28140 56242 28196 56252
rect 27692 55470 27694 55522
rect 27746 55470 27748 55522
rect 27692 55458 27748 55470
rect 27804 55804 27972 55860
rect 27020 54402 27076 54414
rect 27020 54350 27022 54402
rect 27074 54350 27076 54402
rect 27020 54292 27076 54350
rect 27020 54226 27076 54236
rect 27356 54290 27412 54302
rect 27356 54238 27358 54290
rect 27410 54238 27412 54290
rect 27356 53956 27412 54238
rect 27692 54292 27748 54302
rect 27692 54198 27748 54236
rect 27356 53890 27412 53900
rect 27020 53508 27076 53518
rect 27020 53506 27412 53508
rect 27020 53454 27022 53506
rect 27074 53454 27412 53506
rect 27020 53452 27412 53454
rect 27020 53442 27076 53452
rect 27356 53058 27412 53452
rect 27356 53006 27358 53058
rect 27410 53006 27412 53058
rect 27356 52994 27412 53006
rect 27692 51380 27748 51390
rect 27692 50708 27748 51324
rect 27580 50652 27692 50708
rect 27244 50596 27300 50606
rect 26908 49980 27076 50036
rect 26908 49812 26964 49822
rect 26908 49718 26964 49756
rect 26684 49644 26852 49700
rect 26460 49586 26516 49598
rect 26460 49534 26462 49586
rect 26514 49534 26516 49586
rect 26460 48580 26516 49534
rect 26460 48514 26516 48524
rect 26460 47908 26516 47918
rect 26460 46452 26516 47852
rect 26684 46788 26740 49644
rect 27020 49588 27076 49980
rect 27244 49924 27300 50540
rect 27244 49858 27300 49868
rect 27356 49700 27412 49710
rect 26908 49532 27076 49588
rect 27244 49644 27356 49700
rect 26796 48580 26852 48590
rect 26796 48354 26852 48524
rect 26796 48302 26798 48354
rect 26850 48302 26852 48354
rect 26796 48290 26852 48302
rect 26796 48132 26852 48142
rect 26796 46788 26852 48076
rect 26908 47236 26964 49532
rect 27020 49364 27076 49374
rect 27020 49138 27076 49308
rect 27020 49086 27022 49138
rect 27074 49086 27076 49138
rect 27020 49074 27076 49086
rect 27132 48468 27188 48478
rect 27244 48468 27300 49644
rect 27356 49634 27412 49644
rect 27580 48916 27636 50652
rect 27692 50614 27748 50652
rect 27692 49700 27748 49710
rect 27692 49606 27748 49644
rect 27692 49476 27748 49486
rect 27692 49026 27748 49420
rect 27692 48974 27694 49026
rect 27746 48974 27748 49026
rect 27692 48962 27748 48974
rect 27132 48466 27300 48468
rect 27132 48414 27134 48466
rect 27186 48414 27300 48466
rect 27132 48412 27300 48414
rect 27468 48860 27636 48916
rect 27132 48402 27188 48412
rect 27468 48244 27524 48860
rect 27468 47570 27524 48188
rect 27692 48692 27748 48702
rect 27468 47518 27470 47570
rect 27522 47518 27524 47570
rect 27468 47506 27524 47518
rect 27580 48130 27636 48142
rect 27580 48078 27582 48130
rect 27634 48078 27636 48130
rect 26908 47170 26964 47180
rect 27020 47236 27076 47246
rect 27580 47236 27636 48078
rect 27020 47234 27188 47236
rect 27020 47182 27022 47234
rect 27074 47182 27188 47234
rect 27020 47180 27188 47182
rect 27020 47170 27076 47180
rect 26796 46732 27076 46788
rect 26684 46722 26740 46732
rect 26796 46564 26852 46574
rect 26684 46562 26852 46564
rect 26684 46510 26798 46562
rect 26850 46510 26852 46562
rect 26684 46508 26852 46510
rect 26572 46452 26628 46462
rect 26460 46396 26572 46452
rect 26572 46358 26628 46396
rect 26684 46116 26740 46508
rect 26796 46498 26852 46508
rect 26348 45106 26404 45164
rect 26348 45054 26350 45106
rect 26402 45054 26404 45106
rect 26348 45042 26404 45054
rect 26460 46060 26740 46116
rect 25788 42550 25844 42588
rect 26124 43484 26292 43540
rect 26348 43652 26404 43662
rect 25340 42532 25396 42542
rect 25228 41972 25284 41982
rect 25228 41878 25284 41916
rect 25116 41298 25284 41300
rect 25116 41246 25118 41298
rect 25170 41246 25284 41298
rect 25116 41244 25284 41246
rect 25116 41234 25172 41244
rect 24556 38834 24724 38836
rect 24556 38782 24558 38834
rect 24610 38782 24724 38834
rect 24556 38780 24724 38782
rect 24892 39228 25060 39284
rect 25116 39732 25172 39742
rect 24556 37156 24612 38780
rect 24668 37492 24724 37502
rect 24724 37436 24836 37492
rect 24668 37426 24724 37436
rect 24556 37090 24612 37100
rect 24332 36372 24388 36382
rect 24332 36278 24388 36316
rect 24220 35970 24276 35980
rect 24332 34804 24388 34814
rect 24332 34802 24612 34804
rect 24332 34750 24334 34802
rect 24386 34750 24612 34802
rect 24332 34748 24612 34750
rect 24332 34738 24388 34748
rect 24108 34524 24388 34580
rect 23884 34132 23940 34142
rect 24220 34132 24276 34142
rect 23884 34130 24276 34132
rect 23884 34078 23886 34130
rect 23938 34078 24222 34130
rect 24274 34078 24276 34130
rect 23884 34076 24276 34078
rect 23884 34066 23940 34076
rect 24220 34066 24276 34076
rect 22988 31164 23268 31220
rect 23324 32060 23492 32116
rect 23660 33516 23828 33572
rect 23996 33684 24052 33694
rect 23324 31220 23380 32060
rect 23436 31892 23492 31902
rect 23436 31798 23492 31836
rect 22876 30882 22932 30894
rect 22876 30830 22878 30882
rect 22930 30830 22932 30882
rect 22876 30436 22932 30830
rect 22876 30370 22932 30380
rect 22764 30146 22820 30156
rect 22764 29986 22820 29998
rect 22764 29934 22766 29986
rect 22818 29934 22820 29986
rect 22764 29538 22820 29934
rect 22764 29486 22766 29538
rect 22818 29486 22820 29538
rect 22764 29474 22820 29486
rect 22988 26908 23044 31164
rect 23212 30884 23268 30894
rect 23324 30884 23380 31164
rect 23212 30882 23380 30884
rect 23212 30830 23214 30882
rect 23266 30830 23380 30882
rect 23212 30828 23380 30830
rect 23212 30818 23268 30828
rect 23436 30770 23492 30782
rect 23436 30718 23438 30770
rect 23490 30718 23492 30770
rect 23436 30436 23492 30718
rect 23436 30370 23492 30380
rect 23436 30212 23492 30222
rect 22540 26852 22820 26908
rect 20748 24612 20804 24622
rect 20748 23826 20804 24556
rect 20748 23774 20750 23826
rect 20802 23774 20804 23826
rect 20748 23762 20804 23774
rect 20524 22990 20526 23042
rect 20578 22990 20580 23042
rect 20300 21422 20302 21474
rect 20354 21422 20356 21474
rect 20300 21410 20356 21422
rect 20412 22372 20468 22382
rect 20412 20916 20468 22316
rect 20524 21700 20580 22990
rect 21532 22484 21588 22494
rect 21644 22484 21700 26852
rect 22652 26516 22708 26526
rect 22092 26404 22148 26414
rect 22092 26402 22260 26404
rect 22092 26350 22094 26402
rect 22146 26350 22260 26402
rect 22092 26348 22260 26350
rect 22092 26338 22148 26348
rect 22092 25506 22148 25518
rect 22092 25454 22094 25506
rect 22146 25454 22148 25506
rect 22092 24836 22148 25454
rect 21980 24780 22148 24836
rect 21980 24164 22036 24780
rect 22092 24612 22148 24622
rect 22092 24518 22148 24556
rect 21980 24098 22036 24108
rect 21868 23938 21924 23950
rect 22204 23940 22260 26348
rect 22652 26402 22708 26460
rect 22652 26350 22654 26402
rect 22706 26350 22708 26402
rect 22652 26338 22708 26350
rect 21868 23886 21870 23938
rect 21922 23886 21924 23938
rect 21868 22594 21924 23886
rect 21980 23884 22260 23940
rect 21980 23268 22036 23884
rect 22092 23714 22148 23726
rect 22092 23662 22094 23714
rect 22146 23662 22148 23714
rect 22092 23380 22148 23662
rect 22092 23324 22708 23380
rect 21980 23212 22484 23268
rect 21868 22542 21870 22594
rect 21922 22542 21924 22594
rect 21868 22530 21924 22542
rect 21588 22428 21700 22484
rect 22204 22484 22260 22494
rect 21532 22390 21588 22428
rect 22204 22390 22260 22428
rect 22428 22370 22484 23212
rect 22652 23266 22708 23324
rect 22652 23214 22654 23266
rect 22706 23214 22708 23266
rect 22652 23202 22708 23214
rect 22428 22318 22430 22370
rect 22482 22318 22484 22370
rect 21420 21812 21476 21822
rect 20524 21634 20580 21644
rect 20972 21810 21476 21812
rect 20972 21758 21422 21810
rect 21474 21758 21476 21810
rect 20972 21756 21476 21758
rect 20524 20916 20580 20926
rect 20412 20914 20580 20916
rect 20412 20862 20526 20914
rect 20578 20862 20580 20914
rect 20412 20860 20580 20862
rect 20524 20850 20580 20860
rect 20636 20130 20692 20142
rect 20636 20078 20638 20130
rect 20690 20078 20692 20130
rect 20636 18676 20692 20078
rect 20972 20130 21028 21756
rect 21420 21746 21476 21756
rect 21532 21700 21588 21710
rect 20972 20078 20974 20130
rect 21026 20078 21028 20130
rect 20972 20066 21028 20078
rect 21084 21474 21140 21486
rect 21084 21422 21086 21474
rect 21138 21422 21140 21474
rect 21084 20580 21140 21422
rect 21532 20914 21588 21644
rect 21980 21700 22036 21710
rect 21980 21606 22036 21644
rect 22428 21476 22484 22318
rect 22428 21410 22484 21420
rect 21532 20862 21534 20914
rect 21586 20862 21588 20914
rect 21532 20850 21588 20862
rect 21756 21362 21812 21374
rect 21756 21310 21758 21362
rect 21810 21310 21812 21362
rect 21756 20580 21812 21310
rect 21084 20524 21812 20580
rect 20636 18610 20692 18620
rect 21084 18788 21140 20524
rect 20412 18452 20468 18462
rect 20468 18396 20580 18452
rect 20412 18358 20468 18396
rect 20188 16380 20356 16436
rect 19740 16146 19796 16156
rect 20300 15876 20356 16380
rect 20524 16100 20580 18396
rect 20972 18338 21028 18350
rect 20972 18286 20974 18338
rect 21026 18286 21028 18338
rect 20748 17668 20804 17678
rect 20972 17668 21028 18286
rect 20804 17612 21028 17668
rect 20748 17574 20804 17612
rect 20524 15986 20580 16044
rect 20524 15934 20526 15986
rect 20578 15934 20580 15986
rect 20188 15820 20356 15876
rect 20412 15876 20468 15886
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 19628 15374 19630 15426
rect 19682 15374 19684 15426
rect 19628 12404 19684 15374
rect 19740 15314 19796 15326
rect 19740 15262 19742 15314
rect 19794 15262 19796 15314
rect 19740 15092 19796 15262
rect 19740 15026 19796 15036
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19628 12348 20132 12404
rect 19516 12236 19908 12292
rect 19068 12198 19124 12236
rect 18732 12124 18900 12180
rect 18284 12066 18340 12078
rect 18284 12014 18286 12066
rect 18338 12014 18340 12066
rect 18284 10836 18340 12014
rect 18620 11508 18676 12124
rect 18844 11732 18900 12124
rect 19292 12178 19348 12190
rect 19292 12126 19294 12178
rect 19346 12126 19348 12178
rect 18956 12066 19012 12078
rect 18956 12014 18958 12066
rect 19010 12014 19012 12066
rect 18956 11956 19012 12014
rect 18956 11890 19012 11900
rect 19292 11844 19348 12126
rect 19740 12066 19796 12078
rect 19740 12014 19742 12066
rect 19794 12014 19796 12066
rect 19292 11778 19348 11788
rect 19628 11956 19684 11966
rect 18844 11676 19124 11732
rect 18732 11508 18788 11518
rect 18620 11506 18788 11508
rect 18620 11454 18734 11506
rect 18786 11454 18788 11506
rect 18620 11452 18788 11454
rect 19068 11508 19124 11676
rect 19180 11508 19236 11518
rect 19068 11506 19236 11508
rect 19068 11454 19182 11506
rect 19234 11454 19236 11506
rect 19068 11452 19236 11454
rect 18732 11442 18788 11452
rect 19180 11442 19236 11452
rect 19628 11394 19684 11900
rect 19740 11844 19796 12014
rect 19740 11778 19796 11788
rect 19628 11342 19630 11394
rect 19682 11342 19684 11394
rect 19628 11330 19684 11342
rect 19740 11620 19796 11630
rect 19740 11282 19796 11564
rect 19852 11508 19908 12236
rect 19852 11442 19908 11452
rect 19740 11230 19742 11282
rect 19794 11230 19796 11282
rect 19740 11218 19796 11230
rect 19964 11284 20020 11294
rect 19964 11190 20020 11228
rect 20076 11172 20132 12348
rect 20188 12068 20244 15820
rect 20412 15782 20468 15820
rect 20300 15428 20356 15438
rect 20300 15314 20356 15372
rect 20300 15262 20302 15314
rect 20354 15262 20356 15314
rect 20300 15148 20356 15262
rect 20524 15148 20580 15934
rect 20300 15092 20580 15148
rect 20748 16098 20804 16110
rect 20748 16046 20750 16098
rect 20802 16046 20804 16098
rect 20748 15148 20804 16046
rect 20860 15204 20916 15214
rect 20748 15092 20916 15148
rect 20188 12002 20244 12012
rect 20412 11732 20468 11742
rect 20188 11620 20244 11630
rect 20244 11564 20356 11620
rect 20188 11554 20244 11564
rect 20188 11396 20244 11406
rect 20188 11302 20244 11340
rect 20076 11116 20244 11172
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 20188 10836 20244 11116
rect 18284 10770 18340 10780
rect 20076 10780 20244 10836
rect 19068 10724 19124 10734
rect 18844 10668 19068 10724
rect 18508 10612 18564 10622
rect 18508 10518 18564 10556
rect 18620 10610 18676 10622
rect 18620 10558 18622 10610
rect 18674 10558 18676 10610
rect 18284 9940 18340 9950
rect 18172 9938 18340 9940
rect 18172 9886 18286 9938
rect 18338 9886 18340 9938
rect 18172 9884 18340 9886
rect 17724 9826 18116 9828
rect 17724 9774 17726 9826
rect 17778 9774 18116 9826
rect 17724 9772 18116 9774
rect 17724 9762 17780 9772
rect 17388 9604 17444 9614
rect 17388 9510 17444 9548
rect 17612 9604 17668 9614
rect 17612 9602 17892 9604
rect 17612 9550 17614 9602
rect 17666 9550 17892 9602
rect 17612 9548 17892 9550
rect 17612 9538 17668 9548
rect 16828 9042 16996 9044
rect 16828 8990 16830 9042
rect 16882 8990 16996 9042
rect 16828 8988 16996 8990
rect 16828 8978 16884 8988
rect 16604 8820 16660 8830
rect 16604 8036 16660 8764
rect 16604 7970 16660 7980
rect 15708 7186 15764 7196
rect 15820 7644 16548 7700
rect 14588 6750 14590 6802
rect 14642 6750 14644 6802
rect 14588 6738 14644 6750
rect 15036 6692 15092 6702
rect 12348 6690 12516 6692
rect 12348 6638 12350 6690
rect 12402 6638 12516 6690
rect 12348 6636 12516 6638
rect 12348 6626 12404 6636
rect 12460 5794 12516 6636
rect 13020 6636 13524 6692
rect 14924 6690 15092 6692
rect 14924 6638 15038 6690
rect 15090 6638 15092 6690
rect 14924 6636 15092 6638
rect 13020 6132 13076 6636
rect 14028 6468 14084 6478
rect 14028 6466 14532 6468
rect 14028 6414 14030 6466
rect 14082 6414 14532 6466
rect 14028 6412 14532 6414
rect 14028 6402 14084 6412
rect 13020 5908 13076 6076
rect 12460 5742 12462 5794
rect 12514 5742 12516 5794
rect 12460 5730 12516 5742
rect 12796 5906 13076 5908
rect 12796 5854 13022 5906
rect 13074 5854 13076 5906
rect 12796 5852 13076 5854
rect 12796 5234 12852 5852
rect 13020 5842 13076 5852
rect 13692 5796 13748 5806
rect 13692 5794 14308 5796
rect 13692 5742 13694 5794
rect 13746 5742 14308 5794
rect 13692 5740 14308 5742
rect 13692 5730 13748 5740
rect 12796 5182 12798 5234
rect 12850 5182 12852 5234
rect 12796 5170 12852 5182
rect 14252 5010 14308 5740
rect 14476 5122 14532 6412
rect 14476 5070 14478 5122
rect 14530 5070 14532 5122
rect 14476 5058 14532 5070
rect 14924 5124 14980 6636
rect 15036 6626 15092 6636
rect 15148 6692 15204 6702
rect 14924 5058 14980 5068
rect 15036 5122 15092 5134
rect 15036 5070 15038 5122
rect 15090 5070 15092 5122
rect 14252 4958 14254 5010
rect 14306 4958 14308 5010
rect 14252 4946 14308 4958
rect 11900 4898 12292 4900
rect 11900 4846 11902 4898
rect 11954 4846 12292 4898
rect 11900 4844 12292 4846
rect 14028 4900 14084 4910
rect 15036 4900 15092 5070
rect 15148 5124 15204 6636
rect 15708 6578 15764 6590
rect 15708 6526 15710 6578
rect 15762 6526 15764 6578
rect 15708 5460 15764 6526
rect 15820 5796 15876 7644
rect 17836 6802 17892 9548
rect 18060 9268 18116 9772
rect 18172 9604 18228 9884
rect 18284 9874 18340 9884
rect 18620 9940 18676 10558
rect 18844 10610 18900 10668
rect 19068 10658 19124 10668
rect 19740 10724 19796 10734
rect 19740 10630 19796 10668
rect 18844 10558 18846 10610
rect 18898 10558 18900 10610
rect 18844 10546 18900 10558
rect 19180 10612 19236 10622
rect 18620 9874 18676 9884
rect 18956 10500 19012 10510
rect 18956 9938 19012 10444
rect 18956 9886 18958 9938
rect 19010 9886 19012 9938
rect 18956 9874 19012 9886
rect 18172 9538 18228 9548
rect 18396 9828 18452 9838
rect 18172 9268 18228 9278
rect 18060 9266 18228 9268
rect 18060 9214 18174 9266
rect 18226 9214 18228 9266
rect 18060 9212 18228 9214
rect 18172 9202 18228 9212
rect 17836 6750 17838 6802
rect 17890 6750 17892 6802
rect 16380 6692 16436 6702
rect 16268 6132 16324 6142
rect 16268 6038 16324 6076
rect 15820 5794 15988 5796
rect 15820 5742 15822 5794
rect 15874 5742 15988 5794
rect 15820 5740 15988 5742
rect 15820 5730 15876 5740
rect 15708 5404 15876 5460
rect 15708 5124 15764 5134
rect 15148 5068 15708 5124
rect 15148 4900 15204 5068
rect 15708 5030 15764 5068
rect 14028 4898 14196 4900
rect 14028 4846 14030 4898
rect 14082 4846 14196 4898
rect 14028 4844 14196 4846
rect 15036 4844 15204 4900
rect 15372 4900 15428 4910
rect 15372 4898 15764 4900
rect 15372 4846 15374 4898
rect 15426 4846 15764 4898
rect 15372 4844 15764 4846
rect 11900 4834 11956 4844
rect 14028 4834 14084 4844
rect 11340 4510 11342 4562
rect 11394 4510 11396 4562
rect 11340 4498 11396 4510
rect 10892 4398 10894 4450
rect 10946 4398 10948 4450
rect 10892 4386 10948 4398
rect 12908 4452 12964 4462
rect 10444 4338 10500 4350
rect 10444 4286 10446 4338
rect 10498 4286 10500 4338
rect 10444 3666 10500 4286
rect 10556 4340 10612 4350
rect 10612 4284 10724 4340
rect 10556 4274 10612 4284
rect 10444 3614 10446 3666
rect 10498 3614 10500 3666
rect 10444 3602 10500 3614
rect 10556 4116 10612 4126
rect 10332 3556 10388 3566
rect 10332 3462 10388 3500
rect 9996 3332 10052 3342
rect 9996 2996 10052 3276
rect 10108 3332 10276 3388
rect 10108 3108 10164 3332
rect 10108 3052 10276 3108
rect 9996 2940 10164 2996
rect 10108 2882 10164 2940
rect 10108 2830 10110 2882
rect 10162 2830 10164 2882
rect 10108 2818 10164 2830
rect 9772 1874 9940 1876
rect 9772 1822 9774 1874
rect 9826 1822 9940 1874
rect 9772 1820 9940 1822
rect 10220 1874 10276 3052
rect 10556 2994 10612 4060
rect 10556 2942 10558 2994
rect 10610 2942 10612 2994
rect 10556 2930 10612 2942
rect 10556 2770 10612 2782
rect 10556 2718 10558 2770
rect 10610 2718 10612 2770
rect 10444 2660 10500 2670
rect 10444 1988 10500 2604
rect 10556 2548 10612 2718
rect 10556 2482 10612 2492
rect 10220 1822 10222 1874
rect 10274 1822 10276 1874
rect 9772 1810 9828 1820
rect 10220 1810 10276 1822
rect 10332 1986 10500 1988
rect 10332 1934 10446 1986
rect 10498 1934 10500 1986
rect 10332 1932 10500 1934
rect 10332 1540 10388 1932
rect 10444 1922 10500 1932
rect 10668 1876 10724 4284
rect 10780 4338 10836 4350
rect 10780 4286 10782 4338
rect 10834 4286 10836 4338
rect 10780 2884 10836 4286
rect 12572 3668 12628 3678
rect 12908 3668 12964 4396
rect 14028 4450 14084 4462
rect 14028 4398 14030 4450
rect 14082 4398 14084 4450
rect 14028 4340 14084 4398
rect 14140 4452 14196 4844
rect 15372 4834 15428 4844
rect 14196 4396 14644 4452
rect 14140 4358 14196 4396
rect 14028 4274 14084 4284
rect 14588 4338 14644 4396
rect 14588 4286 14590 4338
rect 14642 4286 14644 4338
rect 14588 4274 14644 4286
rect 15708 4340 15764 4844
rect 15820 4562 15876 5404
rect 15932 5234 15988 5740
rect 15932 5182 15934 5234
rect 15986 5182 15988 5234
rect 15932 5170 15988 5182
rect 16380 5122 16436 6636
rect 17388 6020 17444 6030
rect 17052 6018 17444 6020
rect 17052 5966 17390 6018
rect 17442 5966 17444 6018
rect 17052 5964 17444 5966
rect 17052 5234 17108 5964
rect 17388 5954 17444 5964
rect 17612 5908 17668 5918
rect 17052 5182 17054 5234
rect 17106 5182 17108 5234
rect 17052 5170 17108 5182
rect 17500 5906 17668 5908
rect 17500 5854 17614 5906
rect 17666 5854 17668 5906
rect 17500 5852 17668 5854
rect 16380 5070 16382 5122
rect 16434 5070 16436 5122
rect 16380 5012 16436 5070
rect 16380 4946 16436 4956
rect 16828 5124 16884 5134
rect 15820 4510 15822 4562
rect 15874 4510 15876 4562
rect 15820 4498 15876 4510
rect 16828 4562 16884 5068
rect 16828 4510 16830 4562
rect 16882 4510 16884 4562
rect 16828 4498 16884 4510
rect 17388 4564 17444 4574
rect 17500 4564 17556 5852
rect 17612 5842 17668 5852
rect 17388 4562 17556 4564
rect 17388 4510 17390 4562
rect 17442 4510 17556 4562
rect 17388 4508 17556 4510
rect 17724 5124 17780 5134
rect 17388 4498 17444 4508
rect 16044 4340 16100 4350
rect 15708 4338 16100 4340
rect 15708 4286 16046 4338
rect 16098 4286 16100 4338
rect 15708 4284 16100 4286
rect 16044 4274 16100 4284
rect 17724 4338 17780 5068
rect 17724 4286 17726 4338
rect 17778 4286 17780 4338
rect 17724 4274 17780 4286
rect 17836 4340 17892 6750
rect 18284 6692 18340 6702
rect 18396 6692 18452 9772
rect 19068 7364 19124 7374
rect 19068 7270 19124 7308
rect 18340 6636 18676 6692
rect 18284 6598 18340 6636
rect 18620 5124 18676 6636
rect 18956 5908 19012 5918
rect 18956 5814 19012 5852
rect 19180 5234 19236 10556
rect 19292 10612 19348 10622
rect 19628 10612 19684 10622
rect 19292 10610 19628 10612
rect 19292 10558 19294 10610
rect 19346 10558 19628 10610
rect 19292 10556 19628 10558
rect 19292 10546 19348 10556
rect 19180 5182 19182 5234
rect 19234 5182 19236 5234
rect 19180 5170 19236 5182
rect 19292 10164 19348 10174
rect 18620 5068 19124 5124
rect 19068 4562 19124 5068
rect 19068 4510 19070 4562
rect 19122 4510 19124 4562
rect 19068 4498 19124 4510
rect 17948 4340 18004 4350
rect 17836 4338 18004 4340
rect 17836 4286 17950 4338
rect 18002 4286 18004 4338
rect 17836 4284 18004 4286
rect 17948 4274 18004 4284
rect 12572 3666 12964 3668
rect 12572 3614 12574 3666
rect 12626 3614 12964 3666
rect 12572 3612 12964 3614
rect 12572 3602 12628 3612
rect 11116 3442 11172 3454
rect 11116 3390 11118 3442
rect 11170 3390 11172 3442
rect 11116 3332 11172 3390
rect 11452 3332 11508 3342
rect 12124 3332 12180 3342
rect 11116 3266 11172 3276
rect 11228 3330 11508 3332
rect 11228 3278 11454 3330
rect 11506 3278 11508 3330
rect 11228 3276 11508 3278
rect 10892 2884 10948 2894
rect 10780 2828 10892 2884
rect 10892 2818 10948 2828
rect 11116 2770 11172 2782
rect 11116 2718 11118 2770
rect 11170 2718 11172 2770
rect 11116 2660 11172 2718
rect 11116 2594 11172 2604
rect 11228 1988 11284 3276
rect 11452 3266 11508 3276
rect 11676 3330 12180 3332
rect 11676 3278 12126 3330
rect 12178 3278 12180 3330
rect 11676 3276 12180 3278
rect 11564 2884 11620 2894
rect 11564 2212 11620 2828
rect 11564 2146 11620 2156
rect 11004 1986 11284 1988
rect 11004 1934 11230 1986
rect 11282 1934 11284 1986
rect 11004 1932 11284 1934
rect 10892 1876 10948 1886
rect 10668 1874 10948 1876
rect 10668 1822 10894 1874
rect 10946 1822 10948 1874
rect 10668 1820 10948 1822
rect 10892 1810 10948 1820
rect 10108 1484 10388 1540
rect 10108 400 10164 1484
rect 11004 400 11060 1932
rect 11228 1922 11284 1932
rect 11676 1988 11732 3276
rect 12124 3266 12180 3276
rect 12796 2882 12852 2894
rect 12796 2830 12798 2882
rect 12850 2830 12852 2882
rect 11900 2772 11956 2782
rect 11676 1986 11844 1988
rect 11676 1934 11678 1986
rect 11730 1934 11844 1986
rect 11676 1932 11844 1934
rect 11676 1922 11732 1932
rect 11788 1652 11844 1932
rect 11900 1874 11956 2716
rect 12684 2772 12740 2782
rect 12684 2678 12740 2716
rect 12460 2658 12516 2670
rect 12460 2606 12462 2658
rect 12514 2606 12516 2658
rect 11900 1822 11902 1874
rect 11954 1822 11956 1874
rect 11900 1810 11956 1822
rect 12348 1988 12404 1998
rect 12460 1988 12516 2606
rect 12796 2324 12852 2830
rect 12908 2660 12964 3612
rect 14476 4228 14532 4238
rect 15036 4228 15092 4238
rect 13692 3442 13748 3454
rect 13916 3444 13972 3454
rect 13692 3390 13694 3442
rect 13746 3390 13748 3442
rect 13692 3388 13748 3390
rect 13804 3442 13972 3444
rect 13804 3390 13918 3442
rect 13970 3390 13972 3442
rect 13804 3388 13972 3390
rect 12908 2594 12964 2604
rect 13468 3332 13524 3342
rect 13692 3332 13860 3388
rect 13916 3378 13972 3388
rect 14252 3442 14308 3454
rect 14252 3390 14254 3442
rect 14306 3390 14308 3442
rect 12348 1986 12516 1988
rect 12348 1934 12350 1986
rect 12402 1934 12516 1986
rect 12348 1932 12516 1934
rect 12572 2268 12852 2324
rect 11788 1596 11956 1652
rect 11900 400 11956 1596
rect 12348 1540 12404 1932
rect 12572 1874 12628 2268
rect 13244 2212 13300 2222
rect 13244 2118 13300 2156
rect 13468 1986 13524 3276
rect 13468 1934 13470 1986
rect 13522 1934 13524 1986
rect 13468 1922 13524 1934
rect 13692 2994 13748 3006
rect 13692 2942 13694 2994
rect 13746 2942 13748 2994
rect 12572 1822 12574 1874
rect 12626 1822 12628 1874
rect 12572 1810 12628 1822
rect 13692 1874 13748 2942
rect 13692 1822 13694 1874
rect 13746 1822 13748 1874
rect 13692 1810 13748 1822
rect 13804 1652 13860 3332
rect 14252 2884 14308 3390
rect 14252 2818 14308 2828
rect 14476 2548 14532 4172
rect 14812 4226 15092 4228
rect 14812 4174 15038 4226
rect 15090 4174 15092 4226
rect 14812 4172 15092 4174
rect 14812 3554 14868 4172
rect 15036 4162 15092 4172
rect 15484 4226 15540 4238
rect 18396 4228 18452 4238
rect 15484 4174 15486 4226
rect 15538 4174 15540 4226
rect 14812 3502 14814 3554
rect 14866 3502 14868 3554
rect 14812 3388 14868 3502
rect 15484 3554 15540 4174
rect 18060 4226 18452 4228
rect 18060 4174 18398 4226
rect 18450 4174 18452 4226
rect 18060 4172 18452 4174
rect 18060 3892 18116 4172
rect 18396 4162 18452 4172
rect 19292 4116 19348 10108
rect 19404 9938 19460 10556
rect 19628 10518 19684 10556
rect 19964 10610 20020 10622
rect 19964 10558 19966 10610
rect 20018 10558 20020 10610
rect 19404 9886 19406 9938
rect 19458 9886 19460 9938
rect 19404 9874 19460 9886
rect 19852 10500 19908 10510
rect 19852 9938 19908 10444
rect 19852 9886 19854 9938
rect 19906 9886 19908 9938
rect 19852 9874 19908 9886
rect 19964 9604 20020 10558
rect 20076 9938 20132 10780
rect 20188 10612 20244 10622
rect 20300 10612 20356 11564
rect 20188 10610 20356 10612
rect 20188 10558 20190 10610
rect 20242 10558 20356 10610
rect 20188 10556 20356 10558
rect 20188 10500 20244 10556
rect 20188 10434 20244 10444
rect 20076 9886 20078 9938
rect 20130 9886 20132 9938
rect 20076 9874 20132 9886
rect 20300 9828 20356 9838
rect 20412 9828 20468 11676
rect 20524 11172 20580 15092
rect 20860 12066 20916 15092
rect 20860 12014 20862 12066
rect 20914 12014 20916 12066
rect 20860 12002 20916 12014
rect 20748 11620 20804 11630
rect 20748 11508 20804 11564
rect 20748 11506 21028 11508
rect 20748 11454 20750 11506
rect 20802 11454 21028 11506
rect 20748 11452 21028 11454
rect 20748 11442 20804 11452
rect 20524 10722 20580 11116
rect 20636 10836 20692 10846
rect 20636 10742 20692 10780
rect 20524 10670 20526 10722
rect 20578 10670 20580 10722
rect 20524 10612 20580 10670
rect 20524 10546 20580 10556
rect 20748 10610 20804 10622
rect 20748 10558 20750 10610
rect 20802 10558 20804 10610
rect 19964 9538 20020 9548
rect 20188 9826 20468 9828
rect 20188 9774 20302 9826
rect 20354 9774 20468 9826
rect 20188 9772 20468 9774
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 19740 8932 19796 8942
rect 20188 8932 20244 9772
rect 20300 9762 20356 9772
rect 20636 9604 20692 9614
rect 20300 9602 20692 9604
rect 20300 9550 20638 9602
rect 20690 9550 20692 9602
rect 20300 9548 20692 9550
rect 20300 9042 20356 9548
rect 20636 9538 20692 9548
rect 20748 9380 20804 10558
rect 20972 10610 21028 11452
rect 20972 10558 20974 10610
rect 21026 10558 21028 10610
rect 20972 10546 21028 10558
rect 20300 8990 20302 9042
rect 20354 8990 20356 9042
rect 20300 8978 20356 8990
rect 20412 9324 20804 9380
rect 19740 8930 20244 8932
rect 19740 8878 19742 8930
rect 19794 8878 20244 8930
rect 19740 8876 20244 8878
rect 19740 8820 19796 8876
rect 19740 8754 19796 8764
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 19628 5794 19684 5806
rect 19628 5742 19630 5794
rect 19682 5742 19684 5794
rect 19516 4900 19572 4910
rect 19404 4844 19516 4900
rect 19404 4338 19460 4844
rect 19516 4834 19572 4844
rect 19628 4562 19684 5742
rect 20188 5348 20244 8876
rect 20412 7364 20468 9324
rect 21084 9268 21140 18732
rect 21196 20020 21252 20030
rect 21196 11732 21252 19964
rect 22764 19460 22820 26852
rect 22876 26852 23044 26908
rect 23100 29988 23156 29998
rect 23212 29988 23268 29998
rect 23156 29986 23268 29988
rect 23156 29934 23214 29986
rect 23266 29934 23268 29986
rect 23156 29932 23268 29934
rect 22876 26404 22932 26852
rect 22876 26290 22932 26348
rect 22876 26238 22878 26290
rect 22930 26238 22932 26290
rect 22876 26226 22932 26238
rect 22988 26180 23044 26190
rect 22988 26086 23044 26124
rect 23100 25620 23156 29932
rect 23212 29922 23268 29932
rect 23436 29652 23492 30156
rect 23100 25396 23156 25564
rect 23100 25330 23156 25340
rect 23212 29596 23436 29652
rect 23212 20132 23268 29596
rect 23436 29558 23492 29596
rect 23548 26964 23604 26974
rect 23436 26516 23492 26526
rect 23548 26516 23604 26908
rect 23660 26908 23716 33516
rect 23996 33124 24052 33628
rect 24108 33124 24164 33134
rect 23996 33122 24164 33124
rect 23996 33070 24110 33122
rect 24162 33070 24164 33122
rect 23996 33068 24164 33070
rect 23996 30996 24052 33068
rect 24108 33058 24164 33068
rect 24220 31780 24276 31790
rect 24220 31686 24276 31724
rect 24220 31220 24276 31230
rect 24220 31126 24276 31164
rect 23996 30940 24276 30996
rect 23772 30772 23828 30782
rect 23772 30770 24164 30772
rect 23772 30718 23774 30770
rect 23826 30718 24164 30770
rect 23772 30716 24164 30718
rect 23772 30706 23828 30716
rect 24108 30210 24164 30716
rect 24108 30158 24110 30210
rect 24162 30158 24164 30210
rect 24108 30146 24164 30158
rect 24108 29652 24164 29662
rect 24108 29426 24164 29596
rect 24108 29374 24110 29426
rect 24162 29374 24164 29426
rect 24108 29362 24164 29374
rect 23772 29202 23828 29214
rect 23772 29150 23774 29202
rect 23826 29150 23828 29202
rect 23772 28868 23828 29150
rect 24220 28980 24276 30940
rect 24332 29426 24388 34524
rect 24556 34354 24612 34748
rect 24556 34302 24558 34354
rect 24610 34302 24612 34354
rect 24556 34290 24612 34302
rect 24668 31780 24724 31790
rect 24668 31686 24724 31724
rect 24444 29988 24500 29998
rect 24444 29986 24612 29988
rect 24444 29934 24446 29986
rect 24498 29934 24612 29986
rect 24444 29932 24612 29934
rect 24444 29922 24500 29932
rect 24332 29374 24334 29426
rect 24386 29374 24388 29426
rect 24332 29362 24388 29374
rect 23772 28802 23828 28812
rect 24108 28924 24276 28980
rect 24444 29316 24500 29326
rect 23996 28642 24052 28654
rect 23996 28590 23998 28642
rect 24050 28590 24052 28642
rect 23996 28196 24052 28590
rect 23996 28130 24052 28140
rect 23660 26852 23940 26908
rect 23492 26460 23604 26516
rect 23436 26422 23492 26460
rect 23772 26404 23828 26414
rect 23772 26310 23828 26348
rect 23548 25396 23604 25406
rect 23436 25394 23604 25396
rect 23436 25342 23550 25394
rect 23602 25342 23604 25394
rect 23436 25340 23604 25342
rect 23436 25284 23492 25340
rect 23548 25330 23604 25340
rect 23436 25218 23492 25228
rect 22764 19394 22820 19404
rect 22876 20076 23268 20132
rect 23324 23828 23380 23838
rect 23324 22484 23380 23772
rect 23436 23492 23492 23502
rect 23436 23154 23492 23436
rect 23884 23268 23940 26852
rect 24108 24948 24164 28924
rect 24444 27748 24500 29260
rect 24556 28980 24612 29932
rect 24780 29316 24836 37436
rect 24780 29250 24836 29260
rect 24556 28924 24836 28980
rect 24780 28754 24836 28924
rect 24780 28702 24782 28754
rect 24834 28702 24836 28754
rect 24780 28690 24836 28702
rect 24668 28196 24724 28206
rect 24444 27746 24612 27748
rect 24444 27694 24446 27746
rect 24498 27694 24612 27746
rect 24444 27692 24612 27694
rect 24444 27682 24500 27692
rect 24220 26964 24276 26974
rect 24332 26964 24388 26974
rect 24220 26962 24332 26964
rect 24220 26910 24222 26962
rect 24274 26910 24332 26962
rect 24220 26908 24332 26910
rect 24220 26898 24276 26908
rect 24332 26514 24388 26908
rect 24332 26462 24334 26514
rect 24386 26462 24388 26514
rect 24332 26450 24388 26462
rect 24444 26180 24500 26190
rect 24108 24882 24164 24892
rect 24220 25396 24276 25406
rect 24220 24610 24276 25340
rect 24444 25394 24500 26124
rect 24444 25342 24446 25394
rect 24498 25342 24500 25394
rect 24444 25330 24500 25342
rect 24220 24558 24222 24610
rect 24274 24558 24276 24610
rect 24220 24546 24276 24558
rect 24444 24164 24500 24174
rect 24332 24108 24444 24164
rect 24108 23492 24164 23502
rect 23436 23102 23438 23154
rect 23490 23102 23492 23154
rect 23436 23090 23492 23102
rect 23772 23212 23940 23268
rect 23996 23436 24108 23492
rect 22652 17668 22708 17678
rect 21308 17554 21364 17566
rect 21308 17502 21310 17554
rect 21362 17502 21364 17554
rect 21308 15538 21364 17502
rect 21644 17444 21700 17454
rect 21644 17442 21924 17444
rect 21644 17390 21646 17442
rect 21698 17390 21924 17442
rect 21644 17388 21924 17390
rect 21644 17378 21700 17388
rect 21868 16994 21924 17388
rect 21868 16942 21870 16994
rect 21922 16942 21924 16994
rect 21868 16930 21924 16942
rect 22652 16996 22708 17612
rect 22652 16884 22708 16940
rect 22652 16882 22820 16884
rect 22652 16830 22654 16882
rect 22706 16830 22820 16882
rect 22652 16828 22820 16830
rect 22652 16818 22708 16828
rect 21644 16324 21700 16334
rect 21420 16100 21476 16110
rect 21420 16006 21476 16044
rect 21308 15486 21310 15538
rect 21362 15486 21364 15538
rect 21308 15474 21364 15486
rect 21644 15314 21700 16268
rect 22092 16324 22148 16334
rect 22092 16230 22148 16268
rect 21868 16212 21924 16222
rect 21868 16118 21924 16156
rect 21644 15262 21646 15314
rect 21698 15262 21700 15314
rect 21644 15250 21700 15262
rect 22428 15874 22484 15886
rect 22428 15822 22430 15874
rect 22482 15822 22484 15874
rect 22428 15314 22484 15822
rect 22428 15262 22430 15314
rect 22482 15262 22484 15314
rect 22428 15250 22484 15262
rect 22652 15426 22708 15438
rect 22652 15374 22654 15426
rect 22706 15374 22708 15426
rect 21868 15204 21924 15242
rect 22652 15148 22708 15374
rect 21868 15138 21924 15148
rect 22540 15092 22708 15148
rect 22540 14642 22596 15092
rect 22540 14590 22542 14642
rect 22594 14590 22596 14642
rect 22540 14578 22596 14590
rect 21868 14532 21924 14542
rect 21868 14438 21924 14476
rect 22764 14532 22820 16828
rect 22876 16324 22932 20076
rect 23324 20020 23380 22428
rect 23212 19908 23268 19918
rect 23324 19908 23380 19964
rect 23212 19906 23380 19908
rect 23212 19854 23214 19906
rect 23266 19854 23380 19906
rect 23212 19852 23380 19854
rect 23212 19842 23268 19852
rect 23548 19796 23604 19806
rect 23324 19794 23604 19796
rect 23324 19742 23550 19794
rect 23602 19742 23604 19794
rect 23324 19740 23604 19742
rect 23212 19236 23268 19246
rect 23324 19236 23380 19740
rect 23548 19730 23604 19740
rect 23772 19346 23828 23212
rect 23884 23044 23940 23054
rect 23996 23044 24052 23436
rect 24108 23426 24164 23436
rect 23884 23042 24276 23044
rect 23884 22990 23886 23042
rect 23938 22990 24276 23042
rect 23884 22988 24276 22990
rect 23884 22978 23940 22988
rect 24220 22370 24276 22988
rect 24220 22318 24222 22370
rect 24274 22318 24276 22370
rect 24220 22306 24276 22318
rect 24332 20244 24388 24108
rect 24444 24098 24500 24108
rect 24444 23940 24500 23950
rect 24444 23154 24500 23884
rect 24444 23102 24446 23154
rect 24498 23102 24500 23154
rect 24444 23090 24500 23102
rect 23996 20188 24388 20244
rect 23884 20020 23940 20030
rect 23884 19926 23940 19964
rect 23772 19294 23774 19346
rect 23826 19294 23828 19346
rect 23772 19282 23828 19294
rect 23212 19234 23380 19236
rect 23212 19182 23214 19234
rect 23266 19182 23380 19234
rect 23212 19180 23380 19182
rect 23212 19170 23268 19180
rect 23436 19010 23492 19022
rect 23436 18958 23438 19010
rect 23490 18958 23492 19010
rect 23436 17778 23492 18958
rect 23996 18004 24052 20188
rect 24556 20132 24612 27692
rect 24668 27186 24724 28140
rect 24668 27134 24670 27186
rect 24722 27134 24724 27186
rect 24668 24946 24724 27134
rect 24780 26292 24836 26302
rect 24780 26198 24836 26236
rect 24668 24894 24670 24946
rect 24722 24894 24724 24946
rect 24668 23492 24724 24894
rect 24892 23940 24948 39228
rect 25116 38668 25172 39676
rect 25228 38946 25284 41244
rect 25340 40290 25396 42476
rect 25676 42420 25732 42430
rect 25452 42196 25508 42206
rect 25452 42102 25508 42140
rect 25676 42194 25732 42364
rect 25676 42142 25678 42194
rect 25730 42142 25732 42194
rect 25676 42130 25732 42142
rect 25452 41858 25508 41870
rect 25452 41806 25454 41858
rect 25506 41806 25508 41858
rect 25452 41186 25508 41806
rect 25900 41300 25956 41310
rect 26124 41300 26180 43484
rect 26348 42754 26404 43596
rect 26348 42702 26350 42754
rect 26402 42702 26404 42754
rect 26236 42530 26292 42542
rect 26236 42478 26238 42530
rect 26290 42478 26292 42530
rect 26236 42308 26292 42478
rect 26236 42242 26292 42252
rect 26348 42084 26404 42702
rect 26460 43428 26516 46060
rect 26684 45892 26740 45902
rect 26572 45220 26628 45230
rect 26572 45106 26628 45164
rect 26572 45054 26574 45106
rect 26626 45054 26628 45106
rect 26572 44660 26628 45054
rect 26572 44594 26628 44604
rect 26460 42194 26516 43372
rect 26460 42142 26462 42194
rect 26514 42142 26516 42194
rect 26460 42130 26516 42142
rect 26572 43540 26628 43550
rect 26684 43540 26740 45836
rect 26796 45780 26852 45790
rect 26796 45686 26852 45724
rect 26796 45444 26908 45556
rect 27020 45444 27076 46732
rect 26796 45388 27076 45444
rect 26796 44322 26852 45388
rect 27132 45332 27188 47180
rect 27244 47180 27636 47236
rect 27244 47012 27300 47180
rect 27692 47012 27748 48636
rect 27244 46898 27300 46956
rect 27244 46846 27246 46898
rect 27298 46846 27300 46898
rect 27244 46834 27300 46846
rect 27468 46956 27748 47012
rect 27468 46788 27524 46956
rect 27468 46732 27636 46788
rect 27580 46676 27636 46732
rect 27692 46676 27748 46686
rect 27580 46674 27748 46676
rect 27580 46622 27694 46674
rect 27746 46622 27748 46674
rect 27580 46620 27748 46622
rect 27692 46610 27748 46620
rect 27804 45666 27860 55804
rect 28028 55522 28084 55534
rect 28028 55470 28030 55522
rect 28082 55470 28084 55522
rect 27916 55300 27972 55310
rect 28028 55300 28084 55470
rect 28140 55300 28196 55310
rect 28028 55298 28196 55300
rect 28028 55246 28142 55298
rect 28194 55246 28196 55298
rect 28028 55244 28196 55246
rect 27916 55206 27972 55244
rect 28140 55234 28196 55244
rect 28476 55300 28532 55310
rect 28364 55074 28420 55086
rect 28364 55022 28366 55074
rect 28418 55022 28420 55074
rect 28364 54740 28420 55022
rect 28364 54674 28420 54684
rect 27916 54628 27972 54638
rect 27916 54534 27972 54572
rect 28364 54292 28420 54302
rect 28028 52946 28084 52958
rect 28028 52894 28030 52946
rect 28082 52894 28084 52946
rect 28028 52836 28084 52894
rect 28028 50596 28084 52780
rect 28028 50530 28084 50540
rect 28252 48804 28308 48814
rect 28252 48710 28308 48748
rect 28028 48468 28084 48478
rect 28028 48374 28084 48412
rect 28364 47460 28420 54236
rect 28476 53844 28532 55244
rect 28476 53778 28532 53788
rect 28588 52836 28644 52846
rect 28588 52742 28644 52780
rect 28252 47404 28420 47460
rect 28476 49476 28532 49486
rect 28476 48242 28532 49420
rect 28476 48190 28478 48242
rect 28530 48190 28532 48242
rect 28476 47460 28532 48190
rect 27916 47234 27972 47246
rect 27916 47182 27918 47234
rect 27970 47182 27972 47234
rect 27916 46900 27972 47182
rect 27916 46834 27972 46844
rect 28140 46564 28196 46574
rect 28140 46470 28196 46508
rect 27804 45614 27806 45666
rect 27858 45614 27860 45666
rect 27804 45602 27860 45614
rect 28140 45666 28196 45678
rect 28140 45614 28142 45666
rect 28194 45614 28196 45666
rect 27020 45276 27188 45332
rect 26908 45108 26964 45118
rect 26908 45014 26964 45052
rect 26796 44270 26798 44322
rect 26850 44270 26852 44322
rect 26796 43652 26852 44270
rect 26796 43586 26852 43596
rect 27020 43652 27076 45276
rect 27580 45220 27636 45230
rect 26628 43484 26740 43540
rect 26348 42018 26404 42028
rect 26236 41972 26292 41982
rect 26572 41972 26628 43484
rect 27020 43316 27076 43596
rect 27132 45162 27188 45174
rect 27132 45110 27134 45162
rect 27186 45110 27188 45162
rect 28140 45220 28196 45614
rect 28252 45444 28308 47404
rect 28476 47394 28532 47404
rect 28588 48468 28644 48478
rect 28364 47234 28420 47246
rect 28364 47182 28366 47234
rect 28418 47182 28420 47234
rect 28364 46452 28420 47182
rect 28588 47124 28644 48412
rect 28364 46386 28420 46396
rect 28476 47068 28644 47124
rect 28476 46004 28532 47068
rect 28588 46676 28644 46686
rect 28588 46582 28644 46620
rect 28364 45892 28420 45902
rect 28364 45778 28420 45836
rect 28476 45890 28532 45948
rect 28476 45838 28478 45890
rect 28530 45838 28532 45890
rect 28476 45826 28532 45838
rect 28364 45726 28366 45778
rect 28418 45726 28420 45778
rect 28364 45714 28420 45726
rect 28252 45378 28308 45388
rect 28588 45332 28644 45342
rect 28252 45220 28308 45230
rect 28140 45218 28308 45220
rect 28140 45166 28254 45218
rect 28306 45166 28308 45218
rect 28140 45164 28308 45166
rect 27132 44322 27188 45110
rect 27356 45108 27412 45118
rect 27132 44270 27134 44322
rect 27186 44270 27188 44322
rect 27132 43428 27188 44270
rect 27244 44882 27300 44894
rect 27244 44830 27246 44882
rect 27298 44830 27300 44882
rect 27244 43652 27300 44830
rect 27356 44436 27412 45052
rect 27580 45106 27636 45164
rect 28252 45154 28308 45164
rect 28364 45220 28420 45230
rect 27580 45054 27582 45106
rect 27634 45054 27636 45106
rect 27580 45042 27636 45054
rect 27356 44322 27412 44380
rect 27356 44270 27358 44322
rect 27410 44270 27412 44322
rect 27356 44258 27412 44270
rect 27580 44660 27636 44670
rect 27580 44322 27636 44604
rect 27580 44270 27582 44322
rect 27634 44270 27636 44322
rect 27580 44258 27636 44270
rect 27916 44100 27972 44110
rect 27916 44006 27972 44044
rect 27356 43652 27412 43662
rect 27244 43596 27356 43652
rect 27356 43586 27412 43596
rect 27916 43652 27972 43662
rect 27692 43428 27748 43438
rect 27132 43362 27188 43372
rect 27356 43426 27748 43428
rect 27356 43374 27694 43426
rect 27746 43374 27748 43426
rect 27356 43372 27748 43374
rect 27020 43250 27076 43260
rect 26684 43092 26740 43102
rect 26684 42420 26740 43036
rect 27020 43036 27300 43092
rect 27020 42754 27076 43036
rect 27020 42702 27022 42754
rect 27074 42702 27076 42754
rect 27020 42690 27076 42702
rect 27132 42866 27188 42878
rect 27132 42814 27134 42866
rect 27186 42814 27188 42866
rect 26684 42194 26740 42364
rect 26684 42142 26686 42194
rect 26738 42142 26740 42194
rect 26684 42130 26740 42142
rect 26796 42642 26852 42654
rect 26796 42590 26798 42642
rect 26850 42590 26852 42642
rect 26236 41748 26292 41916
rect 26236 41682 26292 41692
rect 26460 41916 26628 41972
rect 26796 41970 26852 42590
rect 27020 41972 27076 41982
rect 26796 41918 26798 41970
rect 26850 41918 26852 41970
rect 25900 41298 26180 41300
rect 25900 41246 25902 41298
rect 25954 41246 26180 41298
rect 25900 41244 26180 41246
rect 26236 41524 26292 41534
rect 25900 41234 25956 41244
rect 25452 41134 25454 41186
rect 25506 41134 25508 41186
rect 25452 41122 25508 41134
rect 25676 41188 25732 41198
rect 25676 41094 25732 41132
rect 25900 40628 25956 40638
rect 25900 40534 25956 40572
rect 26236 40626 26292 41468
rect 26236 40574 26238 40626
rect 26290 40574 26292 40626
rect 26236 40562 26292 40574
rect 26460 40404 26516 41916
rect 26796 41906 26852 41918
rect 26908 41970 27076 41972
rect 26908 41918 27022 41970
rect 27074 41918 27076 41970
rect 26908 41916 27076 41918
rect 26572 41076 26628 41086
rect 26572 40982 26628 41020
rect 26572 40626 26628 40638
rect 26572 40574 26574 40626
rect 26626 40574 26628 40626
rect 26572 40516 26628 40574
rect 26908 40516 26964 41916
rect 27020 41906 27076 41916
rect 27132 41748 27188 42814
rect 27244 41972 27300 43036
rect 27356 42194 27412 43372
rect 27692 43362 27748 43372
rect 27356 42142 27358 42194
rect 27410 42142 27412 42194
rect 27356 42130 27412 42142
rect 27468 43204 27524 43214
rect 27244 41906 27300 41916
rect 26572 40460 26964 40516
rect 27020 41692 27188 41748
rect 26460 40348 26628 40404
rect 25340 40238 25342 40290
rect 25394 40238 25396 40290
rect 25340 40178 25396 40238
rect 25340 40126 25342 40178
rect 25394 40126 25396 40178
rect 25340 40114 25396 40126
rect 25788 40178 25844 40190
rect 25788 40126 25790 40178
rect 25842 40126 25844 40178
rect 25676 39620 25732 39630
rect 25564 39564 25676 39620
rect 25228 38894 25230 38946
rect 25282 38894 25284 38946
rect 25228 38882 25284 38894
rect 25340 39508 25396 39518
rect 25116 38612 25284 38668
rect 25228 38162 25284 38612
rect 25228 38110 25230 38162
rect 25282 38110 25284 38162
rect 25228 38098 25284 38110
rect 25228 37828 25284 37838
rect 25228 37492 25284 37772
rect 25116 37436 25284 37492
rect 25116 36596 25172 37436
rect 25340 37380 25396 39452
rect 25564 38668 25620 39564
rect 25676 39554 25732 39564
rect 25788 39396 25844 40126
rect 26460 39620 26516 39630
rect 26460 39526 26516 39564
rect 26012 39508 26068 39518
rect 25228 37324 25396 37380
rect 25452 38612 25620 38668
rect 25676 39340 25844 39396
rect 25900 39396 25956 39406
rect 25228 36708 25284 37324
rect 25340 37156 25396 37166
rect 25340 37062 25396 37100
rect 25228 36652 25396 36708
rect 25116 36540 25284 36596
rect 25228 36482 25284 36540
rect 25228 36430 25230 36482
rect 25282 36430 25284 36482
rect 25004 36260 25060 36270
rect 25004 24164 25060 36204
rect 25116 34916 25172 34926
rect 25228 34916 25284 36430
rect 25116 34914 25228 34916
rect 25116 34862 25118 34914
rect 25170 34862 25228 34914
rect 25116 34860 25228 34862
rect 25116 34850 25172 34860
rect 25228 34822 25284 34860
rect 25228 33012 25284 33022
rect 25116 32956 25228 33012
rect 25116 25508 25172 32956
rect 25228 32946 25284 32956
rect 25340 32788 25396 36652
rect 25228 32732 25396 32788
rect 25228 25730 25284 32732
rect 25452 32676 25508 38612
rect 25564 34916 25620 34926
rect 25564 34822 25620 34860
rect 25340 32620 25508 32676
rect 25340 28082 25396 32620
rect 25676 31948 25732 39340
rect 25788 39060 25844 39070
rect 25900 39060 25956 39340
rect 25844 39004 25956 39060
rect 25788 38834 25844 39004
rect 26012 38946 26068 39452
rect 26012 38894 26014 38946
rect 26066 38894 26068 38946
rect 26012 38882 26068 38894
rect 26460 39172 26516 39182
rect 25788 38782 25790 38834
rect 25842 38782 25844 38834
rect 25788 38770 25844 38782
rect 26236 38834 26292 38846
rect 26236 38782 26238 38834
rect 26290 38782 26292 38834
rect 26012 38050 26068 38062
rect 26012 37998 26014 38050
rect 26066 37998 26068 38050
rect 26012 37828 26068 37998
rect 26012 37762 26068 37772
rect 25788 37492 25844 37502
rect 25788 37398 25844 37436
rect 25452 31892 25732 31948
rect 25788 37156 25844 37166
rect 25452 28532 25508 31892
rect 25676 31780 25732 31790
rect 25676 31686 25732 31724
rect 25452 28466 25508 28476
rect 25788 28308 25844 37100
rect 26012 36372 26068 36382
rect 26012 36278 26068 36316
rect 26236 31892 26292 38782
rect 26460 38834 26516 39116
rect 26460 38782 26462 38834
rect 26514 38782 26516 38834
rect 26460 38770 26516 38782
rect 26460 38274 26516 38286
rect 26460 38222 26462 38274
rect 26514 38222 26516 38274
rect 26460 38162 26516 38222
rect 26460 38110 26462 38162
rect 26514 38110 26516 38162
rect 26460 38098 26516 38110
rect 26348 33570 26404 33582
rect 26348 33518 26350 33570
rect 26402 33518 26404 33570
rect 26348 33458 26404 33518
rect 26348 33406 26350 33458
rect 26402 33406 26404 33458
rect 26348 33394 26404 33406
rect 26012 31836 26292 31892
rect 26460 33124 26516 33134
rect 26460 31890 26516 33068
rect 26460 31838 26462 31890
rect 26514 31838 26516 31890
rect 25900 29652 25956 29662
rect 25900 29558 25956 29596
rect 25340 28030 25342 28082
rect 25394 28030 25396 28082
rect 25340 28018 25396 28030
rect 25452 28252 25844 28308
rect 25452 27860 25508 28252
rect 25564 27972 25620 27982
rect 25564 27878 25620 27916
rect 25228 25678 25230 25730
rect 25282 25678 25284 25730
rect 25228 25666 25284 25678
rect 25340 27804 25508 27860
rect 25676 27858 25732 27870
rect 25676 27806 25678 27858
rect 25730 27806 25732 27858
rect 25116 25414 25172 25452
rect 25004 24098 25060 24108
rect 24892 23884 25172 23940
rect 24668 23426 24724 23436
rect 24668 23266 24724 23278
rect 24668 23214 24670 23266
rect 24722 23214 24724 23266
rect 24668 22708 24724 23214
rect 24668 22652 25060 22708
rect 25004 22482 25060 22652
rect 25004 22430 25006 22482
rect 25058 22430 25060 22482
rect 25004 22418 25060 22430
rect 24108 20130 24612 20132
rect 24108 20078 24558 20130
rect 24610 20078 24612 20130
rect 24108 20076 24612 20078
rect 24108 20018 24164 20076
rect 24556 20066 24612 20076
rect 24108 19966 24110 20018
rect 24162 19966 24164 20018
rect 24108 19954 24164 19966
rect 23436 17726 23438 17778
rect 23490 17726 23492 17778
rect 23436 17714 23492 17726
rect 23884 17948 24052 18004
rect 23100 16996 23156 17006
rect 23100 16902 23156 16940
rect 22876 16212 22932 16268
rect 23436 16212 23492 16222
rect 23884 16212 23940 17948
rect 22876 16210 23156 16212
rect 22876 16158 22878 16210
rect 22930 16158 23156 16210
rect 22876 16156 23156 16158
rect 22876 16146 22932 16156
rect 22764 14466 22820 14476
rect 23100 15538 23156 16156
rect 23436 16210 23940 16212
rect 23436 16158 23438 16210
rect 23490 16158 23940 16210
rect 23436 16156 23940 16158
rect 23436 16146 23492 16156
rect 23100 15486 23102 15538
rect 23154 15486 23156 15538
rect 22988 12068 23044 12078
rect 21196 11666 21252 11676
rect 22540 12066 23044 12068
rect 22540 12014 22990 12066
rect 23042 12014 23044 12066
rect 22540 12012 23044 12014
rect 21756 11620 21812 11630
rect 21420 11396 21476 11406
rect 21420 11302 21476 11340
rect 21756 11394 21812 11564
rect 21756 11342 21758 11394
rect 21810 11342 21812 11394
rect 21756 11330 21812 11342
rect 22316 11396 22372 11406
rect 22316 11394 22484 11396
rect 22316 11342 22318 11394
rect 22370 11342 22484 11394
rect 22316 11340 22484 11342
rect 22316 11330 22372 11340
rect 21308 11282 21364 11294
rect 21308 11230 21310 11282
rect 21362 11230 21364 11282
rect 21196 11172 21252 11182
rect 21308 11172 21364 11230
rect 21644 11282 21700 11294
rect 21644 11230 21646 11282
rect 21698 11230 21700 11282
rect 21252 11116 21588 11172
rect 21196 11106 21252 11116
rect 21532 10834 21588 11116
rect 21532 10782 21534 10834
rect 21586 10782 21588 10834
rect 21532 10770 21588 10782
rect 21644 10500 21700 11230
rect 22428 10834 22484 11340
rect 22540 11282 22596 12012
rect 22988 12002 23044 12012
rect 22540 11230 22542 11282
rect 22594 11230 22596 11282
rect 22540 11218 22596 11230
rect 23100 10948 23156 15486
rect 23884 15540 23940 16156
rect 23884 15446 23940 15484
rect 23996 17780 24052 17790
rect 23996 15652 24052 17724
rect 25116 17108 25172 23884
rect 25228 23828 25284 23838
rect 25228 23734 25284 23772
rect 25340 23604 25396 27804
rect 25452 26852 25508 26862
rect 25452 26758 25508 26796
rect 25676 26516 25732 27806
rect 25676 26450 25732 26460
rect 25900 26964 25956 27002
rect 25900 26514 25956 26908
rect 25900 26462 25902 26514
rect 25954 26462 25956 26514
rect 25900 26450 25956 26462
rect 26012 26514 26068 31836
rect 26460 31826 26516 31838
rect 26572 29540 26628 40348
rect 26908 40180 26964 40190
rect 26908 38274 26964 40124
rect 27020 39618 27076 41692
rect 27468 41636 27524 43148
rect 27916 42866 27972 43596
rect 28364 43538 28420 45164
rect 28588 44884 28644 45276
rect 28476 44828 28644 44884
rect 28476 44434 28532 44828
rect 28476 44382 28478 44434
rect 28530 44382 28532 44434
rect 28476 44370 28532 44382
rect 28364 43486 28366 43538
rect 28418 43486 28420 43538
rect 28364 43474 28420 43486
rect 27916 42814 27918 42866
rect 27970 42814 27972 42866
rect 27916 42802 27972 42814
rect 28140 42756 28196 42766
rect 28140 42662 28196 42700
rect 28476 42196 28532 42206
rect 27132 41580 27524 41636
rect 27692 41972 27748 41982
rect 27132 41298 27188 41580
rect 27132 41246 27134 41298
rect 27186 41246 27188 41298
rect 27132 41234 27188 41246
rect 27468 41300 27524 41310
rect 27524 41244 27636 41300
rect 27468 41206 27524 41244
rect 27580 40626 27636 41244
rect 27580 40574 27582 40626
rect 27634 40574 27636 40626
rect 27580 40562 27636 40574
rect 27020 39566 27022 39618
rect 27074 39566 27076 39618
rect 27020 39554 27076 39566
rect 27132 40290 27188 40302
rect 27132 40238 27134 40290
rect 27186 40238 27188 40290
rect 27132 39284 27188 40238
rect 27468 39508 27524 39518
rect 27468 39414 27524 39452
rect 27132 39218 27188 39228
rect 27244 38836 27300 38846
rect 27244 38742 27300 38780
rect 27692 38668 27748 41916
rect 27804 41858 27860 41870
rect 27804 41806 27806 41858
rect 27858 41806 27860 41858
rect 27804 40628 27860 41806
rect 28252 41860 28308 41870
rect 28252 41766 28308 41804
rect 28364 41412 28420 41422
rect 28364 41298 28420 41356
rect 28364 41246 28366 41298
rect 28418 41246 28420 41298
rect 28364 41234 28420 41246
rect 28140 41076 28196 41086
rect 27916 40964 27972 40974
rect 27916 40870 27972 40908
rect 27804 40562 27860 40572
rect 28028 40292 28084 40302
rect 28140 40292 28196 41020
rect 28476 40626 28532 42140
rect 28476 40574 28478 40626
rect 28530 40574 28532 40626
rect 28476 40562 28532 40574
rect 28028 40290 28196 40292
rect 28028 40238 28030 40290
rect 28082 40238 28196 40290
rect 28028 40236 28196 40238
rect 28588 40292 28644 40302
rect 28028 40226 28084 40236
rect 28476 39396 28532 39406
rect 28588 39396 28644 40236
rect 28476 39394 28644 39396
rect 28476 39342 28478 39394
rect 28530 39342 28644 39394
rect 28476 39340 28644 39342
rect 28476 39330 28532 39340
rect 26908 38222 26910 38274
rect 26962 38222 26964 38274
rect 26908 38210 26964 38222
rect 27468 38612 27748 38668
rect 28028 38722 28084 38734
rect 28028 38670 28030 38722
rect 28082 38670 28084 38722
rect 28028 38668 28084 38670
rect 28028 38612 28308 38668
rect 26908 37828 26964 37838
rect 26908 37734 26964 37772
rect 27132 37380 27188 37390
rect 26684 35812 26740 35822
rect 26684 35308 26740 35756
rect 27020 35698 27076 35710
rect 27020 35646 27022 35698
rect 27074 35646 27076 35698
rect 26684 35252 26964 35308
rect 26684 34916 26740 34926
rect 26684 31948 26740 34860
rect 26908 34356 26964 35252
rect 27020 34692 27076 35646
rect 27020 34626 27076 34636
rect 27020 34356 27076 34366
rect 26908 34354 27076 34356
rect 26908 34302 27022 34354
rect 27074 34302 27076 34354
rect 26908 34300 27076 34302
rect 27020 34290 27076 34300
rect 26796 33572 26852 33582
rect 27020 33572 27076 33582
rect 27132 33572 27188 37324
rect 27356 35476 27412 35486
rect 27356 34242 27412 35420
rect 27356 34190 27358 34242
rect 27410 34190 27412 34242
rect 27356 34178 27412 34190
rect 26796 33570 27132 33572
rect 26796 33518 26798 33570
rect 26850 33518 27022 33570
rect 27074 33518 27132 33570
rect 26796 33516 27132 33518
rect 26796 33458 26852 33516
rect 27020 33478 27076 33516
rect 27132 33478 27188 33516
rect 26796 33406 26798 33458
rect 26850 33406 26852 33458
rect 26796 33394 26852 33406
rect 27356 33346 27412 33358
rect 27356 33294 27358 33346
rect 27410 33294 27412 33346
rect 27356 33236 27412 33294
rect 27356 33170 27412 33180
rect 27132 33124 27188 33134
rect 27132 33030 27188 33068
rect 26908 32562 26964 32574
rect 26908 32510 26910 32562
rect 26962 32510 26964 32562
rect 26908 32004 26964 32510
rect 27468 32452 27524 38612
rect 28252 37490 28308 38612
rect 28252 37438 28254 37490
rect 28306 37438 28308 37490
rect 28252 37426 28308 37438
rect 27804 37380 27860 37390
rect 28140 37380 28196 37390
rect 27804 37378 28140 37380
rect 27804 37326 27806 37378
rect 27858 37326 28140 37378
rect 27804 37324 28140 37326
rect 27804 37314 27860 37324
rect 28140 37286 28196 37324
rect 28476 37266 28532 37278
rect 28476 37214 28478 37266
rect 28530 37214 28532 37266
rect 28140 36594 28196 36606
rect 28140 36542 28142 36594
rect 28194 36542 28196 36594
rect 28140 35924 28196 36542
rect 28140 35858 28196 35868
rect 28364 36260 28420 36270
rect 28252 35698 28308 35710
rect 28252 35646 28254 35698
rect 28306 35646 28308 35698
rect 28252 34692 28308 35646
rect 28252 34626 28308 34636
rect 28140 34132 28196 34142
rect 27692 33572 27748 33582
rect 27692 33478 27748 33516
rect 28028 33348 28084 33358
rect 28028 33254 28084 33292
rect 27804 33122 27860 33134
rect 27804 33070 27806 33122
rect 27858 33070 27860 33122
rect 27804 32788 27860 33070
rect 27580 32732 27860 32788
rect 27580 32674 27636 32732
rect 27580 32622 27582 32674
rect 27634 32622 27636 32674
rect 27580 32610 27636 32622
rect 27468 32396 27748 32452
rect 26684 31892 26964 31948
rect 26684 31780 26740 31892
rect 26684 31714 26740 31724
rect 26908 31668 26964 31678
rect 26908 30212 26964 31612
rect 26908 30210 27188 30212
rect 26908 30158 26910 30210
rect 26962 30158 27188 30210
rect 26908 30156 27188 30158
rect 26908 30146 26964 30156
rect 26572 29474 26628 29484
rect 26348 29428 26404 29438
rect 26236 29316 26292 29326
rect 26348 29316 26404 29372
rect 26684 29428 26740 29438
rect 27020 29428 27076 29438
rect 26684 29334 26740 29372
rect 26908 29426 27076 29428
rect 26908 29374 27022 29426
rect 27074 29374 27076 29426
rect 26908 29372 27076 29374
rect 26236 29314 26404 29316
rect 26236 29262 26238 29314
rect 26290 29262 26404 29314
rect 26236 29260 26404 29262
rect 26236 29250 26292 29260
rect 26348 27858 26404 29260
rect 26796 29204 26852 29214
rect 26684 29148 26796 29204
rect 26348 27806 26350 27858
rect 26402 27806 26404 27858
rect 26348 27412 26404 27806
rect 26572 27858 26628 27870
rect 26572 27806 26574 27858
rect 26626 27806 26628 27858
rect 26348 27356 26516 27412
rect 26460 27074 26516 27356
rect 26460 27022 26462 27074
rect 26514 27022 26516 27074
rect 26348 26962 26404 26974
rect 26348 26910 26350 26962
rect 26402 26910 26404 26962
rect 26012 26462 26014 26514
rect 26066 26462 26068 26514
rect 26012 26450 26068 26462
rect 26124 26740 26180 26750
rect 25452 26292 25508 26302
rect 25452 26198 25508 26236
rect 25676 26292 25732 26302
rect 25676 26290 26068 26292
rect 25676 26238 25678 26290
rect 25730 26238 26068 26290
rect 25676 26236 26068 26238
rect 25676 26226 25732 26236
rect 25900 26068 25956 26078
rect 25900 25618 25956 26012
rect 25900 25566 25902 25618
rect 25954 25566 25956 25618
rect 25900 25554 25956 25566
rect 25676 25508 25732 25518
rect 25676 24946 25732 25452
rect 25676 24894 25678 24946
rect 25730 24894 25732 24946
rect 25676 24882 25732 24894
rect 26012 24052 26068 26236
rect 26124 25396 26180 26684
rect 26348 26404 26404 26910
rect 26348 26338 26404 26348
rect 26460 26292 26516 27022
rect 26572 26740 26628 27806
rect 26684 27746 26740 29148
rect 26796 29138 26852 29148
rect 26908 28756 26964 29372
rect 27020 29362 27076 29372
rect 27132 29092 27188 30156
rect 27244 29652 27300 29662
rect 27244 29558 27300 29596
rect 27356 29316 27412 29326
rect 27580 29316 27636 29326
rect 27356 29314 27636 29316
rect 27356 29262 27358 29314
rect 27410 29262 27582 29314
rect 27634 29262 27636 29314
rect 27356 29260 27636 29262
rect 27356 29250 27412 29260
rect 27580 29250 27636 29260
rect 27132 29036 27524 29092
rect 27468 28868 27524 29036
rect 27468 28774 27524 28812
rect 27244 28756 27300 28766
rect 26908 28754 27300 28756
rect 26908 28702 26910 28754
rect 26962 28702 27246 28754
rect 27298 28702 27300 28754
rect 26908 28700 27300 28702
rect 26908 28690 26964 28700
rect 27244 28690 27300 28700
rect 26796 28532 26852 28542
rect 26796 28084 26852 28476
rect 27468 28196 27524 28206
rect 26796 28082 26964 28084
rect 26796 28030 26798 28082
rect 26850 28030 26964 28082
rect 26796 28028 26964 28030
rect 26796 28018 26852 28028
rect 26684 27694 26686 27746
rect 26738 27694 26740 27746
rect 26684 27682 26740 27694
rect 26908 27186 26964 28028
rect 27468 27858 27524 28140
rect 27468 27806 27470 27858
rect 27522 27806 27524 27858
rect 27468 27524 27524 27806
rect 27692 27748 27748 32396
rect 28140 29650 28196 34076
rect 28364 33236 28420 36204
rect 28476 35700 28532 37214
rect 28476 35138 28532 35644
rect 28476 35086 28478 35138
rect 28530 35086 28532 35138
rect 28476 35074 28532 35086
rect 28588 36258 28644 36270
rect 28588 36206 28590 36258
rect 28642 36206 28644 36258
rect 28588 35028 28644 36206
rect 28700 35922 28756 58604
rect 28812 57540 28868 57550
rect 29036 57540 29092 61404
rect 29148 61394 29204 61404
rect 29148 60900 29204 60910
rect 29148 60786 29204 60844
rect 29148 60734 29150 60786
rect 29202 60734 29204 60786
rect 29148 60722 29204 60734
rect 29148 60562 29204 60574
rect 29148 60510 29150 60562
rect 29202 60510 29204 60562
rect 29148 60004 29204 60510
rect 29148 59938 29204 59948
rect 28812 57538 29092 57540
rect 28812 57486 28814 57538
rect 28866 57486 29092 57538
rect 28812 57484 29092 57486
rect 29260 59892 29316 59902
rect 29372 59892 29428 61628
rect 29260 59890 29428 59892
rect 29260 59838 29262 59890
rect 29314 59838 29428 59890
rect 29260 59836 29428 59838
rect 29484 61572 29540 61582
rect 29932 61572 29988 61964
rect 30156 61908 30212 64092
rect 30268 62188 30324 65996
rect 30380 65986 30436 65996
rect 30380 64036 30436 64046
rect 30492 64036 30548 66332
rect 30716 66164 30772 66174
rect 30716 66070 30772 66108
rect 30828 65940 30884 70028
rect 30940 69748 30996 69758
rect 30940 68850 30996 69692
rect 30940 68798 30942 68850
rect 30994 68798 30996 68850
rect 30940 68786 30996 68798
rect 30940 66946 30996 66958
rect 30940 66894 30942 66946
rect 30994 66894 30996 66946
rect 30940 66836 30996 66894
rect 30940 66164 30996 66780
rect 30940 66098 30996 66108
rect 30716 65884 30884 65940
rect 30604 65492 30660 65502
rect 30604 65398 30660 65436
rect 30380 64034 30660 64036
rect 30380 63982 30382 64034
rect 30434 63982 30660 64034
rect 30380 63980 30660 63982
rect 30380 63970 30436 63980
rect 30604 63138 30660 63980
rect 30716 63362 30772 65884
rect 30940 65604 30996 65614
rect 30940 65510 30996 65548
rect 30828 64484 30884 64494
rect 30828 63922 30884 64428
rect 30940 64036 30996 64046
rect 31052 64036 31108 70588
rect 31164 70196 31220 70206
rect 31164 70102 31220 70140
rect 31164 68964 31220 68974
rect 31164 67844 31220 68908
rect 31276 68068 31332 70924
rect 31612 70588 31668 75404
rect 31724 75516 31836 75572
rect 31724 75124 31780 75516
rect 31836 75506 31892 75516
rect 32172 75572 32228 75582
rect 32396 75572 32452 75582
rect 32172 75570 32340 75572
rect 32172 75518 32174 75570
rect 32226 75518 32340 75570
rect 32172 75516 32340 75518
rect 32172 75506 32228 75516
rect 32284 75348 32340 75516
rect 32396 75478 32452 75516
rect 33292 75348 33348 75854
rect 32284 75292 32900 75348
rect 31724 75030 31780 75068
rect 31836 75236 31892 75246
rect 32844 75236 32900 75292
rect 33292 75282 33348 75292
rect 33404 76244 33460 76254
rect 32844 75180 33124 75236
rect 31388 70532 31668 70588
rect 31724 70978 31780 70990
rect 31724 70926 31726 70978
rect 31778 70926 31780 70978
rect 31724 70756 31780 70926
rect 31388 69524 31444 70532
rect 31724 69636 31780 70700
rect 31836 70420 31892 75180
rect 32508 75124 32564 75134
rect 31948 73892 32004 73902
rect 31948 72660 32004 73836
rect 31948 72658 32452 72660
rect 31948 72606 31950 72658
rect 32002 72606 32452 72658
rect 31948 72604 32452 72606
rect 31948 72594 32004 72604
rect 31836 70354 31892 70364
rect 32172 72100 32228 72110
rect 31836 70196 31892 70206
rect 31836 70102 31892 70140
rect 32172 70194 32228 72044
rect 32396 71988 32452 72604
rect 32396 71894 32452 71932
rect 32508 71204 32564 75068
rect 33068 75122 33124 75180
rect 33068 75070 33070 75122
rect 33122 75070 33124 75122
rect 33068 75058 33124 75070
rect 33404 75010 33460 76188
rect 33516 75572 33572 75582
rect 33516 75478 33572 75516
rect 33628 75124 33684 76636
rect 34412 76580 34468 77196
rect 34748 77476 34804 77486
rect 35084 77476 35140 77756
rect 35644 77700 35700 78542
rect 35868 78596 35924 78606
rect 35868 78502 35924 78540
rect 35980 78594 36036 78606
rect 35980 78542 35982 78594
rect 36034 78542 36036 78594
rect 35756 78148 35812 78158
rect 35756 77812 35812 78092
rect 35868 78036 35924 78046
rect 35868 77942 35924 77980
rect 35756 77756 35924 77812
rect 35196 77644 35460 77654
rect 35644 77644 35812 77700
rect 35252 77588 35300 77644
rect 35356 77588 35404 77644
rect 35196 77578 35460 77588
rect 35756 77588 35812 77644
rect 35196 77476 35252 77486
rect 35084 77474 35252 77476
rect 35084 77422 35198 77474
rect 35250 77422 35252 77474
rect 35084 77420 35252 77422
rect 34748 77250 34804 77420
rect 35196 77410 35252 77420
rect 34748 77198 34750 77250
rect 34802 77198 34804 77250
rect 34748 77186 34804 77198
rect 35420 77362 35476 77374
rect 35420 77310 35422 77362
rect 35474 77310 35476 77362
rect 34524 77140 34580 77150
rect 34524 77138 34692 77140
rect 34524 77086 34526 77138
rect 34578 77086 34692 77138
rect 34524 77084 34692 77086
rect 34524 77074 34580 77084
rect 34636 76580 34692 77084
rect 35420 77028 35476 77310
rect 35644 77364 35700 77374
rect 35644 77270 35700 77308
rect 35756 77250 35812 77532
rect 35756 77198 35758 77250
rect 35810 77198 35812 77250
rect 35756 77186 35812 77198
rect 35420 76962 35476 76972
rect 35420 76804 35476 76814
rect 34636 76524 34916 76580
rect 34412 76514 34468 76524
rect 33964 76468 34020 76478
rect 33964 76374 34020 76412
rect 34748 76356 34804 76366
rect 34636 76354 34804 76356
rect 34636 76302 34750 76354
rect 34802 76302 34804 76354
rect 34636 76300 34804 76302
rect 34188 76244 34244 76254
rect 34188 76150 34244 76188
rect 34524 76244 34580 76254
rect 34524 76150 34580 76188
rect 34076 75908 34132 75918
rect 34076 75814 34132 75852
rect 34636 75796 34692 76300
rect 34748 76290 34804 76300
rect 34524 75740 34692 75796
rect 34412 75684 34468 75694
rect 33964 75628 34412 75684
rect 33964 75570 34020 75628
rect 33964 75518 33966 75570
rect 34018 75518 34020 75570
rect 33964 75506 34020 75518
rect 33740 75460 33796 75470
rect 33740 75366 33796 75404
rect 33964 75348 34020 75358
rect 33740 75124 33796 75134
rect 33964 75124 34020 75292
rect 33404 74958 33406 75010
rect 33458 74958 33460 75010
rect 33404 74946 33460 74958
rect 33516 75122 33796 75124
rect 33516 75070 33742 75122
rect 33794 75070 33796 75122
rect 33516 75068 33796 75070
rect 32508 71090 32564 71148
rect 32508 71038 32510 71090
rect 32562 71038 32564 71090
rect 32508 71026 32564 71038
rect 32732 74788 32788 74798
rect 32732 74116 32788 74732
rect 32732 70980 32788 74060
rect 33516 74002 33572 75068
rect 33740 75058 33796 75068
rect 33852 75122 34020 75124
rect 33852 75070 33966 75122
rect 34018 75070 34020 75122
rect 33852 75068 34020 75070
rect 33740 74116 33796 74126
rect 33852 74116 33908 75068
rect 33964 75058 34020 75068
rect 34076 75124 34132 75134
rect 34076 75010 34132 75068
rect 34076 74958 34078 75010
rect 34130 74958 34132 75010
rect 34076 74946 34132 74958
rect 34412 74900 34468 75628
rect 34524 75682 34580 75740
rect 34860 75684 34916 76524
rect 35308 76468 35364 76478
rect 35084 76412 35308 76468
rect 35420 76468 35476 76748
rect 35868 76578 35924 77756
rect 35980 77474 36036 78542
rect 36092 78594 36148 78606
rect 36092 78542 36094 78594
rect 36146 78542 36148 78594
rect 36092 78484 36148 78542
rect 37996 78596 38052 78606
rect 36092 78428 36596 78484
rect 36540 78036 36596 78428
rect 37324 78260 37380 78270
rect 37100 78148 37156 78158
rect 37100 78054 37156 78092
rect 36764 78036 36820 78046
rect 36540 78034 36820 78036
rect 36540 77982 36766 78034
rect 36818 77982 36820 78034
rect 36540 77980 36820 77982
rect 35980 77422 35982 77474
rect 36034 77422 36036 77474
rect 35980 77410 36036 77422
rect 36092 77924 36148 77934
rect 36092 76804 36148 77868
rect 36316 77924 36372 77934
rect 36316 77830 36372 77868
rect 36204 77810 36260 77822
rect 36204 77758 36206 77810
rect 36258 77758 36260 77810
rect 36204 77476 36260 77758
rect 36540 77812 36596 77822
rect 36540 77718 36596 77756
rect 36204 77410 36260 77420
rect 36652 77476 36708 77486
rect 36428 77252 36484 77262
rect 36428 77158 36484 77196
rect 36316 77138 36372 77150
rect 36316 77086 36318 77138
rect 36370 77086 36372 77138
rect 36316 76916 36372 77086
rect 36316 76860 36484 76916
rect 36428 76804 36484 76860
rect 36092 76748 36260 76804
rect 35868 76526 35870 76578
rect 35922 76526 35924 76578
rect 35644 76468 35700 76478
rect 35420 76466 35700 76468
rect 35420 76414 35646 76466
rect 35698 76414 35700 76466
rect 35420 76412 35700 76414
rect 35084 75908 35140 76412
rect 35308 76374 35364 76412
rect 35644 76402 35700 76412
rect 35532 76244 35588 76254
rect 35196 76076 35460 76086
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35196 76010 35460 76020
rect 35084 75852 35476 75908
rect 34524 75630 34526 75682
rect 34578 75630 34580 75682
rect 34524 75618 34580 75630
rect 34748 75628 34916 75684
rect 35196 75682 35252 75694
rect 35196 75630 35198 75682
rect 35250 75630 35252 75682
rect 34636 75570 34692 75582
rect 34636 75518 34638 75570
rect 34690 75518 34692 75570
rect 34636 75460 34692 75518
rect 34636 75012 34692 75404
rect 34636 74946 34692 74956
rect 34748 74900 34804 75628
rect 34972 75572 35028 75582
rect 35028 75516 35140 75572
rect 34972 75478 35028 75516
rect 34972 75012 35028 75022
rect 34412 74844 34580 74900
rect 34412 74676 34468 74686
rect 34076 74674 34468 74676
rect 34076 74622 34414 74674
rect 34466 74622 34468 74674
rect 34076 74620 34468 74622
rect 33740 74114 33908 74116
rect 33740 74062 33742 74114
rect 33794 74062 33908 74114
rect 33740 74060 33908 74062
rect 33964 74116 34020 74126
rect 34076 74116 34132 74620
rect 34412 74610 34468 74620
rect 33964 74114 34132 74116
rect 33964 74062 33966 74114
rect 34018 74062 34132 74114
rect 33964 74060 34132 74062
rect 33740 74050 33796 74060
rect 33964 74050 34020 74060
rect 33516 73950 33518 74002
rect 33570 73950 33572 74002
rect 33516 73938 33572 73950
rect 34524 73948 34580 74844
rect 34748 74898 34916 74900
rect 34748 74846 34750 74898
rect 34802 74846 34916 74898
rect 34748 74844 34916 74846
rect 34748 74834 34804 74844
rect 34860 74116 34916 74844
rect 34972 74898 35028 74956
rect 34972 74846 34974 74898
rect 35026 74846 35028 74898
rect 34972 74834 35028 74846
rect 35084 74340 35140 75516
rect 35196 75124 35252 75630
rect 35308 75682 35364 75694
rect 35308 75630 35310 75682
rect 35362 75630 35364 75682
rect 35308 75460 35364 75630
rect 35308 75394 35364 75404
rect 35308 75124 35364 75134
rect 35252 75122 35364 75124
rect 35252 75070 35310 75122
rect 35362 75070 35364 75122
rect 35252 75068 35364 75070
rect 35196 75030 35252 75068
rect 35308 75058 35364 75068
rect 35420 75010 35476 75852
rect 35532 75794 35588 76188
rect 35532 75742 35534 75794
rect 35586 75742 35588 75794
rect 35532 75730 35588 75742
rect 35420 74958 35422 75010
rect 35474 74958 35476 75010
rect 35420 74946 35476 74958
rect 35644 75570 35700 75582
rect 35644 75518 35646 75570
rect 35698 75518 35700 75570
rect 35644 74788 35700 75518
rect 35868 75458 35924 76526
rect 36092 76580 36148 76590
rect 36092 75684 36148 76524
rect 36092 75590 36148 75628
rect 36204 76580 36260 76748
rect 36428 76738 36484 76748
rect 36316 76580 36372 76590
rect 36204 76524 36316 76580
rect 36204 75682 36260 76524
rect 36316 76514 36372 76524
rect 36428 76578 36484 76590
rect 36428 76526 36430 76578
rect 36482 76526 36484 76578
rect 36204 75630 36206 75682
rect 36258 75630 36260 75682
rect 35868 75406 35870 75458
rect 35922 75406 35924 75458
rect 35868 75348 35924 75406
rect 36092 75460 36148 75470
rect 35980 75348 36036 75358
rect 35868 75292 35980 75348
rect 35980 75282 36036 75292
rect 35980 75124 36036 75134
rect 35756 74788 35812 74798
rect 35644 74786 35812 74788
rect 35644 74734 35758 74786
rect 35810 74734 35812 74786
rect 35644 74732 35812 74734
rect 35756 74676 35812 74732
rect 35756 74610 35812 74620
rect 35980 74674 36036 75068
rect 35980 74622 35982 74674
rect 36034 74622 36036 74674
rect 35196 74508 35460 74518
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35196 74442 35460 74452
rect 35308 74340 35364 74350
rect 35084 74284 35308 74340
rect 34972 74116 35028 74126
rect 34860 74114 35028 74116
rect 34860 74062 34974 74114
rect 35026 74062 35028 74114
rect 34860 74060 35028 74062
rect 34972 74050 35028 74060
rect 35308 74114 35364 74284
rect 35756 74340 35812 74350
rect 35756 74246 35812 74284
rect 35308 74062 35310 74114
rect 35362 74062 35364 74114
rect 35308 74050 35364 74062
rect 35420 74116 35476 74126
rect 35196 74002 35252 74014
rect 35196 73950 35198 74002
rect 35250 73950 35252 74002
rect 35196 73948 35252 73950
rect 35420 73948 35476 74060
rect 35644 74116 35700 74126
rect 35980 74116 36036 74622
rect 35644 74114 36036 74116
rect 35644 74062 35646 74114
rect 35698 74062 36036 74114
rect 35644 74060 36036 74062
rect 36092 74116 36148 75404
rect 36204 74338 36260 75630
rect 36428 76468 36484 76526
rect 36316 75124 36372 75134
rect 36316 75030 36372 75068
rect 36428 74676 36484 76412
rect 36652 75010 36708 77420
rect 36764 75122 36820 77980
rect 37212 78036 37268 78046
rect 37212 77476 37268 77980
rect 37212 77382 37268 77420
rect 36876 77252 36932 77262
rect 36876 76578 36932 77196
rect 37100 77252 37156 77262
rect 37324 77252 37380 78204
rect 37884 77476 37940 77486
rect 37884 77382 37940 77420
rect 37996 77362 38052 78540
rect 37996 77310 37998 77362
rect 38050 77310 38052 77362
rect 37996 77298 38052 77310
rect 37436 77252 37492 77262
rect 37100 77250 37268 77252
rect 37100 77198 37102 77250
rect 37154 77198 37268 77250
rect 37100 77196 37268 77198
rect 37100 77186 37156 77196
rect 36988 77140 37044 77150
rect 36988 76690 37044 77084
rect 37100 77028 37156 77038
rect 37100 76934 37156 76972
rect 37212 76804 37268 77196
rect 37212 76738 37268 76748
rect 37324 77196 37436 77252
rect 36988 76638 36990 76690
rect 37042 76638 37044 76690
rect 36988 76626 37044 76638
rect 36876 76526 36878 76578
rect 36930 76526 36932 76578
rect 36876 76514 36932 76526
rect 37100 76468 37156 76478
rect 37324 76468 37380 77196
rect 37436 77158 37492 77196
rect 38108 77252 38164 77262
rect 38108 77138 38164 77196
rect 38108 77086 38110 77138
rect 38162 77086 38164 77138
rect 38108 77074 38164 77086
rect 37660 76916 37716 76926
rect 37660 76690 37716 76860
rect 37660 76638 37662 76690
rect 37714 76638 37716 76690
rect 37660 76626 37716 76638
rect 37884 76580 37940 76590
rect 37884 76486 37940 76524
rect 37156 76412 37380 76468
rect 37436 76466 37492 76478
rect 37436 76414 37438 76466
rect 37490 76414 37492 76466
rect 37100 76374 37156 76412
rect 37436 76356 37492 76414
rect 37436 76290 37492 76300
rect 37996 76466 38052 76478
rect 37996 76414 37998 76466
rect 38050 76414 38052 76466
rect 37996 75908 38052 76414
rect 37996 75842 38052 75852
rect 37100 75796 37156 75806
rect 37100 75702 37156 75740
rect 37212 75684 37268 75694
rect 36988 75572 37044 75582
rect 36988 75478 37044 75516
rect 37212 75570 37268 75628
rect 37212 75518 37214 75570
rect 37266 75518 37268 75570
rect 36764 75070 36766 75122
rect 36818 75070 36820 75122
rect 36764 75058 36820 75070
rect 36652 74958 36654 75010
rect 36706 74958 36708 75010
rect 36652 74946 36708 74958
rect 37212 75010 37268 75518
rect 37436 75458 37492 75470
rect 37436 75406 37438 75458
rect 37490 75406 37492 75458
rect 37436 75124 37492 75406
rect 37436 75058 37492 75068
rect 37212 74958 37214 75010
rect 37266 74958 37268 75010
rect 37212 74946 37268 74958
rect 36428 74610 36484 74620
rect 36876 74898 36932 74910
rect 36876 74846 36878 74898
rect 36930 74846 36932 74898
rect 36876 74676 36932 74846
rect 38220 74900 38276 74910
rect 38276 74844 38388 74900
rect 38220 74806 38276 74844
rect 37660 74788 37716 74798
rect 37660 74694 37716 74732
rect 36876 74610 36932 74620
rect 36204 74286 36206 74338
rect 36258 74286 36260 74338
rect 36204 74274 36260 74286
rect 38332 74226 38388 74844
rect 38332 74174 38334 74226
rect 38386 74174 38388 74226
rect 38332 74162 38388 74174
rect 36316 74116 36372 74126
rect 36148 74114 36372 74116
rect 36148 74062 36318 74114
rect 36370 74062 36372 74114
rect 36148 74060 36372 74062
rect 35644 74050 35700 74060
rect 33852 73890 33908 73902
rect 34524 73892 35252 73948
rect 35308 73892 35476 73948
rect 35756 73892 35812 73902
rect 33852 73838 33854 73890
rect 33906 73838 33908 73890
rect 33628 72322 33684 72334
rect 33628 72270 33630 72322
rect 33682 72270 33684 72322
rect 33628 72212 33684 72270
rect 33292 72156 33628 72212
rect 33292 71876 33348 72156
rect 33628 72146 33684 72156
rect 33740 72324 33796 72334
rect 32732 70886 32788 70924
rect 33068 71874 33348 71876
rect 33068 71822 33294 71874
rect 33346 71822 33348 71874
rect 33068 71820 33348 71822
rect 32172 70142 32174 70194
rect 32226 70142 32228 70194
rect 32172 70130 32228 70142
rect 32284 70868 32340 70878
rect 32620 70868 32676 70878
rect 32340 70866 32676 70868
rect 32340 70814 32622 70866
rect 32674 70814 32676 70866
rect 32340 70812 32676 70814
rect 32172 69970 32228 69982
rect 32172 69918 32174 69970
rect 32226 69918 32228 69970
rect 31724 69580 32004 69636
rect 31388 69522 31556 69524
rect 31388 69470 31390 69522
rect 31442 69470 31556 69522
rect 31388 69468 31556 69470
rect 31388 69458 31444 69468
rect 31500 69412 31556 69468
rect 31836 69412 31892 69422
rect 31500 69410 31892 69412
rect 31500 69358 31838 69410
rect 31890 69358 31892 69410
rect 31500 69356 31892 69358
rect 31836 69346 31892 69356
rect 31948 69188 32004 69580
rect 32172 69634 32228 69918
rect 32172 69582 32174 69634
rect 32226 69582 32228 69634
rect 32172 69570 32228 69582
rect 32284 69412 32340 70812
rect 32620 70802 32676 70812
rect 33068 70194 33124 71820
rect 33292 71810 33348 71820
rect 33740 71988 33796 72268
rect 33852 72100 33908 73838
rect 33852 72034 33908 72044
rect 34076 73556 34132 73566
rect 34076 72322 34132 73500
rect 34972 72436 35028 73892
rect 35308 73780 35364 73892
rect 35084 73724 35364 73780
rect 35084 72658 35140 73724
rect 35196 72940 35460 72950
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35196 72874 35460 72884
rect 35084 72606 35086 72658
rect 35138 72606 35140 72658
rect 35084 72594 35140 72606
rect 34972 72380 35140 72436
rect 34076 72270 34078 72322
rect 34130 72270 34132 72322
rect 34076 72212 34132 72270
rect 34076 71988 34132 72156
rect 34636 72322 34692 72334
rect 34636 72270 34638 72322
rect 34690 72270 34692 72322
rect 34076 71932 34356 71988
rect 33068 70142 33070 70194
rect 33122 70142 33124 70194
rect 33068 69748 33124 70142
rect 33292 71540 33348 71550
rect 33292 70194 33348 71484
rect 33404 71538 33460 71550
rect 33404 71486 33406 71538
rect 33458 71486 33460 71538
rect 33404 70868 33460 71486
rect 33404 70802 33460 70812
rect 33628 71204 33684 71214
rect 33628 70418 33684 71148
rect 33740 70978 33796 71932
rect 34300 71876 34356 71932
rect 34412 71876 34468 71886
rect 34300 71820 34412 71876
rect 34412 71782 34468 71820
rect 34188 71762 34244 71774
rect 34188 71710 34190 71762
rect 34242 71710 34244 71762
rect 33740 70926 33742 70978
rect 33794 70926 33796 70978
rect 33740 70914 33796 70926
rect 33964 71650 34020 71662
rect 33964 71598 33966 71650
rect 34018 71598 34020 71650
rect 33628 70366 33630 70418
rect 33682 70366 33684 70418
rect 33628 70354 33684 70366
rect 33292 70142 33294 70194
rect 33346 70142 33348 70194
rect 33292 70130 33348 70142
rect 33516 70194 33572 70206
rect 33516 70142 33518 70194
rect 33570 70142 33572 70194
rect 33404 69972 33460 69982
rect 33068 69682 33124 69692
rect 33292 69916 33404 69972
rect 32956 69522 33012 69534
rect 32956 69470 32958 69522
rect 33010 69470 33012 69522
rect 32844 69412 32900 69422
rect 31724 69132 32004 69188
rect 32060 69186 32116 69198
rect 32060 69134 32062 69186
rect 32114 69134 32116 69186
rect 31612 68626 31668 68638
rect 31612 68574 31614 68626
rect 31666 68574 31668 68626
rect 31276 68012 31556 68068
rect 31276 67844 31332 67854
rect 31164 67842 31332 67844
rect 31164 67790 31278 67842
rect 31330 67790 31332 67842
rect 31164 67788 31332 67790
rect 31276 67778 31332 67788
rect 31164 67172 31220 67182
rect 31164 66386 31220 67116
rect 31388 66948 31444 66958
rect 31164 66334 31166 66386
rect 31218 66334 31220 66386
rect 31164 66052 31220 66334
rect 31164 65986 31220 65996
rect 31276 66946 31444 66948
rect 31276 66894 31390 66946
rect 31442 66894 31444 66946
rect 31276 66892 31444 66894
rect 31276 66164 31332 66892
rect 31388 66882 31444 66892
rect 30940 64034 31108 64036
rect 30940 63982 30942 64034
rect 30994 63982 31108 64034
rect 30940 63980 31108 63982
rect 31164 64708 31220 64718
rect 31276 64708 31332 66108
rect 31164 64706 31332 64708
rect 31164 64654 31166 64706
rect 31218 64654 31332 64706
rect 31164 64652 31332 64654
rect 31388 65380 31444 65390
rect 30940 63970 30996 63980
rect 30828 63870 30830 63922
rect 30882 63870 30884 63922
rect 30828 63858 30884 63870
rect 30716 63310 30718 63362
rect 30770 63310 30772 63362
rect 30716 63298 30772 63310
rect 30828 63700 30884 63710
rect 30604 63086 30606 63138
rect 30658 63086 30660 63138
rect 30492 62580 30548 62590
rect 30492 62486 30548 62524
rect 30604 62188 30660 63086
rect 30828 63138 30884 63644
rect 30828 63086 30830 63138
rect 30882 63086 30884 63138
rect 30828 63074 30884 63086
rect 31052 62242 31108 62254
rect 31052 62190 31054 62242
rect 31106 62190 31108 62242
rect 30268 62132 30436 62188
rect 30604 62132 30996 62188
rect 30156 61842 30212 61852
rect 29484 61570 29988 61572
rect 29484 61518 29486 61570
rect 29538 61518 29988 61570
rect 29484 61516 29988 61518
rect 29484 60900 29540 61516
rect 29260 59780 29316 59836
rect 29484 59780 29540 60844
rect 29596 60786 29652 60798
rect 29596 60734 29598 60786
rect 29650 60734 29652 60786
rect 29596 60226 29652 60734
rect 29596 60174 29598 60226
rect 29650 60174 29652 60226
rect 29596 60162 29652 60174
rect 29596 60002 29652 60014
rect 29596 59950 29598 60002
rect 29650 59950 29652 60002
rect 29596 59780 29652 59950
rect 29932 60004 29988 60014
rect 30268 60004 30324 60014
rect 29932 59910 29988 59948
rect 30156 59948 30268 60004
rect 28812 57474 28868 57484
rect 29148 56868 29204 56878
rect 29148 56774 29204 56812
rect 29148 55298 29204 55310
rect 29148 55246 29150 55298
rect 29202 55246 29204 55298
rect 28812 54516 28868 54526
rect 28812 54422 28868 54460
rect 29148 54516 29204 55246
rect 29148 54450 29204 54460
rect 28924 53732 28980 53742
rect 28812 48804 28868 48814
rect 28812 46564 28868 48748
rect 28812 46498 28868 46508
rect 28924 43204 28980 53676
rect 29148 53730 29204 53742
rect 29148 53678 29150 53730
rect 29202 53678 29204 53730
rect 29148 52836 29204 53678
rect 29148 52770 29204 52780
rect 29260 50428 29316 59724
rect 29372 59724 29596 59780
rect 29372 58434 29428 59724
rect 29596 59714 29652 59724
rect 30156 59780 30212 59948
rect 30268 59938 30324 59948
rect 29820 59444 29876 59454
rect 29820 59350 29876 59388
rect 29484 59220 29540 59230
rect 29484 58658 29540 59164
rect 29484 58606 29486 58658
rect 29538 58606 29540 58658
rect 29484 58594 29540 58606
rect 29708 59218 29764 59230
rect 29708 59166 29710 59218
rect 29762 59166 29764 59218
rect 29372 58382 29374 58434
rect 29426 58382 29428 58434
rect 29372 58370 29428 58382
rect 29484 58212 29540 58222
rect 29484 58118 29540 58156
rect 29708 57316 29764 59166
rect 29708 57250 29764 57260
rect 29820 58324 29876 58334
rect 29932 58324 29988 58334
rect 29876 58322 29988 58324
rect 29876 58270 29934 58322
rect 29986 58270 29988 58322
rect 29876 58268 29988 58270
rect 29596 55970 29652 55982
rect 29596 55918 29598 55970
rect 29650 55918 29652 55970
rect 29372 55300 29428 55310
rect 29596 55300 29652 55918
rect 29372 55298 29652 55300
rect 29372 55246 29374 55298
rect 29426 55246 29652 55298
rect 29372 55244 29652 55246
rect 29372 54628 29428 55244
rect 29372 54562 29428 54572
rect 29148 50372 29316 50428
rect 29372 53844 29428 53854
rect 29372 52164 29428 53788
rect 29484 53732 29540 53742
rect 29820 53732 29876 58268
rect 29932 58258 29988 58268
rect 30156 58324 30212 59724
rect 30268 58548 30324 58558
rect 30268 58454 30324 58492
rect 30156 58322 30324 58324
rect 30156 58270 30158 58322
rect 30210 58270 30324 58322
rect 30156 58268 30324 58270
rect 30156 58258 30212 58268
rect 30156 56866 30212 56878
rect 30156 56814 30158 56866
rect 30210 56814 30212 56866
rect 30044 55972 30100 55982
rect 30156 55972 30212 56814
rect 30268 56754 30324 58268
rect 30380 57652 30436 62132
rect 30716 61908 30772 61918
rect 30492 61572 30548 61582
rect 30492 61478 30548 61516
rect 30492 60786 30548 60798
rect 30492 60734 30494 60786
rect 30546 60734 30548 60786
rect 30492 60004 30548 60734
rect 30492 59938 30548 59948
rect 30492 59220 30548 59230
rect 30492 59126 30548 59164
rect 30604 58548 30660 58558
rect 30604 58434 30660 58492
rect 30604 58382 30606 58434
rect 30658 58382 30660 58434
rect 30604 58370 30660 58382
rect 30604 57652 30660 57662
rect 30380 57650 30660 57652
rect 30380 57598 30606 57650
rect 30658 57598 30660 57650
rect 30380 57596 30660 57598
rect 30268 56702 30270 56754
rect 30322 56702 30324 56754
rect 30268 56690 30324 56702
rect 30380 57316 30436 57326
rect 29932 55970 30212 55972
rect 29932 55918 30046 55970
rect 30098 55918 30212 55970
rect 29932 55916 30212 55918
rect 29932 54068 29988 55916
rect 30044 55906 30100 55916
rect 30380 55522 30436 57260
rect 30604 56980 30660 57596
rect 30604 56914 30660 56924
rect 30716 56866 30772 61852
rect 30940 61458 30996 62132
rect 31052 61572 31108 62190
rect 31052 61506 31108 61516
rect 30940 61406 30942 61458
rect 30994 61406 30996 61458
rect 30828 60788 30884 60798
rect 30828 60694 30884 60732
rect 30940 59330 30996 61406
rect 30940 59278 30942 59330
rect 30994 59278 30996 59330
rect 30940 59266 30996 59278
rect 31052 57650 31108 57662
rect 31052 57598 31054 57650
rect 31106 57598 31108 57650
rect 30940 57316 30996 57326
rect 31052 57316 31108 57598
rect 30996 57260 31108 57316
rect 30940 57250 30996 57260
rect 30716 56814 30718 56866
rect 30770 56814 30772 56866
rect 30716 56802 30772 56814
rect 30940 56756 30996 56766
rect 30828 56754 30996 56756
rect 30828 56702 30942 56754
rect 30994 56702 30996 56754
rect 30828 56700 30996 56702
rect 30492 55972 30548 55982
rect 30828 55972 30884 56700
rect 30940 56690 30996 56700
rect 30940 56308 30996 56318
rect 30940 56214 30996 56252
rect 30492 55970 30884 55972
rect 30492 55918 30494 55970
rect 30546 55918 30884 55970
rect 30492 55916 30884 55918
rect 30492 55906 30548 55916
rect 30380 55470 30382 55522
rect 30434 55470 30436 55522
rect 30380 55458 30436 55470
rect 30044 54740 30100 54750
rect 30044 54646 30100 54684
rect 30156 54404 30212 54414
rect 30156 54310 30212 54348
rect 29932 54012 30212 54068
rect 29540 53676 29876 53732
rect 29484 53666 29540 53676
rect 29932 53620 29988 53630
rect 29708 53618 29988 53620
rect 29708 53566 29934 53618
rect 29986 53566 29988 53618
rect 29708 53564 29988 53566
rect 29372 52162 29652 52164
rect 29372 52110 29374 52162
rect 29426 52110 29652 52162
rect 29372 52108 29652 52110
rect 29036 46562 29092 46574
rect 29036 46510 29038 46562
rect 29090 46510 29092 46562
rect 29036 46116 29092 46510
rect 29036 46050 29092 46060
rect 29148 45892 29204 50372
rect 29260 48804 29316 48814
rect 29260 48710 29316 48748
rect 29372 48468 29428 52108
rect 29484 51938 29540 51950
rect 29484 51886 29486 51938
rect 29538 51886 29540 51938
rect 29484 50428 29540 51886
rect 29596 51940 29652 52108
rect 29708 52162 29764 53564
rect 29932 53554 29988 53564
rect 29708 52110 29710 52162
rect 29762 52110 29764 52162
rect 29708 52098 29764 52110
rect 30044 51940 30100 51950
rect 29596 51938 30100 51940
rect 29596 51886 30046 51938
rect 30098 51886 30100 51938
rect 29596 51884 30100 51886
rect 30044 51874 30100 51884
rect 30156 51492 30212 54012
rect 30492 53732 30548 53742
rect 30492 52162 30548 53676
rect 30492 52110 30494 52162
rect 30546 52110 30548 52162
rect 30492 52098 30548 52110
rect 30156 51436 30324 51492
rect 30156 51268 30212 51278
rect 29820 51266 30212 51268
rect 29820 51214 30158 51266
rect 30210 51214 30212 51266
rect 29820 51212 30212 51214
rect 29484 50372 29652 50428
rect 29372 48402 29428 48412
rect 29260 48132 29316 48142
rect 29260 48130 29540 48132
rect 29260 48078 29262 48130
rect 29314 48078 29540 48130
rect 29260 48076 29540 48078
rect 29260 48066 29316 48076
rect 29484 47346 29540 48076
rect 29596 47684 29652 50372
rect 29820 49700 29876 51212
rect 30156 51202 30212 51212
rect 30268 51044 30324 51436
rect 30380 51380 30436 51390
rect 30380 51286 30436 51324
rect 30156 50988 30324 51044
rect 29820 49698 30100 49700
rect 29820 49646 29822 49698
rect 29874 49646 30100 49698
rect 29820 49644 30100 49646
rect 29820 49634 29876 49644
rect 29708 49476 29764 49486
rect 29708 49138 29764 49420
rect 29708 49086 29710 49138
rect 29762 49086 29764 49138
rect 29708 49074 29764 49086
rect 30044 49026 30100 49644
rect 30044 48974 30046 49026
rect 30098 48974 30100 49026
rect 30044 48962 30100 48974
rect 29596 47628 29876 47684
rect 29708 47460 29764 47470
rect 29484 47294 29486 47346
rect 29538 47294 29540 47346
rect 29484 47282 29540 47294
rect 29596 47458 29764 47460
rect 29596 47406 29710 47458
rect 29762 47406 29764 47458
rect 29596 47404 29764 47406
rect 29596 46898 29652 47404
rect 29708 47394 29764 47404
rect 29596 46846 29598 46898
rect 29650 46846 29652 46898
rect 29596 46834 29652 46846
rect 29148 45836 29428 45892
rect 29036 45780 29092 45790
rect 29092 45724 29316 45780
rect 29036 45714 29092 45724
rect 29260 45666 29316 45724
rect 29260 45614 29262 45666
rect 29314 45614 29316 45666
rect 29260 45602 29316 45614
rect 29036 44660 29092 44670
rect 29036 43650 29092 44604
rect 29260 44212 29316 44222
rect 29260 44118 29316 44156
rect 29036 43598 29038 43650
rect 29090 43598 29092 43650
rect 29036 43586 29092 43598
rect 28924 43148 29092 43204
rect 28924 42308 28980 42318
rect 28924 41970 28980 42252
rect 28924 41918 28926 41970
rect 28978 41918 28980 41970
rect 28924 41906 28980 41918
rect 28700 35870 28702 35922
rect 28754 35870 28756 35922
rect 28700 35858 28756 35870
rect 28812 41858 28868 41870
rect 28812 41806 28814 41858
rect 28866 41806 28868 41858
rect 28588 34972 28756 35028
rect 28588 34802 28644 34814
rect 28588 34750 28590 34802
rect 28642 34750 28644 34802
rect 28476 34130 28532 34142
rect 28476 34078 28478 34130
rect 28530 34078 28532 34130
rect 28476 33460 28532 34078
rect 28588 33572 28644 34750
rect 28700 34580 28756 34972
rect 28700 34514 28756 34524
rect 28588 33506 28644 33516
rect 28476 33394 28532 33404
rect 28476 33236 28532 33246
rect 28420 33234 28532 33236
rect 28420 33182 28478 33234
rect 28530 33182 28532 33234
rect 28420 33180 28532 33182
rect 28364 33142 28420 33180
rect 28476 33170 28532 33180
rect 28812 33012 28868 41806
rect 29036 41410 29092 43148
rect 29036 41358 29038 41410
rect 29090 41358 29092 41410
rect 29036 41346 29092 41358
rect 29260 41748 29316 41758
rect 29260 41298 29316 41692
rect 29260 41246 29262 41298
rect 29314 41246 29316 41298
rect 29260 41234 29316 41246
rect 29148 40404 29204 40414
rect 29204 40348 29316 40404
rect 29148 40310 29204 40348
rect 29260 39732 29316 40348
rect 28924 39730 29316 39732
rect 28924 39678 29262 39730
rect 29314 39678 29316 39730
rect 28924 39676 29316 39678
rect 28924 37492 28980 39676
rect 29260 39666 29316 39676
rect 29372 38668 29428 45836
rect 29708 45668 29764 45678
rect 29484 45666 29764 45668
rect 29484 45614 29710 45666
rect 29762 45614 29764 45666
rect 29484 45612 29764 45614
rect 29484 43540 29540 45612
rect 29708 45602 29764 45612
rect 29708 44436 29764 44446
rect 29708 44342 29764 44380
rect 29484 43474 29540 43484
rect 29596 43428 29652 43438
rect 29596 43334 29652 43372
rect 29484 43092 29540 43102
rect 29484 42866 29540 43036
rect 29484 42814 29486 42866
rect 29538 42814 29540 42866
rect 29484 42084 29540 42814
rect 29708 42754 29764 42766
rect 29708 42702 29710 42754
rect 29762 42702 29764 42754
rect 29708 42308 29764 42702
rect 29708 42242 29764 42252
rect 29484 42082 29764 42084
rect 29484 42030 29486 42082
rect 29538 42030 29764 42082
rect 29484 42028 29764 42030
rect 29484 42018 29540 42028
rect 29484 41410 29540 41422
rect 29484 41358 29486 41410
rect 29538 41358 29540 41410
rect 29484 40626 29540 41358
rect 29708 41410 29764 42028
rect 29708 41358 29710 41410
rect 29762 41358 29764 41410
rect 29708 41298 29764 41358
rect 29708 41246 29710 41298
rect 29762 41246 29764 41298
rect 29708 41234 29764 41246
rect 29484 40574 29486 40626
rect 29538 40574 29540 40626
rect 29484 40562 29540 40574
rect 29596 40516 29652 40526
rect 29820 40516 29876 47628
rect 30156 46788 30212 50988
rect 30380 50932 30436 50942
rect 30268 49698 30324 49710
rect 30268 49646 30270 49698
rect 30322 49646 30324 49698
rect 30268 49476 30324 49646
rect 30268 49410 30324 49420
rect 30380 49252 30436 50876
rect 30604 50428 30660 55916
rect 31164 55412 31220 64652
rect 31388 64596 31444 65324
rect 31500 65156 31556 68012
rect 31612 65604 31668 68574
rect 31724 68180 31780 69132
rect 32060 68740 32116 69134
rect 32060 68674 32116 68684
rect 31948 68516 32004 68526
rect 31948 68422 32004 68460
rect 31836 68404 31892 68414
rect 31836 68310 31892 68348
rect 32284 68292 32340 69356
rect 32508 69410 32900 69412
rect 32508 69358 32846 69410
rect 32898 69358 32900 69410
rect 32508 69356 32900 69358
rect 31948 68236 32340 68292
rect 32396 68516 32452 68526
rect 31724 68124 31892 68180
rect 31724 67956 31780 67966
rect 31724 67862 31780 67900
rect 31724 67732 31780 67742
rect 31836 67732 31892 68124
rect 31948 68066 32004 68236
rect 31948 68014 31950 68066
rect 32002 68014 32004 68066
rect 31948 68002 32004 68014
rect 31724 67730 31892 67732
rect 31724 67678 31726 67730
rect 31778 67678 31892 67730
rect 31724 67676 31892 67678
rect 31724 67666 31780 67676
rect 32396 67172 32452 68460
rect 32508 67284 32564 69356
rect 32844 69346 32900 69356
rect 32956 68852 33012 69470
rect 32956 68786 33012 68796
rect 33180 68852 33236 68862
rect 33292 68852 33348 69916
rect 33404 69906 33460 69916
rect 33180 68850 33348 68852
rect 33180 68798 33182 68850
rect 33234 68798 33348 68850
rect 33180 68796 33348 68798
rect 33404 69298 33460 69310
rect 33404 69246 33406 69298
rect 33458 69246 33460 69298
rect 33180 68786 33236 68796
rect 33068 68740 33124 68750
rect 33068 68646 33124 68684
rect 32620 68628 32676 68638
rect 32620 68626 33012 68628
rect 32620 68574 32622 68626
rect 32674 68574 33012 68626
rect 32620 68572 33012 68574
rect 32620 68562 32676 68572
rect 32956 68068 33012 68572
rect 33404 68180 33460 69246
rect 33404 68114 33460 68124
rect 33068 68068 33124 68078
rect 32956 68012 33068 68068
rect 33068 67974 33124 68012
rect 32508 67218 32564 67228
rect 32956 67844 33012 67854
rect 32172 67116 32452 67172
rect 31836 66164 31892 66174
rect 31836 66070 31892 66108
rect 31612 65548 32004 65604
rect 31612 65380 31668 65390
rect 31612 65286 31668 65324
rect 31500 65100 31668 65156
rect 31276 63812 31332 63822
rect 31388 63812 31444 64540
rect 31276 63810 31444 63812
rect 31276 63758 31278 63810
rect 31330 63758 31444 63810
rect 31276 63756 31444 63758
rect 31276 60452 31332 63756
rect 31500 62132 31556 62142
rect 31500 60674 31556 62076
rect 31500 60622 31502 60674
rect 31554 60622 31556 60674
rect 31500 60610 31556 60622
rect 31276 60396 31556 60452
rect 31276 60002 31332 60014
rect 31276 59950 31278 60002
rect 31330 59950 31332 60002
rect 31276 59892 31332 59950
rect 31276 59826 31332 59836
rect 31276 59106 31332 59118
rect 31276 59054 31278 59106
rect 31330 59054 31332 59106
rect 31276 58324 31332 59054
rect 31276 58258 31332 58268
rect 31164 55298 31220 55356
rect 31164 55246 31166 55298
rect 31218 55246 31220 55298
rect 31164 55234 31220 55246
rect 31276 56866 31332 56878
rect 31276 56814 31278 56866
rect 31330 56814 31332 56866
rect 31276 54740 31332 56814
rect 31276 54674 31332 54684
rect 31164 53058 31220 53070
rect 31164 53006 31166 53058
rect 31218 53006 31220 53058
rect 30828 52948 30884 52958
rect 30716 52946 30884 52948
rect 30716 52894 30830 52946
rect 30882 52894 30884 52946
rect 30716 52892 30884 52894
rect 30716 51602 30772 52892
rect 30828 52882 30884 52892
rect 31164 52276 31220 53006
rect 31500 52836 31556 60396
rect 31612 59330 31668 65100
rect 31948 65044 32004 65548
rect 32172 65490 32228 67116
rect 32956 66498 33012 67788
rect 33180 67732 33236 67742
rect 33516 67732 33572 70142
rect 33740 70194 33796 70206
rect 33740 70142 33742 70194
rect 33794 70142 33796 70194
rect 33740 70084 33796 70142
rect 33964 70084 34020 71598
rect 34076 70420 34132 70430
rect 34076 70326 34132 70364
rect 33740 70028 34020 70084
rect 33740 68852 33796 68862
rect 33628 68516 33684 68526
rect 33628 67842 33684 68460
rect 33628 67790 33630 67842
rect 33682 67790 33684 67842
rect 33628 67778 33684 67790
rect 33740 67956 33796 68796
rect 33964 68626 34020 70028
rect 33964 68574 33966 68626
rect 34018 68574 34020 68626
rect 33964 68562 34020 68574
rect 32956 66446 32958 66498
rect 33010 66446 33012 66498
rect 32956 66434 33012 66446
rect 33068 67730 33572 67732
rect 33068 67678 33182 67730
rect 33234 67678 33572 67730
rect 33068 67676 33572 67678
rect 32172 65438 32174 65490
rect 32226 65438 32228 65490
rect 32172 65426 32228 65438
rect 32396 65602 32452 65614
rect 32396 65550 32398 65602
rect 32450 65550 32452 65602
rect 32396 65268 32452 65550
rect 32396 65202 32452 65212
rect 32508 65490 32564 65502
rect 32508 65438 32510 65490
rect 32562 65438 32564 65490
rect 31948 64988 32452 65044
rect 32060 64482 32116 64494
rect 32060 64430 32062 64482
rect 32114 64430 32116 64482
rect 31948 64260 32004 64270
rect 31948 64034 32004 64204
rect 32060 64146 32116 64430
rect 32060 64094 32062 64146
rect 32114 64094 32116 64146
rect 32060 64082 32116 64094
rect 32172 64482 32228 64494
rect 32172 64430 32174 64482
rect 32226 64430 32228 64482
rect 31948 63982 31950 64034
rect 32002 63982 32004 64034
rect 31948 63970 32004 63982
rect 32172 63364 32228 64430
rect 32284 64484 32340 64494
rect 32284 64390 32340 64428
rect 32284 64036 32340 64046
rect 32284 63942 32340 63980
rect 32172 63298 32228 63308
rect 32172 63138 32228 63150
rect 32172 63086 32174 63138
rect 32226 63086 32228 63138
rect 31724 62466 31780 62478
rect 31724 62414 31726 62466
rect 31778 62414 31780 62466
rect 31724 61684 31780 62414
rect 31724 61618 31780 61628
rect 31836 61570 31892 61582
rect 31836 61518 31838 61570
rect 31890 61518 31892 61570
rect 31724 61458 31780 61470
rect 31724 61406 31726 61458
rect 31778 61406 31780 61458
rect 31724 59444 31780 61406
rect 31836 60228 31892 61518
rect 32060 61572 32116 61582
rect 31948 61346 32004 61358
rect 31948 61294 31950 61346
rect 32002 61294 32004 61346
rect 31948 61236 32004 61294
rect 31948 61170 32004 61180
rect 32060 60452 32116 61516
rect 32172 61012 32228 63086
rect 32284 62466 32340 62478
rect 32284 62414 32286 62466
rect 32338 62414 32340 62466
rect 32284 61796 32340 62414
rect 32284 61730 32340 61740
rect 32284 61572 32340 61582
rect 32284 61478 32340 61516
rect 32284 61012 32340 61022
rect 32172 60956 32284 61012
rect 32284 60918 32340 60956
rect 32396 61010 32452 64988
rect 32508 64932 32564 65438
rect 33068 65380 33124 67676
rect 33180 67666 33236 67676
rect 33404 67284 33460 67294
rect 33404 67170 33460 67228
rect 33404 67118 33406 67170
rect 33458 67118 33460 67170
rect 33404 67106 33460 67118
rect 33628 67058 33684 67070
rect 33628 67006 33630 67058
rect 33682 67006 33684 67058
rect 33628 66388 33684 67006
rect 33292 66276 33348 66286
rect 33292 66182 33348 66220
rect 33516 66164 33572 66174
rect 33516 66070 33572 66108
rect 33292 65716 33348 65726
rect 33292 65622 33348 65660
rect 33628 65604 33684 66332
rect 33740 65604 33796 67900
rect 33852 68404 33908 68414
rect 34188 68404 34244 71710
rect 34636 71204 34692 72270
rect 34636 71138 34692 71148
rect 34748 71876 34804 71886
rect 34860 71876 34916 71886
rect 34804 71874 34916 71876
rect 34804 71822 34862 71874
rect 34914 71822 34916 71874
rect 34804 71820 34916 71822
rect 34748 70644 34804 71820
rect 34860 71810 34916 71820
rect 34972 71762 35028 71774
rect 34972 71710 34974 71762
rect 35026 71710 35028 71762
rect 34300 70306 34356 70318
rect 34300 70254 34302 70306
rect 34354 70254 34356 70306
rect 34300 68740 34356 70254
rect 34412 70196 34468 70206
rect 34412 70102 34468 70140
rect 34748 69412 34804 70588
rect 34860 71538 34916 71550
rect 34860 71486 34862 71538
rect 34914 71486 34916 71538
rect 34860 70194 34916 71486
rect 34860 70142 34862 70194
rect 34914 70142 34916 70194
rect 34860 70130 34916 70142
rect 34860 69412 34916 69422
rect 34748 69410 34916 69412
rect 34748 69358 34862 69410
rect 34914 69358 34916 69410
rect 34748 69356 34916 69358
rect 34860 69346 34916 69356
rect 34524 69300 34580 69310
rect 34524 69298 34804 69300
rect 34524 69246 34526 69298
rect 34578 69246 34804 69298
rect 34524 69244 34804 69246
rect 34524 69234 34580 69244
rect 34300 68674 34356 68684
rect 33908 68348 34244 68404
rect 33852 67730 33908 68348
rect 33852 67678 33854 67730
rect 33906 67678 33908 67730
rect 33852 67666 33908 67678
rect 34188 68180 34244 68190
rect 34188 67170 34244 68124
rect 34412 68068 34468 68078
rect 34412 67974 34468 68012
rect 34748 68066 34804 69244
rect 34972 68964 35028 71710
rect 35084 69636 35140 72380
rect 35644 72324 35700 72334
rect 35644 72230 35700 72268
rect 35532 71540 35588 71550
rect 35532 71446 35588 71484
rect 35196 71372 35460 71382
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35196 71306 35460 71316
rect 35308 71092 35364 71102
rect 35308 70978 35364 71036
rect 35308 70926 35310 70978
rect 35362 70926 35364 70978
rect 35308 70914 35364 70926
rect 35420 70868 35476 70878
rect 35420 70774 35476 70812
rect 35756 70588 35812 73836
rect 35644 70532 35812 70588
rect 35196 69804 35460 69814
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35196 69738 35460 69748
rect 35084 69580 35252 69636
rect 34972 68898 35028 68908
rect 35084 69412 35140 69422
rect 34748 68014 34750 68066
rect 34802 68014 34804 68066
rect 34748 68002 34804 68014
rect 34972 68514 35028 68526
rect 34972 68462 34974 68514
rect 35026 68462 35028 68514
rect 34188 67118 34190 67170
rect 34242 67118 34244 67170
rect 34188 67106 34244 67118
rect 34300 67058 34356 67070
rect 34300 67006 34302 67058
rect 34354 67006 34356 67058
rect 33852 65604 33908 65614
rect 33740 65602 34132 65604
rect 33740 65550 33854 65602
rect 33906 65550 34132 65602
rect 33740 65548 34132 65550
rect 33628 65538 33684 65548
rect 33852 65538 33908 65548
rect 33404 65492 33460 65502
rect 33404 65398 33460 65436
rect 33516 65380 33572 65390
rect 33068 65324 33348 65380
rect 32508 64866 32564 64876
rect 32620 64708 32676 64718
rect 32620 64614 32676 64652
rect 33068 64594 33124 64606
rect 33068 64542 33070 64594
rect 33122 64542 33124 64594
rect 32732 64372 32788 64382
rect 32508 64148 32564 64158
rect 32508 64034 32564 64092
rect 32508 63982 32510 64034
rect 32562 63982 32564 64034
rect 32508 63970 32564 63982
rect 32732 64036 32788 64316
rect 32620 63924 32676 63934
rect 32620 62466 32676 63868
rect 32620 62414 32622 62466
rect 32674 62414 32676 62466
rect 32620 62402 32676 62414
rect 32508 62354 32564 62366
rect 32508 62302 32510 62354
rect 32562 62302 32564 62354
rect 32508 62244 32564 62302
rect 32732 62244 32788 63980
rect 33068 62468 33124 64542
rect 32508 62188 32788 62244
rect 32956 62412 33124 62468
rect 32956 62020 33012 62412
rect 32956 61954 33012 61964
rect 33180 61796 33236 61806
rect 32396 60958 32398 61010
rect 32450 60958 32452 61010
rect 32396 60946 32452 60958
rect 33068 61740 33180 61796
rect 33068 61012 33124 61740
rect 33180 61730 33236 61740
rect 33292 61684 33348 65324
rect 33516 65286 33572 65324
rect 33852 65268 33908 65278
rect 33404 64932 33460 64942
rect 33460 64876 33572 64932
rect 33404 64866 33460 64876
rect 33292 61618 33348 61628
rect 33404 64706 33460 64718
rect 33404 64654 33406 64706
rect 33458 64654 33460 64706
rect 33404 63362 33460 64654
rect 33516 64036 33572 64876
rect 33516 63942 33572 63980
rect 33628 64818 33684 64830
rect 33628 64766 33630 64818
rect 33682 64766 33684 64818
rect 33404 63310 33406 63362
rect 33458 63310 33460 63362
rect 33180 61572 33236 61582
rect 33180 61478 33236 61516
rect 33292 61458 33348 61470
rect 33292 61406 33294 61458
rect 33346 61406 33348 61458
rect 33292 61012 33348 61406
rect 33404 61460 33460 63310
rect 33404 61394 33460 61404
rect 33516 63138 33572 63150
rect 33516 63086 33518 63138
rect 33570 63086 33572 63138
rect 33068 60956 33236 61012
rect 32508 60900 32564 60910
rect 32844 60900 32900 60910
rect 32508 60898 32844 60900
rect 32508 60846 32510 60898
rect 32562 60846 32844 60898
rect 32508 60844 32844 60846
rect 32508 60834 32564 60844
rect 32844 60834 32900 60844
rect 33068 60786 33124 60798
rect 33068 60734 33070 60786
rect 33122 60734 33124 60786
rect 33068 60452 33124 60734
rect 32060 60396 32452 60452
rect 31836 60162 31892 60172
rect 32172 60228 32228 60238
rect 32060 60116 32116 60126
rect 32060 60022 32116 60060
rect 31724 59378 31780 59388
rect 31836 60004 31892 60014
rect 31836 59890 31892 59948
rect 31836 59838 31838 59890
rect 31890 59838 31892 59890
rect 31612 59278 31614 59330
rect 31666 59278 31668 59330
rect 31612 59266 31668 59278
rect 31724 59220 31780 59230
rect 31836 59220 31892 59838
rect 31724 59218 31892 59220
rect 31724 59166 31726 59218
rect 31778 59166 31892 59218
rect 31724 59164 31892 59166
rect 31724 58434 31780 59164
rect 31948 58436 32004 58446
rect 31724 58382 31726 58434
rect 31778 58382 31780 58434
rect 31724 58370 31780 58382
rect 31836 58434 32004 58436
rect 31836 58382 31950 58434
rect 32002 58382 32004 58434
rect 31836 58380 32004 58382
rect 31836 58212 31892 58380
rect 31948 58370 32004 58380
rect 31836 57988 31892 58156
rect 31612 57932 31892 57988
rect 31612 57874 31668 57932
rect 31612 57822 31614 57874
rect 31666 57822 31668 57874
rect 31612 57810 31668 57822
rect 32172 57538 32228 60172
rect 32396 59332 32452 60396
rect 32956 60396 33124 60452
rect 32956 60116 33012 60396
rect 33068 60228 33124 60238
rect 33068 60134 33124 60172
rect 32844 59890 32900 59902
rect 32844 59838 32846 59890
rect 32898 59838 32900 59890
rect 32844 59444 32900 59838
rect 32844 59378 32900 59388
rect 32284 57876 32340 57886
rect 32396 57876 32452 59276
rect 32508 58994 32564 59006
rect 32508 58942 32510 58994
rect 32562 58942 32564 58994
rect 32508 58772 32564 58942
rect 32508 58706 32564 58716
rect 32956 58660 33012 60060
rect 32956 58594 33012 58604
rect 32732 58548 32788 58558
rect 32284 57874 32452 57876
rect 32284 57822 32286 57874
rect 32338 57822 32452 57874
rect 32284 57820 32452 57822
rect 32508 58492 32732 58548
rect 32284 57810 32340 57820
rect 32508 57762 32564 58492
rect 32732 58454 32788 58492
rect 33180 58434 33236 60956
rect 33292 60676 33348 60956
rect 33516 60900 33572 63086
rect 33628 62354 33684 64766
rect 33852 63924 33908 65212
rect 34076 64932 34132 65548
rect 34188 65492 34244 65502
rect 34188 65398 34244 65436
rect 34076 64876 34244 64932
rect 33852 63830 33908 63868
rect 34076 64706 34132 64718
rect 34076 64654 34078 64706
rect 34130 64654 34132 64706
rect 33628 62302 33630 62354
rect 33682 62302 33684 62354
rect 33628 62290 33684 62302
rect 33852 63138 33908 63150
rect 33852 63086 33854 63138
rect 33906 63086 33908 63138
rect 33292 60620 33460 60676
rect 33404 60452 33460 60620
rect 33516 60674 33572 60844
rect 33628 61684 33684 61694
rect 33628 61570 33684 61628
rect 33628 61518 33630 61570
rect 33682 61518 33684 61570
rect 33628 60788 33684 61518
rect 33628 60722 33684 60732
rect 33740 61572 33796 61582
rect 33740 60898 33796 61516
rect 33740 60846 33742 60898
rect 33794 60846 33796 60898
rect 33516 60622 33518 60674
rect 33570 60622 33572 60674
rect 33516 60610 33572 60622
rect 33740 60564 33796 60846
rect 33628 60508 33796 60564
rect 33852 61236 33908 63086
rect 34076 62188 34132 64654
rect 34188 64372 34244 64876
rect 34300 64596 34356 67006
rect 34972 66612 35028 68462
rect 35084 67282 35140 69356
rect 35196 68402 35252 69580
rect 35644 69522 35700 70532
rect 35756 69972 35812 69982
rect 35868 69972 35924 74060
rect 36092 74022 36148 74060
rect 36316 74050 36372 74060
rect 36092 72324 36148 72334
rect 36092 72230 36148 72268
rect 36764 72324 36820 72334
rect 35980 71932 36708 71988
rect 35980 71874 36036 71932
rect 35980 71822 35982 71874
rect 36034 71822 36036 71874
rect 35980 71810 36036 71822
rect 36092 71764 36148 71774
rect 36092 71762 36260 71764
rect 36092 71710 36094 71762
rect 36146 71710 36260 71762
rect 36092 71708 36260 71710
rect 36092 71698 36148 71708
rect 35756 69970 35924 69972
rect 35756 69918 35758 69970
rect 35810 69918 35924 69970
rect 35756 69916 35924 69918
rect 36092 70754 36148 70766
rect 36092 70702 36094 70754
rect 36146 70702 36148 70754
rect 36092 70196 36148 70702
rect 35756 69906 35812 69916
rect 35644 69470 35646 69522
rect 35698 69470 35700 69522
rect 35644 69458 35700 69470
rect 35868 69412 35924 69422
rect 35868 69318 35924 69356
rect 35196 68350 35198 68402
rect 35250 68350 35252 68402
rect 35196 68338 35252 68350
rect 35532 68852 35588 68862
rect 35196 68236 35460 68246
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35196 68170 35460 68180
rect 35532 67842 35588 68796
rect 36092 68628 36148 70140
rect 35532 67790 35534 67842
rect 35586 67790 35588 67842
rect 35532 67778 35588 67790
rect 35980 68626 36148 68628
rect 35980 68574 36094 68626
rect 36146 68574 36148 68626
rect 35980 68572 36148 68574
rect 35084 67230 35086 67282
rect 35138 67230 35140 67282
rect 35084 67218 35140 67230
rect 35308 67730 35364 67742
rect 35308 67678 35310 67730
rect 35362 67678 35364 67730
rect 35308 67284 35364 67678
rect 35308 67218 35364 67228
rect 35980 67058 36036 68572
rect 36092 68562 36148 68572
rect 36092 67844 36148 67882
rect 36092 67778 36148 67788
rect 36092 67620 36148 67630
rect 36092 67526 36148 67564
rect 35980 67006 35982 67058
rect 36034 67006 36036 67058
rect 35980 66994 36036 67006
rect 35196 66668 35460 66678
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 34972 66556 35140 66612
rect 35196 66602 35460 66612
rect 34636 66388 34692 66398
rect 34636 66294 34692 66332
rect 34860 66276 34916 66286
rect 34748 66274 34916 66276
rect 34748 66222 34862 66274
rect 34914 66222 34916 66274
rect 34748 66220 34916 66222
rect 34748 66164 34804 66220
rect 34860 66210 34916 66220
rect 34748 65716 34804 66108
rect 34524 65660 34804 65716
rect 34972 66164 35028 66174
rect 34524 65378 34580 65660
rect 34524 65326 34526 65378
rect 34578 65326 34580 65378
rect 34300 64530 34356 64540
rect 34412 64594 34468 64606
rect 34412 64542 34414 64594
rect 34466 64542 34468 64594
rect 34412 64372 34468 64542
rect 34188 64316 34468 64372
rect 34412 64036 34468 64046
rect 34524 64036 34580 65326
rect 34636 65492 34692 65502
rect 34636 64706 34692 65436
rect 34972 64930 35028 66108
rect 34972 64878 34974 64930
rect 35026 64878 35028 64930
rect 34972 64866 35028 64878
rect 34636 64654 34638 64706
rect 34690 64654 34692 64706
rect 34636 64642 34692 64654
rect 34860 64596 34916 64606
rect 35084 64596 35140 66556
rect 35420 66276 35476 66286
rect 35420 66164 35476 66220
rect 36204 66276 36260 71708
rect 36316 71762 36372 71774
rect 36316 71710 36318 71762
rect 36370 71710 36372 71762
rect 36316 71652 36372 71710
rect 36316 71092 36372 71596
rect 36316 71026 36372 71036
rect 36652 69636 36708 71932
rect 36764 71986 36820 72268
rect 36764 71934 36766 71986
rect 36818 71934 36820 71986
rect 36764 71922 36820 71934
rect 37212 71652 37268 71662
rect 37212 71558 37268 71596
rect 37660 71652 37716 71662
rect 37660 71558 37716 71596
rect 37212 71090 37268 71102
rect 37212 71038 37214 71090
rect 37266 71038 37268 71090
rect 37212 70980 37268 71038
rect 37212 70914 37268 70924
rect 38220 70868 38276 70878
rect 38220 70866 38388 70868
rect 38220 70814 38222 70866
rect 38274 70814 38388 70866
rect 38220 70812 38388 70814
rect 38220 70802 38276 70812
rect 38220 70644 38276 70654
rect 36988 70196 37044 70206
rect 36876 70194 37044 70196
rect 36876 70142 36990 70194
rect 37042 70142 37044 70194
rect 36876 70140 37044 70142
rect 36876 69972 36932 70140
rect 36988 70130 37044 70140
rect 37324 70196 37380 70206
rect 37324 70082 37380 70140
rect 37324 70030 37326 70082
rect 37378 70030 37380 70082
rect 37324 70018 37380 70030
rect 36876 69906 36932 69916
rect 36652 69580 36932 69636
rect 36764 68626 36820 68638
rect 36764 68574 36766 68626
rect 36818 68574 36820 68626
rect 36764 67620 36820 68574
rect 36876 68066 36932 69580
rect 38220 69522 38276 70588
rect 38220 69470 38222 69522
rect 38274 69470 38276 69522
rect 38220 69458 38276 69470
rect 36876 68014 36878 68066
rect 36930 68014 36932 68066
rect 36876 68002 36932 68014
rect 36988 69410 37044 69422
rect 36988 69358 36990 69410
rect 37042 69358 37044 69410
rect 36764 67554 36820 67564
rect 36988 67284 37044 69358
rect 37212 69298 37268 69310
rect 37212 69246 37214 69298
rect 37266 69246 37268 69298
rect 37212 67844 37268 69246
rect 37324 69298 37380 69310
rect 37324 69246 37326 69298
rect 37378 69246 37380 69298
rect 37324 68964 37380 69246
rect 37772 69188 37828 69198
rect 37324 68898 37380 68908
rect 37548 69186 37828 69188
rect 37548 69134 37774 69186
rect 37826 69134 37828 69186
rect 37548 69132 37828 69134
rect 37548 68514 37604 69132
rect 37772 69122 37828 69132
rect 37548 68462 37550 68514
rect 37602 68462 37604 68514
rect 37548 68450 37604 68462
rect 37884 68964 37940 68974
rect 37324 67956 37380 67966
rect 37324 67862 37380 67900
rect 37548 67844 37604 67854
rect 37212 67778 37268 67788
rect 37436 67842 37604 67844
rect 37436 67790 37550 67842
rect 37602 67790 37604 67842
rect 37436 67788 37604 67790
rect 37436 67508 37492 67788
rect 37548 67778 37604 67788
rect 37772 67842 37828 67854
rect 37772 67790 37774 67842
rect 37826 67790 37828 67842
rect 36988 67218 37044 67228
rect 37324 67452 37492 67508
rect 37324 66500 37380 67452
rect 37436 67284 37492 67294
rect 37772 67284 37828 67790
rect 37492 67228 37828 67284
rect 37436 67170 37492 67228
rect 37436 67118 37438 67170
rect 37490 67118 37492 67170
rect 37436 67106 37492 67118
rect 37884 67060 37940 68908
rect 37772 67058 37940 67060
rect 37772 67006 37886 67058
rect 37938 67006 37940 67058
rect 37772 67004 37940 67006
rect 37324 66444 37492 66500
rect 36204 66210 36260 66220
rect 37324 66274 37380 66286
rect 37324 66222 37326 66274
rect 37378 66222 37380 66274
rect 35420 66162 35588 66164
rect 35420 66110 35422 66162
rect 35474 66110 35588 66162
rect 35420 66108 35588 66110
rect 35420 66098 35476 66108
rect 35196 65490 35252 65502
rect 35196 65438 35198 65490
rect 35250 65438 35252 65490
rect 35196 65268 35252 65438
rect 35196 65202 35252 65212
rect 35196 65100 35460 65110
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35196 65034 35460 65044
rect 35532 64930 35588 66108
rect 36316 66052 36372 66062
rect 35868 66050 36372 66052
rect 35868 65998 36318 66050
rect 36370 65998 36372 66050
rect 35868 65996 36372 65998
rect 35868 65492 35924 65996
rect 36316 65986 36372 65996
rect 36988 66050 37044 66062
rect 36988 65998 36990 66050
rect 37042 65998 37044 66050
rect 35868 65398 35924 65436
rect 35980 65378 36036 65390
rect 35980 65326 35982 65378
rect 36034 65326 36036 65378
rect 35532 64878 35534 64930
rect 35586 64878 35588 64930
rect 35532 64866 35588 64878
rect 35644 65044 35700 65054
rect 34860 64502 34916 64540
rect 34972 64540 35140 64596
rect 34636 64036 34692 64046
rect 34524 64034 34692 64036
rect 34524 63982 34638 64034
rect 34690 63982 34692 64034
rect 34524 63980 34692 63982
rect 34076 62132 34356 62188
rect 33852 60676 33908 61180
rect 33628 60452 33684 60508
rect 33292 60396 33460 60452
rect 33516 60396 33684 60452
rect 33292 59556 33348 60396
rect 33404 59780 33460 59790
rect 33404 59686 33460 59724
rect 33292 59500 33460 59556
rect 33292 59332 33348 59342
rect 33292 59218 33348 59276
rect 33292 59166 33294 59218
rect 33346 59166 33348 59218
rect 33292 59154 33348 59166
rect 33180 58382 33182 58434
rect 33234 58382 33236 58434
rect 33180 58370 33236 58382
rect 33404 58322 33460 59500
rect 33516 59106 33572 60396
rect 33852 59332 33908 60620
rect 33516 59054 33518 59106
rect 33570 59054 33572 59106
rect 33516 58548 33572 59054
rect 33516 58482 33572 58492
rect 33740 59276 33908 59332
rect 34188 60788 34244 60798
rect 33404 58270 33406 58322
rect 33458 58270 33460 58322
rect 33404 58258 33460 58270
rect 33516 58324 33572 58334
rect 33740 58324 33796 59276
rect 34188 58994 34244 60732
rect 34188 58942 34190 58994
rect 34242 58942 34244 58994
rect 33852 58772 33908 58782
rect 33852 58434 33908 58716
rect 33852 58382 33854 58434
rect 33906 58382 33908 58434
rect 33852 58370 33908 58382
rect 33964 58548 34020 58558
rect 33516 58322 33796 58324
rect 33516 58270 33518 58322
rect 33570 58270 33796 58322
rect 33516 58268 33796 58270
rect 33516 58258 33572 58268
rect 32508 57710 32510 57762
rect 32562 57710 32564 57762
rect 32508 57698 32564 57710
rect 33852 57652 33908 57662
rect 33964 57652 34020 58492
rect 32172 57486 32174 57538
rect 32226 57486 32228 57538
rect 32172 57474 32228 57486
rect 33516 57650 34020 57652
rect 33516 57598 33854 57650
rect 33906 57598 34020 57650
rect 33516 57596 34020 57598
rect 34188 57650 34244 58942
rect 34300 57762 34356 62132
rect 34412 62130 34468 63980
rect 34636 63970 34692 63980
rect 34972 63140 35028 64540
rect 34412 62078 34414 62130
rect 34466 62078 34468 62130
rect 34412 62066 34468 62078
rect 34748 62354 34804 62366
rect 34748 62302 34750 62354
rect 34802 62302 34804 62354
rect 34412 61570 34468 61582
rect 34412 61518 34414 61570
rect 34466 61518 34468 61570
rect 34412 59780 34468 61518
rect 34748 61012 34804 62302
rect 34748 60946 34804 60956
rect 34860 62020 34916 62030
rect 34860 60898 34916 61964
rect 34972 61796 35028 63084
rect 35084 63922 35140 63934
rect 35084 63870 35086 63922
rect 35138 63870 35140 63922
rect 35084 62354 35140 63870
rect 35196 63532 35460 63542
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35196 63466 35460 63476
rect 35196 63364 35252 63374
rect 35196 63026 35252 63308
rect 35532 63140 35588 63150
rect 35644 63140 35700 64988
rect 35868 64708 35924 64718
rect 35868 63924 35924 64652
rect 35868 63858 35924 63868
rect 35980 63250 36036 65326
rect 36764 65380 36820 65390
rect 36316 64820 36372 64830
rect 36092 64708 36148 64718
rect 36092 64706 36260 64708
rect 36092 64654 36094 64706
rect 36146 64654 36260 64706
rect 36092 64652 36260 64654
rect 36092 64642 36148 64652
rect 36204 64484 36260 64652
rect 35980 63198 35982 63250
rect 36034 63198 36036 63250
rect 35980 63186 36036 63198
rect 36092 64148 36148 64158
rect 36092 64034 36148 64092
rect 36092 63982 36094 64034
rect 36146 63982 36148 64034
rect 35532 63138 35700 63140
rect 35532 63086 35534 63138
rect 35586 63086 35700 63138
rect 35532 63084 35700 63086
rect 36092 63140 36148 63982
rect 36204 63588 36260 64428
rect 36316 63922 36372 64764
rect 36316 63870 36318 63922
rect 36370 63870 36372 63922
rect 36316 63858 36372 63870
rect 36204 63532 36484 63588
rect 36092 63138 36372 63140
rect 36092 63086 36094 63138
rect 36146 63086 36372 63138
rect 36092 63084 36372 63086
rect 35532 63074 35588 63084
rect 36092 63074 36148 63084
rect 35196 62974 35198 63026
rect 35250 62974 35252 63026
rect 35196 62962 35252 62974
rect 35084 62302 35086 62354
rect 35138 62302 35140 62354
rect 35084 62132 35140 62302
rect 36316 62188 36372 63084
rect 36428 63028 36484 63532
rect 36428 62934 36484 62972
rect 36652 63364 36708 63374
rect 35084 62066 35140 62076
rect 36092 62132 36372 62188
rect 36428 62354 36484 62366
rect 36428 62302 36430 62354
rect 36482 62302 36484 62354
rect 36428 62188 36484 62302
rect 36652 62354 36708 63308
rect 36652 62302 36654 62354
rect 36706 62302 36708 62354
rect 36652 62290 36708 62302
rect 36764 62188 36820 65324
rect 36988 65044 37044 65998
rect 37324 65380 37380 66222
rect 37324 65314 37380 65324
rect 37436 65490 37492 66444
rect 37436 65438 37438 65490
rect 37490 65438 37492 65490
rect 36988 64978 37044 64988
rect 36988 64820 37044 64830
rect 36988 64726 37044 64764
rect 37100 64706 37156 64718
rect 37100 64654 37102 64706
rect 37154 64654 37156 64706
rect 37100 64260 37156 64654
rect 36428 62132 36820 62188
rect 36876 64204 37100 64260
rect 35196 61964 35460 61974
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35196 61898 35460 61908
rect 34972 61740 35588 61796
rect 35532 61684 35588 61740
rect 35756 61684 35812 61694
rect 35532 61682 35812 61684
rect 35532 61630 35758 61682
rect 35810 61630 35812 61682
rect 35532 61628 35812 61630
rect 35420 61570 35476 61582
rect 35420 61518 35422 61570
rect 35474 61518 35476 61570
rect 34860 60846 34862 60898
rect 34914 60846 34916 60898
rect 34860 60564 34916 60846
rect 35308 61460 35364 61470
rect 35308 60786 35364 61404
rect 35308 60734 35310 60786
rect 35362 60734 35364 60786
rect 35308 60722 35364 60734
rect 35420 60564 35476 61518
rect 34860 60228 34916 60508
rect 34636 60172 34916 60228
rect 35084 60508 35476 60564
rect 34636 60114 34692 60172
rect 34636 60062 34638 60114
rect 34690 60062 34692 60114
rect 34636 60050 34692 60062
rect 34412 59714 34468 59724
rect 34860 60004 34916 60014
rect 35084 60004 35140 60508
rect 35196 60396 35460 60406
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35196 60330 35460 60340
rect 34860 60002 35140 60004
rect 34860 59950 34862 60002
rect 34914 59950 35140 60002
rect 34860 59948 35140 59950
rect 34860 59444 34916 59948
rect 34860 58546 34916 59388
rect 35308 59332 35364 59342
rect 35308 59220 35364 59276
rect 35532 59220 35588 59230
rect 35308 59218 35532 59220
rect 35308 59166 35310 59218
rect 35362 59166 35532 59218
rect 35308 59164 35532 59166
rect 35308 59154 35364 59164
rect 34860 58494 34862 58546
rect 34914 58494 34916 58546
rect 34860 58482 34916 58494
rect 34972 58996 35028 59006
rect 34300 57710 34302 57762
rect 34354 57710 34356 57762
rect 34300 57698 34356 57710
rect 34188 57598 34190 57650
rect 34242 57598 34244 57650
rect 31948 56980 32004 56990
rect 31948 56886 32004 56924
rect 33516 56978 33572 57596
rect 33852 57586 33908 57596
rect 34188 57540 34244 57598
rect 34300 57540 34356 57550
rect 34188 57484 34300 57540
rect 34300 57474 34356 57484
rect 33516 56926 33518 56978
rect 33570 56926 33572 56978
rect 33516 56914 33572 56926
rect 33852 56980 33908 56990
rect 34972 56980 35028 58940
rect 35196 58828 35460 58838
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35196 58762 35460 58772
rect 35532 58434 35588 59164
rect 35532 58382 35534 58434
rect 35586 58382 35588 58434
rect 35532 58370 35588 58382
rect 35532 57650 35588 57662
rect 35532 57598 35534 57650
rect 35586 57598 35588 57650
rect 33852 56978 35028 56980
rect 33852 56926 33854 56978
rect 33906 56926 35028 56978
rect 33852 56924 35028 56926
rect 35084 57540 35140 57550
rect 35084 56980 35140 57484
rect 35196 57260 35460 57270
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35196 57194 35460 57204
rect 35196 56980 35252 56990
rect 35084 56978 35252 56980
rect 35084 56926 35198 56978
rect 35250 56926 35252 56978
rect 35084 56924 35252 56926
rect 35532 56980 35588 57598
rect 35756 57538 35812 61628
rect 35980 60676 36036 60686
rect 36092 60676 36148 62132
rect 35980 60674 36148 60676
rect 35980 60622 35982 60674
rect 36034 60622 36148 60674
rect 35980 60620 36148 60622
rect 36204 61458 36260 61470
rect 36204 61406 36206 61458
rect 36258 61406 36260 61458
rect 35980 60610 36036 60620
rect 35868 59890 35924 59902
rect 35868 59838 35870 59890
rect 35922 59838 35924 59890
rect 35868 59780 35924 59838
rect 35868 59714 35924 59724
rect 36204 59556 36260 61406
rect 36428 60786 36484 62132
rect 36428 60734 36430 60786
rect 36482 60734 36484 60786
rect 36316 59780 36372 59790
rect 36428 59780 36484 60734
rect 36316 59778 36484 59780
rect 36316 59726 36318 59778
rect 36370 59726 36484 59778
rect 36316 59724 36484 59726
rect 36316 59714 36372 59724
rect 36204 59500 36372 59556
rect 36316 59332 36372 59500
rect 36316 59238 36372 59276
rect 36204 59218 36260 59230
rect 36204 59166 36206 59218
rect 36258 59166 36260 59218
rect 36204 58996 36260 59166
rect 36428 59220 36484 59230
rect 36428 59126 36484 59164
rect 35868 58660 35924 58670
rect 35868 57650 35924 58604
rect 36204 58322 36260 58940
rect 36204 58270 36206 58322
rect 36258 58270 36260 58322
rect 36204 58258 36260 58270
rect 36540 57764 36596 57774
rect 36876 57764 36932 64204
rect 37100 64194 37156 64204
rect 37324 64594 37380 64606
rect 37324 64542 37326 64594
rect 37378 64542 37380 64594
rect 37324 64372 37380 64542
rect 37324 62188 37380 64316
rect 37436 64596 37492 65438
rect 37436 64034 37492 64540
rect 37436 63982 37438 64034
rect 37490 63982 37492 64034
rect 37436 63970 37492 63982
rect 37548 66162 37604 66174
rect 37548 66110 37550 66162
rect 37602 66110 37604 66162
rect 37548 65716 37604 66110
rect 37548 63364 37604 65660
rect 37772 65378 37828 67004
rect 37884 66994 37940 67004
rect 37772 65326 37774 65378
rect 37826 65326 37828 65378
rect 37772 65314 37828 65326
rect 37884 65268 37940 65278
rect 37884 64706 37940 65212
rect 37884 64654 37886 64706
rect 37938 64654 37940 64706
rect 37884 64642 37940 64654
rect 38220 64594 38276 64606
rect 38220 64542 38222 64594
rect 38274 64542 38276 64594
rect 38108 64482 38164 64494
rect 38108 64430 38110 64482
rect 38162 64430 38164 64482
rect 37548 63270 37604 63308
rect 37996 63924 38052 63934
rect 38108 63924 38164 64430
rect 38220 64148 38276 64542
rect 38220 64082 38276 64092
rect 38220 63924 38276 63934
rect 38108 63922 38276 63924
rect 38108 63870 38222 63922
rect 38274 63870 38276 63922
rect 38108 63868 38276 63870
rect 37548 63140 37604 63150
rect 37548 63046 37604 63084
rect 37884 63138 37940 63150
rect 37884 63086 37886 63138
rect 37938 63086 37940 63138
rect 37324 62132 37492 62188
rect 36988 61796 37044 61806
rect 36988 61570 37044 61740
rect 36988 61518 36990 61570
rect 37042 61518 37044 61570
rect 36988 61506 37044 61518
rect 37212 61458 37268 61470
rect 37212 61406 37214 61458
rect 37266 61406 37268 61458
rect 37212 61348 37268 61406
rect 37100 60564 37156 60574
rect 36988 59780 37044 59790
rect 36988 58434 37044 59724
rect 36988 58382 36990 58434
rect 37042 58382 37044 58434
rect 36988 58370 37044 58382
rect 37100 59218 37156 60508
rect 37212 59668 37268 61292
rect 37212 59602 37268 59612
rect 37436 61458 37492 62132
rect 37436 61406 37438 61458
rect 37490 61406 37492 61458
rect 37100 59166 37102 59218
rect 37154 59166 37156 59218
rect 36540 57762 36932 57764
rect 36540 57710 36542 57762
rect 36594 57710 36932 57762
rect 36540 57708 36932 57710
rect 37100 58322 37156 59166
rect 37100 58270 37102 58322
rect 37154 58270 37156 58322
rect 36540 57698 36596 57708
rect 35868 57598 35870 57650
rect 35922 57598 35924 57650
rect 35868 57586 35924 57598
rect 35756 57486 35758 57538
rect 35810 57486 35812 57538
rect 35756 57474 35812 57486
rect 37100 57538 37156 58270
rect 37212 58660 37268 58670
rect 37212 57650 37268 58604
rect 37436 58546 37492 61406
rect 37660 62132 37716 62142
rect 37548 61012 37604 61022
rect 37548 60226 37604 60956
rect 37660 60786 37716 62076
rect 37884 62020 37940 63086
rect 37996 62578 38052 63868
rect 37996 62526 37998 62578
rect 38050 62526 38052 62578
rect 37996 62514 38052 62526
rect 38220 63028 38276 63868
rect 38108 62242 38164 62254
rect 38108 62190 38110 62242
rect 38162 62190 38164 62242
rect 38108 62132 38164 62190
rect 38108 62066 38164 62076
rect 37884 61954 37940 61964
rect 37884 61796 37940 61806
rect 37772 61684 37828 61694
rect 37772 61590 37828 61628
rect 37660 60734 37662 60786
rect 37714 60734 37716 60786
rect 37660 60722 37716 60734
rect 37548 60174 37550 60226
rect 37602 60174 37604 60226
rect 37548 60162 37604 60174
rect 37660 60564 37716 60574
rect 37660 60114 37716 60508
rect 37660 60062 37662 60114
rect 37714 60062 37716 60114
rect 37660 60050 37716 60062
rect 37884 60004 37940 61740
rect 38108 61684 38164 61694
rect 38220 61684 38276 62972
rect 38164 61628 38276 61684
rect 38108 61618 38164 61628
rect 37772 60002 37940 60004
rect 37772 59950 37886 60002
rect 37938 59950 37940 60002
rect 37772 59948 37940 59950
rect 37660 59668 37716 59678
rect 37660 59442 37716 59612
rect 37660 59390 37662 59442
rect 37714 59390 37716 59442
rect 37660 59378 37716 59390
rect 37772 58660 37828 59948
rect 37884 59938 37940 59948
rect 37884 59444 37940 59454
rect 37884 59350 37940 59388
rect 37996 59332 38052 59342
rect 37996 59238 38052 59276
rect 37772 58594 37828 58604
rect 38332 58548 38388 70812
rect 37436 58494 37438 58546
rect 37490 58494 37492 58546
rect 37436 58482 37492 58494
rect 37884 58492 38388 58548
rect 37884 57874 37940 58492
rect 37884 57822 37886 57874
rect 37938 57822 37940 57874
rect 37884 57810 37940 57822
rect 38220 58324 38276 58334
rect 38220 57764 38276 58268
rect 38220 57762 38388 57764
rect 38220 57710 38222 57762
rect 38274 57710 38388 57762
rect 38220 57708 38388 57710
rect 38220 57698 38276 57708
rect 37212 57598 37214 57650
rect 37266 57598 37268 57650
rect 37212 57586 37268 57598
rect 37100 57486 37102 57538
rect 37154 57486 37156 57538
rect 37100 57474 37156 57486
rect 35644 56980 35700 56990
rect 35532 56978 35700 56980
rect 35532 56926 35646 56978
rect 35698 56926 35700 56978
rect 35532 56924 35700 56926
rect 33852 56914 33908 56924
rect 34972 56866 35028 56924
rect 35196 56914 35252 56924
rect 35644 56914 35700 56924
rect 38332 56978 38388 57708
rect 38332 56926 38334 56978
rect 38386 56926 38388 56978
rect 38332 56914 38388 56926
rect 34972 56814 34974 56866
rect 35026 56814 35028 56866
rect 34972 56802 35028 56814
rect 31836 56308 31892 56318
rect 31836 53732 31892 56252
rect 35196 55692 35460 55702
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35196 55626 35460 55636
rect 32284 55412 32340 55422
rect 32172 55356 32284 55412
rect 32060 54404 32116 54414
rect 32060 53842 32116 54348
rect 32060 53790 32062 53842
rect 32114 53790 32116 53842
rect 32060 53778 32116 53790
rect 31836 53666 31892 53676
rect 31500 52770 31556 52780
rect 31388 52724 31444 52734
rect 31276 52276 31332 52286
rect 31164 52274 31332 52276
rect 31164 52222 31278 52274
rect 31330 52222 31332 52274
rect 31164 52220 31332 52222
rect 31276 52210 31332 52220
rect 30716 51550 30718 51602
rect 30770 51550 30772 51602
rect 30716 51538 30772 51550
rect 31164 51604 31220 51614
rect 31388 51604 31444 52668
rect 31164 51602 31444 51604
rect 31164 51550 31166 51602
rect 31218 51550 31444 51602
rect 31164 51548 31444 51550
rect 31164 51380 31220 51548
rect 31164 51314 31220 51324
rect 30604 50372 30884 50428
rect 30716 49698 30772 49710
rect 30716 49646 30718 49698
rect 30770 49646 30772 49698
rect 30716 49364 30772 49646
rect 30716 49298 30772 49308
rect 30268 49028 30324 49038
rect 30380 49028 30436 49196
rect 30492 49140 30548 49150
rect 30492 49138 30772 49140
rect 30492 49086 30494 49138
rect 30546 49086 30772 49138
rect 30492 49084 30772 49086
rect 30492 49074 30548 49084
rect 30268 49026 30436 49028
rect 30268 48974 30270 49026
rect 30322 48974 30436 49026
rect 30268 48972 30436 48974
rect 30268 48962 30324 48972
rect 30604 48916 30660 48926
rect 30604 48822 30660 48860
rect 30492 48802 30548 48814
rect 30492 48750 30494 48802
rect 30546 48750 30548 48802
rect 30492 48132 30548 48750
rect 30492 48066 30548 48076
rect 30716 47908 30772 49084
rect 30044 46732 30212 46788
rect 30268 47852 30772 47908
rect 29932 46452 29988 46462
rect 29932 42868 29988 46396
rect 30044 44100 30100 46732
rect 30156 46562 30212 46574
rect 30156 46510 30158 46562
rect 30210 46510 30212 46562
rect 30156 45892 30212 46510
rect 30268 46116 30324 47852
rect 30828 47684 30884 50372
rect 31164 49252 31220 49262
rect 31164 49138 31220 49196
rect 31164 49086 31166 49138
rect 31218 49086 31220 49138
rect 31164 49074 31220 49086
rect 31276 48468 31332 51548
rect 30492 47628 30884 47684
rect 31164 48412 31332 48468
rect 31724 49138 31780 49150
rect 31724 49086 31726 49138
rect 31778 49086 31780 49138
rect 30492 46228 30548 47628
rect 30828 47460 30884 47470
rect 30828 47366 30884 47404
rect 31052 47460 31108 47470
rect 30940 47236 30996 47246
rect 30604 46562 30660 46574
rect 30604 46510 30606 46562
rect 30658 46510 30660 46562
rect 30604 46452 30660 46510
rect 30604 46386 30660 46396
rect 30492 46162 30548 46172
rect 30268 46050 30324 46060
rect 30604 46004 30660 46014
rect 30604 45910 30660 45948
rect 30156 45836 30324 45892
rect 30156 45666 30212 45678
rect 30156 45614 30158 45666
rect 30210 45614 30212 45666
rect 30156 44436 30212 45614
rect 30156 44370 30212 44380
rect 30268 44996 30324 45836
rect 30380 44996 30436 45006
rect 30268 44994 30436 44996
rect 30268 44942 30382 44994
rect 30434 44942 30436 44994
rect 30268 44940 30436 44942
rect 30268 44322 30324 44940
rect 30380 44930 30436 44940
rect 30828 44994 30884 45006
rect 30828 44942 30830 44994
rect 30882 44942 30884 44994
rect 30828 44660 30884 44942
rect 30828 44594 30884 44604
rect 30268 44270 30270 44322
rect 30322 44270 30324 44322
rect 30268 44258 30324 44270
rect 30492 44548 30548 44558
rect 30492 44322 30548 44492
rect 30940 44436 30996 47180
rect 31052 46002 31108 47404
rect 31164 46452 31220 48412
rect 31724 48356 31780 49086
rect 31724 48290 31780 48300
rect 31388 48132 31444 48142
rect 31388 48038 31444 48076
rect 31724 48020 31780 48030
rect 31500 48018 31780 48020
rect 31500 47966 31726 48018
rect 31778 47966 31780 48018
rect 31500 47964 31780 47966
rect 31500 47684 31556 47964
rect 31724 47954 31780 47964
rect 32060 48018 32116 48030
rect 32060 47966 32062 48018
rect 32114 47966 32116 48018
rect 31276 47628 31556 47684
rect 31276 47458 31332 47628
rect 31276 47406 31278 47458
rect 31330 47406 31332 47458
rect 31276 47394 31332 47406
rect 31836 47460 31892 47470
rect 31500 47348 31556 47358
rect 31500 47254 31556 47292
rect 31164 46386 31220 46396
rect 31052 45950 31054 46002
rect 31106 45950 31108 46002
rect 31052 45938 31108 45950
rect 31164 46116 31220 46126
rect 31164 44436 31220 46060
rect 31276 44996 31332 45006
rect 31724 44996 31780 45006
rect 31276 44994 31780 44996
rect 31276 44942 31278 44994
rect 31330 44942 31726 44994
rect 31778 44942 31780 44994
rect 31276 44940 31780 44942
rect 31276 44930 31332 44940
rect 31164 44380 31332 44436
rect 30940 44370 30996 44380
rect 30492 44270 30494 44322
rect 30546 44270 30548 44322
rect 30492 44258 30548 44270
rect 30604 44212 30660 44250
rect 30604 44146 30660 44156
rect 30828 44212 30884 44222
rect 30380 44100 30436 44110
rect 30044 44044 30212 44100
rect 30044 43316 30100 43326
rect 30044 42978 30100 43260
rect 30044 42926 30046 42978
rect 30098 42926 30100 42978
rect 30044 42914 30100 42926
rect 29932 42802 29988 42812
rect 30156 42308 30212 44044
rect 30380 44006 30436 44044
rect 30716 44098 30772 44110
rect 30716 44046 30718 44098
rect 30770 44046 30772 44098
rect 30716 43316 30772 44046
rect 30716 43250 30772 43260
rect 30828 43428 30884 44156
rect 30604 42868 30660 42878
rect 30604 42754 30660 42812
rect 30604 42702 30606 42754
rect 30658 42702 30660 42754
rect 30044 42252 30212 42308
rect 30380 42642 30436 42654
rect 30380 42590 30382 42642
rect 30434 42590 30436 42642
rect 29932 42196 29988 42206
rect 29932 42082 29988 42140
rect 29932 42030 29934 42082
rect 29986 42030 29988 42082
rect 29932 42018 29988 42030
rect 29596 40514 29876 40516
rect 29596 40462 29598 40514
rect 29650 40462 29876 40514
rect 29596 40460 29876 40462
rect 29596 40450 29652 40460
rect 29820 39842 29876 40460
rect 30044 40292 30100 42252
rect 30380 42196 30436 42590
rect 30380 42130 30436 42140
rect 30492 41972 30548 41982
rect 30492 41878 30548 41916
rect 30604 41748 30660 42702
rect 30828 42084 30884 43372
rect 31164 44210 31220 44222
rect 31164 44158 31166 44210
rect 31218 44158 31220 44210
rect 30940 43316 30996 43326
rect 30940 43204 30996 43260
rect 30940 43148 31108 43204
rect 30940 42980 30996 42990
rect 30940 42886 30996 42924
rect 30828 42018 30884 42028
rect 30492 41692 30660 41748
rect 30940 41858 30996 41870
rect 30940 41806 30942 41858
rect 30994 41806 30996 41858
rect 30940 41748 30996 41806
rect 30156 41410 30212 41422
rect 30156 41358 30158 41410
rect 30210 41358 30212 41410
rect 30156 41298 30212 41358
rect 30492 41412 30548 41692
rect 30940 41682 30996 41692
rect 30940 41524 30996 41534
rect 30492 41346 30548 41356
rect 30604 41410 30660 41422
rect 30604 41358 30606 41410
rect 30658 41358 30660 41410
rect 30156 41246 30158 41298
rect 30210 41246 30212 41298
rect 30156 41234 30212 41246
rect 30604 41300 30660 41358
rect 30604 41298 30772 41300
rect 30604 41246 30606 41298
rect 30658 41246 30772 41298
rect 30604 41244 30772 41246
rect 30604 41234 30660 41244
rect 30492 40626 30548 40638
rect 30492 40574 30494 40626
rect 30546 40574 30548 40626
rect 30044 40226 30100 40236
rect 30268 40402 30324 40414
rect 30268 40350 30270 40402
rect 30322 40350 30324 40402
rect 29820 39790 29822 39842
rect 29874 39790 29876 39842
rect 29820 39778 29876 39790
rect 29932 39508 29988 39518
rect 29932 39506 30212 39508
rect 29932 39454 29934 39506
rect 29986 39454 30212 39506
rect 29932 39452 30212 39454
rect 29932 39442 29988 39452
rect 29260 38612 29428 38668
rect 30156 38722 30212 39452
rect 30156 38670 30158 38722
rect 30210 38670 30212 38722
rect 30156 38658 30212 38670
rect 28924 35812 28980 37436
rect 29148 37604 29204 37614
rect 29148 36482 29204 37548
rect 29148 36430 29150 36482
rect 29202 36430 29204 36482
rect 29148 36418 29204 36430
rect 28924 34132 28980 35756
rect 29148 35700 29204 35710
rect 29148 35606 29204 35644
rect 29260 34356 29316 38612
rect 30268 36708 30324 40350
rect 30492 39844 30548 40574
rect 30492 39778 30548 39788
rect 30380 39730 30436 39742
rect 30380 39678 30382 39730
rect 30434 39678 30436 39730
rect 30380 36708 30436 39678
rect 30492 39284 30548 39294
rect 30492 38836 30548 39228
rect 30604 38948 30660 38958
rect 30604 38854 30660 38892
rect 30492 38162 30548 38780
rect 30716 38612 30772 41244
rect 30716 38546 30772 38556
rect 30492 38110 30494 38162
rect 30546 38110 30548 38162
rect 30492 38098 30548 38110
rect 30380 36652 30660 36708
rect 30268 36642 30324 36652
rect 30156 36482 30212 36494
rect 30156 36430 30158 36482
rect 30210 36430 30212 36482
rect 30044 34580 30100 34590
rect 29372 34356 29428 34366
rect 29260 34354 29428 34356
rect 29260 34302 29374 34354
rect 29426 34302 29428 34354
rect 29260 34300 29428 34302
rect 29372 34290 29428 34300
rect 29148 34132 29204 34142
rect 29484 34132 29540 34142
rect 28924 34130 29204 34132
rect 28924 34078 29150 34130
rect 29202 34078 29204 34130
rect 28924 34076 29204 34078
rect 29148 34066 29204 34076
rect 29372 34130 29540 34132
rect 29372 34078 29486 34130
rect 29538 34078 29540 34130
rect 29372 34076 29540 34078
rect 29260 33572 29316 33582
rect 29372 33572 29428 34076
rect 29484 34066 29540 34076
rect 29260 33570 29428 33572
rect 29260 33518 29262 33570
rect 29314 33518 29428 33570
rect 29260 33516 29428 33518
rect 29484 33572 29540 33582
rect 29540 33516 29764 33572
rect 29260 33348 29316 33516
rect 29484 33506 29540 33516
rect 29260 33282 29316 33292
rect 29148 33236 29204 33246
rect 28812 32946 28868 32956
rect 28924 33234 29204 33236
rect 28924 33182 29150 33234
rect 29202 33182 29204 33234
rect 28924 33180 29204 33182
rect 28924 32340 28980 33180
rect 29148 33170 29204 33180
rect 29708 32450 29764 33516
rect 29708 32398 29710 32450
rect 29762 32398 29764 32450
rect 29708 32386 29764 32398
rect 30044 32452 30100 34524
rect 30156 34356 30212 36430
rect 30604 35812 30660 36652
rect 30940 36258 30996 41468
rect 31052 39396 31108 43148
rect 31164 42980 31220 44158
rect 31164 42914 31220 42924
rect 31276 42308 31332 44380
rect 31388 43876 31444 44940
rect 31724 44930 31780 44940
rect 31500 44100 31556 44110
rect 31500 44098 31780 44100
rect 31500 44046 31502 44098
rect 31554 44046 31780 44098
rect 31500 44044 31780 44046
rect 31500 44034 31556 44044
rect 31388 43820 31556 43876
rect 31388 43204 31444 43214
rect 31388 42866 31444 43148
rect 31500 43092 31556 43820
rect 31724 43650 31780 44044
rect 31724 43598 31726 43650
rect 31778 43598 31780 43650
rect 31724 43586 31780 43598
rect 31500 43026 31556 43036
rect 31388 42814 31390 42866
rect 31442 42814 31444 42866
rect 31388 42802 31444 42814
rect 31836 42532 31892 47404
rect 32060 47012 32116 47966
rect 32060 46946 32116 46956
rect 31948 44660 32004 44670
rect 31948 44434 32004 44604
rect 31948 44382 31950 44434
rect 32002 44382 32004 44434
rect 31948 44370 32004 44382
rect 31948 42532 32004 42542
rect 31836 42530 31948 42532
rect 31836 42478 31838 42530
rect 31890 42478 31948 42530
rect 31836 42476 31948 42478
rect 31836 42466 31892 42476
rect 31276 42252 31444 42308
rect 31276 42084 31332 42094
rect 31276 41990 31332 42028
rect 31388 41860 31444 42252
rect 31276 41804 31444 41860
rect 31500 41860 31556 41870
rect 31052 39340 31220 39396
rect 31052 37492 31108 37502
rect 31052 36482 31108 37436
rect 31052 36430 31054 36482
rect 31106 36430 31108 36482
rect 31052 36418 31108 36430
rect 30940 36206 30942 36258
rect 30994 36206 30996 36258
rect 30940 36194 30996 36206
rect 30604 35718 30660 35756
rect 31052 35924 31108 35934
rect 30828 35698 30884 35710
rect 30828 35646 30830 35698
rect 30882 35646 30884 35698
rect 30268 34916 30324 34926
rect 30268 34822 30324 34860
rect 30828 34916 30884 35646
rect 30828 34850 30884 34860
rect 30940 35586 30996 35598
rect 30940 35534 30942 35586
rect 30994 35534 30996 35586
rect 30156 34290 30212 34300
rect 30940 34244 30996 35534
rect 31052 34468 31108 35868
rect 31164 35922 31220 39340
rect 31276 36708 31332 41804
rect 31500 41746 31556 41804
rect 31836 41748 31892 41758
rect 31500 41694 31502 41746
rect 31554 41694 31556 41746
rect 31388 41636 31444 41646
rect 31388 39058 31444 41580
rect 31500 41412 31556 41694
rect 31500 41346 31556 41356
rect 31612 41746 31892 41748
rect 31612 41694 31838 41746
rect 31890 41694 31892 41746
rect 31612 41692 31892 41694
rect 31500 41188 31556 41198
rect 31612 41188 31668 41692
rect 31836 41682 31892 41692
rect 31500 41186 31668 41188
rect 31500 41134 31502 41186
rect 31554 41134 31668 41186
rect 31500 41132 31668 41134
rect 31500 41122 31556 41132
rect 31724 40962 31780 40974
rect 31724 40910 31726 40962
rect 31778 40910 31780 40962
rect 31724 39732 31780 40910
rect 31724 39666 31780 39676
rect 31948 39620 32004 42476
rect 32172 41412 32228 55356
rect 32284 55318 32340 55356
rect 35420 55298 35476 55310
rect 35420 55246 35422 55298
rect 35474 55246 35476 55298
rect 34860 55188 34916 55198
rect 34860 55094 34916 55132
rect 35420 55188 35476 55246
rect 35420 55122 35476 55132
rect 36428 55188 36484 55198
rect 35756 55076 35812 55086
rect 35644 55074 35812 55076
rect 35644 55022 35758 55074
rect 35810 55022 35812 55074
rect 35644 55020 35812 55022
rect 33180 54626 33236 54638
rect 33180 54574 33182 54626
rect 33234 54574 33236 54626
rect 33180 53842 33236 54574
rect 33404 54516 33460 54526
rect 33180 53790 33182 53842
rect 33234 53790 33236 53842
rect 33180 53778 33236 53790
rect 33292 54514 33460 54516
rect 33292 54462 33406 54514
rect 33458 54462 33460 54514
rect 33292 54460 33460 54462
rect 32396 53732 32452 53742
rect 32396 53638 32452 53676
rect 33068 53172 33124 53182
rect 33292 53172 33348 54460
rect 33404 54450 33460 54460
rect 35308 54514 35364 54526
rect 35308 54462 35310 54514
rect 35362 54462 35364 54514
rect 35308 54292 35364 54462
rect 35084 54236 35364 54292
rect 33068 53170 33348 53172
rect 33068 53118 33070 53170
rect 33122 53118 33348 53170
rect 33068 53116 33348 53118
rect 33852 53732 33908 53742
rect 33852 53172 33908 53676
rect 33068 53106 33124 53116
rect 32284 52948 32340 52958
rect 32284 52854 32340 52892
rect 33628 52834 33684 52846
rect 33628 52782 33630 52834
rect 33682 52782 33684 52834
rect 33404 52724 33460 52734
rect 33404 52630 33460 52668
rect 33404 52276 33460 52286
rect 33628 52276 33684 52782
rect 33404 52274 33684 52276
rect 33404 52222 33406 52274
rect 33458 52222 33684 52274
rect 33404 52220 33684 52222
rect 33404 52210 33460 52220
rect 33628 50148 33684 52220
rect 33852 52274 33908 53116
rect 34972 53172 35028 53182
rect 35084 53172 35140 54236
rect 35196 54124 35460 54134
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35196 54058 35460 54068
rect 35028 53116 35140 53172
rect 34972 53078 35028 53116
rect 34076 52834 34132 52846
rect 34076 52782 34078 52834
rect 34130 52782 34132 52834
rect 34076 52724 34132 52782
rect 34076 52658 34132 52668
rect 33852 52222 33854 52274
rect 33906 52222 33908 52274
rect 33852 52210 33908 52222
rect 35084 50708 35140 53116
rect 35308 53842 35364 53854
rect 35308 53790 35310 53842
rect 35362 53790 35364 53842
rect 35308 53060 35364 53790
rect 35308 53004 35588 53060
rect 35308 52836 35364 52846
rect 35308 52742 35364 52780
rect 35196 52556 35460 52566
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35196 52490 35460 52500
rect 35532 52388 35588 53004
rect 35420 52332 35588 52388
rect 35644 52724 35700 55020
rect 35756 55010 35812 55020
rect 36092 54404 36148 54414
rect 36092 54402 36372 54404
rect 36092 54350 36094 54402
rect 36146 54350 36372 54402
rect 36092 54348 36372 54350
rect 36092 54338 36148 54348
rect 35308 52162 35364 52174
rect 35308 52110 35310 52162
rect 35362 52110 35364 52162
rect 35308 51940 35364 52110
rect 35420 51940 35476 52332
rect 35532 52164 35588 52174
rect 35644 52164 35700 52668
rect 35980 53618 36036 53630
rect 35980 53566 35982 53618
rect 36034 53566 36036 53618
rect 35868 52388 35924 52398
rect 35980 52388 36036 53566
rect 36316 53618 36372 54348
rect 36316 53566 36318 53618
rect 36370 53566 36372 53618
rect 36316 53554 36372 53566
rect 35868 52386 36036 52388
rect 35868 52334 35870 52386
rect 35922 52334 36036 52386
rect 35868 52332 36036 52334
rect 35868 52322 35924 52332
rect 35532 52162 35644 52164
rect 35532 52110 35534 52162
rect 35586 52110 35644 52162
rect 35532 52108 35644 52110
rect 35532 52098 35588 52108
rect 35308 51884 35588 51940
rect 35196 50988 35460 50998
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35196 50922 35460 50932
rect 35196 50708 35252 50718
rect 33516 50092 33684 50148
rect 34748 50706 35252 50708
rect 34748 50654 35198 50706
rect 35250 50654 35252 50706
rect 34748 50652 35252 50654
rect 34748 50372 34804 50652
rect 35196 50642 35252 50652
rect 33516 49700 33572 50092
rect 33628 49924 33684 49934
rect 33628 49922 33908 49924
rect 33628 49870 33630 49922
rect 33682 49870 33908 49922
rect 33628 49868 33908 49870
rect 33628 49858 33684 49868
rect 33516 49644 33684 49700
rect 33628 48354 33684 49644
rect 33740 49252 33796 49262
rect 33740 48468 33796 49196
rect 33852 49138 33908 49868
rect 33964 49810 34020 49822
rect 33964 49758 33966 49810
rect 34018 49758 34020 49810
rect 33964 49700 34020 49758
rect 34636 49700 34692 49710
rect 33964 49698 34692 49700
rect 33964 49646 34638 49698
rect 34690 49646 34692 49698
rect 33964 49644 34692 49646
rect 34636 49634 34692 49644
rect 33852 49086 33854 49138
rect 33906 49086 33908 49138
rect 33852 49074 33908 49086
rect 34636 49028 34692 49038
rect 34748 49028 34804 50316
rect 34636 49026 34804 49028
rect 34636 48974 34638 49026
rect 34690 48974 34804 49026
rect 34636 48972 34804 48974
rect 34860 50370 34916 50382
rect 34860 50318 34862 50370
rect 34914 50318 34916 50370
rect 34636 48962 34692 48972
rect 34188 48916 34244 48926
rect 33852 48468 33908 48478
rect 33740 48412 33852 48468
rect 33852 48374 33908 48412
rect 34188 48466 34244 48860
rect 34860 48804 34916 50318
rect 34972 49812 35028 49822
rect 34972 49718 35028 49756
rect 35196 49700 35252 49710
rect 35084 49698 35252 49700
rect 35084 49646 35198 49698
rect 35250 49646 35252 49698
rect 35084 49644 35252 49646
rect 35084 49028 35140 49644
rect 35196 49634 35252 49644
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35196 49354 35460 49364
rect 35308 49028 35364 49038
rect 35084 49026 35364 49028
rect 35084 48974 35310 49026
rect 35362 48974 35364 49026
rect 35084 48972 35364 48974
rect 35532 49028 35588 51884
rect 35644 50034 35700 52108
rect 36316 52164 36372 52174
rect 36316 52070 36372 52108
rect 35644 49982 35646 50034
rect 35698 49982 35700 50034
rect 35644 49812 35700 49982
rect 35644 49746 35700 49756
rect 35756 52052 35812 52062
rect 35532 48972 35700 49028
rect 35196 48804 35252 48814
rect 34860 48738 34916 48748
rect 35084 48748 35196 48804
rect 34748 48468 34804 48478
rect 34188 48414 34190 48466
rect 34242 48414 34244 48466
rect 34188 48402 34244 48414
rect 34636 48412 34748 48468
rect 33628 48302 33630 48354
rect 33682 48302 33684 48354
rect 33628 48290 33684 48302
rect 34076 48242 34132 48254
rect 34076 48190 34078 48242
rect 34130 48190 34132 48242
rect 32284 48132 32340 48142
rect 32284 48038 32340 48076
rect 33180 48130 33236 48142
rect 33180 48078 33182 48130
rect 33234 48078 33236 48130
rect 32620 47348 32676 47358
rect 32620 47254 32676 47292
rect 33180 47012 33236 48078
rect 33180 46946 33236 46956
rect 33964 48130 34020 48142
rect 33964 48078 33966 48130
rect 34018 48078 34020 48130
rect 33404 46900 33460 46910
rect 33404 46806 33460 46844
rect 32396 44324 32452 44334
rect 32396 44230 32452 44268
rect 32844 44100 32900 44110
rect 32844 44006 32900 44044
rect 33180 43652 33236 43662
rect 32396 43538 32452 43550
rect 32396 43486 32398 43538
rect 32450 43486 32452 43538
rect 32284 43092 32340 43102
rect 32284 42866 32340 43036
rect 32284 42814 32286 42866
rect 32338 42814 32340 42866
rect 32284 42802 32340 42814
rect 32396 42532 32452 43486
rect 33068 43428 33124 43438
rect 33068 42866 33124 43372
rect 33068 42814 33070 42866
rect 33122 42814 33124 42866
rect 33068 42802 33124 42814
rect 33180 43426 33236 43596
rect 33180 43374 33182 43426
rect 33234 43374 33236 43426
rect 32396 42466 32452 42476
rect 32732 42530 32788 42542
rect 32732 42478 32734 42530
rect 32786 42478 32788 42530
rect 32284 41860 32340 41870
rect 32732 41860 32788 42478
rect 33180 42532 33236 43374
rect 33180 42466 33236 42476
rect 32340 41804 32788 41860
rect 32284 41766 32340 41804
rect 32172 41346 32228 41356
rect 32732 41300 32788 41804
rect 32732 41234 32788 41244
rect 33628 39842 33684 39854
rect 33628 39790 33630 39842
rect 33682 39790 33684 39842
rect 32508 39732 32564 39742
rect 32508 39638 32564 39676
rect 31948 39554 32004 39564
rect 33180 39620 33236 39630
rect 31388 39006 31390 39058
rect 31442 39006 31444 39058
rect 31388 38724 31444 39006
rect 31388 38658 31444 38668
rect 31612 39004 32452 39060
rect 31612 38612 31668 39004
rect 32396 38946 32452 39004
rect 32396 38894 32398 38946
rect 32450 38894 32452 38946
rect 32396 38882 32452 38894
rect 33180 38948 33236 39564
rect 33628 39058 33684 39790
rect 33740 39620 33796 39630
rect 33740 39526 33796 39564
rect 33628 39006 33630 39058
rect 33682 39006 33684 39058
rect 33628 38994 33684 39006
rect 33180 38882 33236 38892
rect 31836 38834 31892 38846
rect 31836 38782 31838 38834
rect 31890 38782 31892 38834
rect 31836 38724 31892 38782
rect 32172 38836 32228 38846
rect 32172 38742 32228 38780
rect 32508 38724 32564 38734
rect 33068 38724 33124 38734
rect 32508 38722 33124 38724
rect 32508 38670 32510 38722
rect 32562 38670 33070 38722
rect 33122 38670 33124 38722
rect 32508 38668 33124 38670
rect 33964 38668 34020 48078
rect 34076 47572 34132 48190
rect 34076 47506 34132 47516
rect 34636 46898 34692 48412
rect 34748 48374 34804 48412
rect 34748 47572 34804 47582
rect 34748 47478 34804 47516
rect 34636 46846 34638 46898
rect 34690 46846 34692 46898
rect 34636 46834 34692 46846
rect 35084 47458 35140 48748
rect 35196 48710 35252 48748
rect 35308 48130 35364 48972
rect 35308 48078 35310 48130
rect 35362 48078 35364 48130
rect 35308 48066 35364 48078
rect 35420 48802 35476 48814
rect 35420 48750 35422 48802
rect 35474 48750 35476 48802
rect 35420 48132 35476 48750
rect 35532 48802 35588 48814
rect 35532 48750 35534 48802
rect 35586 48750 35588 48802
rect 35532 48692 35588 48750
rect 35644 48804 35700 48972
rect 35756 49026 35812 51996
rect 36428 50428 36484 55132
rect 38220 54404 38276 54414
rect 38108 54402 38276 54404
rect 38108 54350 38222 54402
rect 38274 54350 38276 54402
rect 38108 54348 38276 54350
rect 36988 53618 37044 53630
rect 36988 53566 36990 53618
rect 37042 53566 37044 53618
rect 36988 52386 37044 53566
rect 37324 53506 37380 53518
rect 37324 53454 37326 53506
rect 37378 53454 37380 53506
rect 37324 53060 37380 53454
rect 37436 53060 37492 53070
rect 37324 53058 37492 53060
rect 37324 53006 37438 53058
rect 37490 53006 37492 53058
rect 37324 53004 37492 53006
rect 37436 52994 37492 53004
rect 36988 52334 36990 52386
rect 37042 52334 37044 52386
rect 36988 52322 37044 52334
rect 37324 52164 37380 52174
rect 36652 52162 37380 52164
rect 36652 52110 37326 52162
rect 37378 52110 37380 52162
rect 36652 52108 37380 52110
rect 36652 51602 36708 52108
rect 36652 51550 36654 51602
rect 36706 51550 36708 51602
rect 36652 51538 36708 51550
rect 35756 48974 35758 49026
rect 35810 48974 35812 49026
rect 35756 48962 35812 48974
rect 36316 50372 36484 50428
rect 35644 48748 35812 48804
rect 35532 48626 35588 48636
rect 35420 48076 35700 48132
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 35084 47406 35086 47458
rect 35138 47406 35140 47458
rect 35084 46900 35140 47406
rect 35532 47684 35588 47694
rect 35532 47458 35588 47628
rect 35532 47406 35534 47458
rect 35586 47406 35588 47458
rect 35532 47394 35588 47406
rect 35084 46806 35140 46844
rect 35308 47234 35364 47246
rect 35308 47182 35310 47234
rect 35362 47182 35364 47234
rect 35308 46562 35364 47182
rect 35420 47236 35476 47246
rect 35420 47234 35588 47236
rect 35420 47182 35422 47234
rect 35474 47182 35588 47234
rect 35420 47180 35588 47182
rect 35420 47170 35476 47180
rect 35308 46510 35310 46562
rect 35362 46510 35364 46562
rect 35308 46452 35364 46510
rect 35308 46386 35364 46396
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 34972 45668 35028 45678
rect 34972 43652 35028 45612
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 34972 43586 35028 43596
rect 34636 43428 34692 43438
rect 34636 43334 34692 43372
rect 34524 43314 34580 43326
rect 34524 43262 34526 43314
rect 34578 43262 34580 43314
rect 34524 42756 34580 43262
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 35532 42980 35588 47180
rect 35644 44324 35700 48076
rect 35756 47458 35812 48748
rect 36204 48802 36260 48814
rect 36204 48750 36206 48802
rect 36258 48750 36260 48802
rect 36204 48692 36260 48750
rect 36204 47684 36260 48636
rect 36204 47618 36260 47628
rect 35756 47406 35758 47458
rect 35810 47406 35812 47458
rect 35756 47394 35812 47406
rect 36204 47458 36260 47470
rect 36204 47406 36206 47458
rect 36258 47406 36260 47458
rect 36204 47348 36260 47406
rect 36204 47282 36260 47292
rect 35644 44268 35812 44324
rect 35532 42914 35588 42924
rect 35644 44100 35700 44110
rect 34524 42690 34580 42700
rect 35196 42644 35252 42654
rect 34860 42642 35252 42644
rect 34860 42590 35198 42642
rect 35250 42590 35252 42642
rect 34860 42588 35252 42590
rect 34860 42194 34916 42588
rect 35196 42578 35252 42588
rect 34860 42142 34862 42194
rect 34914 42142 34916 42194
rect 34860 42130 34916 42142
rect 35308 42196 35364 42206
rect 34636 41972 34692 41982
rect 34636 41970 35028 41972
rect 34636 41918 34638 41970
rect 34690 41918 35028 41970
rect 34636 41916 35028 41918
rect 34636 41906 34692 41916
rect 34972 41410 35028 41916
rect 35308 41858 35364 42140
rect 35308 41806 35310 41858
rect 35362 41806 35364 41858
rect 35308 41794 35364 41806
rect 35644 41636 35700 44044
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 35532 41580 35700 41636
rect 34972 41358 34974 41410
rect 35026 41358 35028 41410
rect 34972 41346 35028 41358
rect 35308 41300 35364 41310
rect 35532 41300 35588 41580
rect 35756 41524 35812 44268
rect 35868 43652 35924 43662
rect 35868 42868 35924 43596
rect 35868 42754 35924 42812
rect 35868 42702 35870 42754
rect 35922 42702 35924 42754
rect 35868 42690 35924 42702
rect 35308 41206 35364 41244
rect 35420 41244 35588 41300
rect 35644 41468 35812 41524
rect 35308 40628 35364 40638
rect 35420 40628 35476 41244
rect 35308 40626 35420 40628
rect 35308 40574 35310 40626
rect 35362 40574 35420 40626
rect 35308 40572 35420 40574
rect 34972 40292 35028 40302
rect 34076 39842 34132 39854
rect 34076 39790 34078 39842
rect 34130 39790 34132 39842
rect 34076 39620 34132 39790
rect 34300 39844 34356 39854
rect 34300 39750 34356 39788
rect 34524 39620 34580 39630
rect 34076 39618 34580 39620
rect 34076 39566 34526 39618
rect 34578 39566 34580 39618
rect 34076 39564 34580 39566
rect 34524 39554 34580 39564
rect 34972 39618 35028 40236
rect 35308 40180 35364 40572
rect 35420 40534 35476 40572
rect 35532 41074 35588 41086
rect 35532 41022 35534 41074
rect 35586 41022 35588 41074
rect 34972 39566 34974 39618
rect 35026 39566 35028 39618
rect 34972 39554 35028 39566
rect 35084 40124 35364 40180
rect 35532 40180 35588 41022
rect 35644 40292 35700 41468
rect 35756 41300 35812 41310
rect 35756 40626 35812 41244
rect 36092 41300 36148 41310
rect 36092 41206 36148 41244
rect 36316 41188 36372 50372
rect 36428 47234 36484 47246
rect 36428 47182 36430 47234
rect 36482 47182 36484 47234
rect 36428 46788 36484 47182
rect 36876 47124 36932 52108
rect 37324 52098 37380 52108
rect 37548 52162 37604 52174
rect 37548 52110 37550 52162
rect 37602 52110 37604 52162
rect 37548 52052 37604 52110
rect 37548 51986 37604 51996
rect 38108 52052 38164 54348
rect 38220 54338 38276 54348
rect 38108 51986 38164 51996
rect 38220 53506 38276 53518
rect 38220 53454 38222 53506
rect 38274 53454 38276 53506
rect 38220 52946 38276 53454
rect 38220 52894 38222 52946
rect 38274 52894 38276 52946
rect 38220 52162 38276 52894
rect 38220 52110 38222 52162
rect 38274 52110 38276 52162
rect 38220 50428 38276 52110
rect 37884 50372 38276 50428
rect 37100 49028 37156 49038
rect 37100 49026 37268 49028
rect 37100 48974 37102 49026
rect 37154 48974 37268 49026
rect 37100 48972 37268 48974
rect 37100 48962 37156 48972
rect 37212 47684 37268 48972
rect 37324 48802 37380 48814
rect 37324 48750 37326 48802
rect 37378 48750 37380 48802
rect 37324 48356 37380 48750
rect 37436 48356 37492 48366
rect 37324 48354 37492 48356
rect 37324 48302 37438 48354
rect 37490 48302 37492 48354
rect 37324 48300 37492 48302
rect 37436 48290 37492 48300
rect 37212 47628 37492 47684
rect 37324 47458 37380 47470
rect 37324 47406 37326 47458
rect 37378 47406 37380 47458
rect 36988 47348 37044 47358
rect 36988 47254 37044 47292
rect 37324 47124 37380 47406
rect 37436 47236 37492 47628
rect 37548 47572 37604 47582
rect 37548 47478 37604 47516
rect 37436 47180 37604 47236
rect 36876 47068 37380 47124
rect 36428 46722 36484 46732
rect 37212 47012 37268 47068
rect 36988 46452 37044 46462
rect 36988 46002 37044 46396
rect 36988 45950 36990 46002
rect 37042 45950 37044 46002
rect 36988 45938 37044 45950
rect 37212 45890 37268 46956
rect 37436 46788 37492 46798
rect 37436 46694 37492 46732
rect 37548 46114 37604 47180
rect 37548 46062 37550 46114
rect 37602 46062 37604 46114
rect 37548 46050 37604 46062
rect 37212 45838 37214 45890
rect 37266 45838 37268 45890
rect 36428 45666 36484 45678
rect 36428 45614 36430 45666
rect 36482 45614 36484 45666
rect 36428 45556 36484 45614
rect 37212 45556 37268 45838
rect 36428 45500 37268 45556
rect 36428 42868 36484 42878
rect 36428 42774 36484 42812
rect 36428 42644 36484 42654
rect 36428 41410 36484 42588
rect 36428 41358 36430 41410
rect 36482 41358 36484 41410
rect 36428 41346 36484 41358
rect 36316 41132 36708 41188
rect 35756 40574 35758 40626
rect 35810 40574 35812 40626
rect 35756 40562 35812 40574
rect 35868 41074 35924 41086
rect 35868 41022 35870 41074
rect 35922 41022 35924 41074
rect 35644 40226 35700 40236
rect 31836 38612 32116 38668
rect 32508 38658 32564 38668
rect 33068 38658 33124 38668
rect 31612 37154 31668 38556
rect 31612 37102 31614 37154
rect 31666 37102 31668 37154
rect 31276 36652 31444 36708
rect 31388 36260 31444 36652
rect 31164 35870 31166 35922
rect 31218 35870 31220 35922
rect 31164 35252 31220 35870
rect 31164 35186 31220 35196
rect 31276 36204 31444 36260
rect 31052 34412 31220 34468
rect 31052 34244 31108 34254
rect 30940 34242 31108 34244
rect 30940 34190 31054 34242
rect 31106 34190 31108 34242
rect 30940 34188 31108 34190
rect 31052 34178 31108 34188
rect 30940 34020 30996 34030
rect 30604 34018 30996 34020
rect 30604 33966 30942 34018
rect 30994 33966 30996 34018
rect 30604 33964 30996 33966
rect 30156 32452 30212 32462
rect 30044 32450 30212 32452
rect 30044 32398 30158 32450
rect 30210 32398 30212 32450
rect 30044 32396 30212 32398
rect 28588 32284 28980 32340
rect 28588 31890 28644 32284
rect 28588 31838 28590 31890
rect 28642 31838 28644 31890
rect 28588 31826 28644 31838
rect 29260 32004 29316 32014
rect 29260 31890 29316 31948
rect 29260 31838 29262 31890
rect 29314 31838 29316 31890
rect 29260 31826 29316 31838
rect 30044 32004 30100 32396
rect 30156 32386 30212 32396
rect 30044 30324 30100 31948
rect 30492 30884 30548 30894
rect 30492 30790 30548 30828
rect 28140 29598 28142 29650
rect 28194 29598 28196 29650
rect 28140 29586 28196 29598
rect 29708 30268 30100 30324
rect 29708 29426 29764 30268
rect 29708 29374 29710 29426
rect 29762 29374 29764 29426
rect 29708 29362 29764 29374
rect 29820 30100 29876 30110
rect 29820 29428 29876 30044
rect 30044 29764 30100 30268
rect 30492 30098 30548 30110
rect 30492 30046 30494 30098
rect 30546 30046 30548 30098
rect 30156 29988 30212 29998
rect 30156 29986 30436 29988
rect 30156 29934 30158 29986
rect 30210 29934 30436 29986
rect 30156 29932 30436 29934
rect 30156 29922 30212 29932
rect 30044 29708 30212 29764
rect 27804 29204 27860 29214
rect 27804 29110 27860 29148
rect 27804 28644 27860 28654
rect 28364 28644 28420 28654
rect 27804 28642 28420 28644
rect 27804 28590 27806 28642
rect 27858 28590 28366 28642
rect 28418 28590 28420 28642
rect 27804 28588 28420 28590
rect 27804 28578 27860 28588
rect 28364 28578 28420 28588
rect 29260 28642 29316 28654
rect 29260 28590 29262 28642
rect 29314 28590 29316 28642
rect 28140 28418 28196 28430
rect 28140 28366 28142 28418
rect 28194 28366 28196 28418
rect 28140 27970 28196 28366
rect 28140 27918 28142 27970
rect 28194 27918 28196 27970
rect 28140 27906 28196 27918
rect 29260 28084 29316 28590
rect 27692 27692 28196 27748
rect 27468 27458 27524 27468
rect 28028 27524 28084 27534
rect 26908 27134 26910 27186
rect 26962 27134 26964 27186
rect 26908 26964 26964 27134
rect 26908 26898 26964 26908
rect 26572 26674 26628 26684
rect 26348 26180 26404 26190
rect 26460 26180 26516 26236
rect 26348 26178 26516 26180
rect 26348 26126 26350 26178
rect 26402 26126 26516 26178
rect 26348 26124 26516 26126
rect 26572 26516 26628 26526
rect 26348 26114 26404 26124
rect 26348 25620 26404 25630
rect 26348 25526 26404 25564
rect 26124 25302 26180 25340
rect 26124 24052 26180 24062
rect 26012 24050 26180 24052
rect 26012 23998 26126 24050
rect 26178 23998 26180 24050
rect 26012 23996 26180 23998
rect 25564 23940 25620 23950
rect 25564 23846 25620 23884
rect 25900 23938 25956 23950
rect 25900 23886 25902 23938
rect 25954 23886 25956 23938
rect 25676 23828 25732 23838
rect 25900 23828 25956 23886
rect 25732 23772 25956 23828
rect 25676 23762 25732 23772
rect 25340 23548 25620 23604
rect 25564 23482 25620 23492
rect 25228 23044 25284 23054
rect 25228 22950 25284 22988
rect 26012 23044 26068 23996
rect 26124 23986 26180 23996
rect 26012 22978 26068 22988
rect 25900 19122 25956 19134
rect 25900 19070 25902 19122
rect 25954 19070 25956 19122
rect 25564 17780 25620 17790
rect 25564 17686 25620 17724
rect 25900 17554 25956 19070
rect 26124 17668 26180 17678
rect 25900 17502 25902 17554
rect 25954 17502 25956 17554
rect 25900 17490 25956 17502
rect 26012 17666 26180 17668
rect 26012 17614 26126 17666
rect 26178 17614 26180 17666
rect 26012 17612 26180 17614
rect 25900 17108 25956 17118
rect 26012 17108 26068 17612
rect 26124 17602 26180 17612
rect 25116 17052 25396 17108
rect 23996 15596 24836 15652
rect 23996 15538 24052 15596
rect 23996 15486 23998 15538
rect 24050 15486 24052 15538
rect 23996 15474 24052 15486
rect 24220 15428 24276 15438
rect 24220 15334 24276 15372
rect 24108 15316 24164 15326
rect 24108 15222 24164 15260
rect 24444 15314 24500 15326
rect 24444 15262 24446 15314
rect 24498 15262 24500 15314
rect 24444 15148 24500 15262
rect 24444 15092 24724 15148
rect 24668 14642 24724 15092
rect 24668 14590 24670 14642
rect 24722 14590 24724 14642
rect 24556 13188 24612 13198
rect 24556 13094 24612 13132
rect 24220 12740 24276 12750
rect 24668 12740 24724 14590
rect 24780 13074 24836 15596
rect 25340 15538 25396 17052
rect 25900 17106 26068 17108
rect 25900 17054 25902 17106
rect 25954 17054 26068 17106
rect 25900 17052 26068 17054
rect 26236 17108 26292 17118
rect 25900 17042 25956 17052
rect 26236 16882 26292 17052
rect 26236 16830 26238 16882
rect 26290 16830 26292 16882
rect 26236 16818 26292 16830
rect 25676 16772 25732 16782
rect 26460 16772 26516 16782
rect 25676 16210 25732 16716
rect 25676 16158 25678 16210
rect 25730 16158 25732 16210
rect 25676 16146 25732 16158
rect 26348 16770 26516 16772
rect 26348 16718 26462 16770
rect 26514 16718 26516 16770
rect 26348 16716 26516 16718
rect 25340 15486 25342 15538
rect 25394 15486 25396 15538
rect 25340 15428 25396 15486
rect 25340 15148 25396 15372
rect 26012 15540 26068 15550
rect 26012 15314 26068 15484
rect 26012 15262 26014 15314
rect 26066 15262 26068 15314
rect 26012 15148 26068 15262
rect 25340 15092 25508 15148
rect 25452 14644 25508 15092
rect 25900 15092 26068 15148
rect 26236 15540 26292 15550
rect 26348 15540 26404 16716
rect 26460 16706 26516 16716
rect 26236 15538 26404 15540
rect 26236 15486 26238 15538
rect 26290 15486 26404 15538
rect 26236 15484 26404 15486
rect 25900 14754 25956 15092
rect 25900 14702 25902 14754
rect 25954 14702 25956 14754
rect 25452 14642 25844 14644
rect 25452 14590 25454 14642
rect 25506 14590 25844 14642
rect 25452 14588 25844 14590
rect 25452 14578 25508 14588
rect 25340 13634 25396 13646
rect 25340 13582 25342 13634
rect 25394 13582 25396 13634
rect 25340 13524 25396 13582
rect 24780 13022 24782 13074
rect 24834 13022 24836 13074
rect 24780 13010 24836 13022
rect 25116 13468 25396 13524
rect 24220 12738 24388 12740
rect 24220 12686 24222 12738
rect 24274 12686 24388 12738
rect 24220 12684 24388 12686
rect 24220 12674 24276 12684
rect 23772 12292 23828 12302
rect 23772 12178 23828 12236
rect 24220 12292 24276 12302
rect 24220 12198 24276 12236
rect 23772 12126 23774 12178
rect 23826 12126 23828 12178
rect 23772 12114 23828 12126
rect 24332 11394 24388 12684
rect 24332 11342 24334 11394
rect 24386 11342 24388 11394
rect 24332 11330 24388 11342
rect 24444 12684 24724 12740
rect 24108 11172 24164 11182
rect 23884 11170 24164 11172
rect 23884 11118 24110 11170
rect 24162 11118 24164 11170
rect 23884 11116 24164 11118
rect 22876 10892 23492 10948
rect 22876 10836 22932 10892
rect 22428 10782 22430 10834
rect 22482 10782 22484 10834
rect 22428 10770 22484 10782
rect 22540 10834 22932 10836
rect 22540 10782 22878 10834
rect 22930 10782 22932 10834
rect 22540 10780 22932 10782
rect 22092 10612 22148 10622
rect 22540 10612 22596 10780
rect 22876 10770 22932 10780
rect 22092 10610 22596 10612
rect 22092 10558 22094 10610
rect 22146 10558 22596 10610
rect 22092 10556 22596 10558
rect 22092 10546 22148 10556
rect 21868 10500 21924 10510
rect 21644 10498 21924 10500
rect 21644 10446 21870 10498
rect 21922 10446 21924 10498
rect 21644 10444 21924 10446
rect 21868 10164 21924 10444
rect 21868 10098 21924 10108
rect 23100 9826 23156 9838
rect 23100 9774 23102 9826
rect 23154 9774 23156 9826
rect 21756 9604 21812 9614
rect 21084 9212 21364 9268
rect 20524 9156 20580 9166
rect 20524 9154 21252 9156
rect 20524 9102 20526 9154
rect 20578 9102 21252 9154
rect 20524 9100 21252 9102
rect 20524 9090 20580 9100
rect 21196 7586 21252 9100
rect 21196 7534 21198 7586
rect 21250 7534 21252 7586
rect 21196 7522 21252 7534
rect 20468 7308 20692 7364
rect 20412 7298 20468 7308
rect 20188 5282 20244 5292
rect 20412 6692 20468 6702
rect 20412 5346 20468 6636
rect 20412 5294 20414 5346
rect 20466 5294 20468 5346
rect 19740 5236 19796 5246
rect 19740 5142 19796 5180
rect 20412 5236 20468 5294
rect 20412 5170 20468 5180
rect 20636 5234 20692 7308
rect 21308 6692 21364 9212
rect 21308 6626 21364 6636
rect 21756 5796 21812 9548
rect 21980 7474 22036 7486
rect 21980 7422 21982 7474
rect 22034 7422 22036 7474
rect 21980 7364 22036 7422
rect 22428 7364 22484 7374
rect 23100 7364 23156 9774
rect 21980 7362 23156 7364
rect 21980 7310 22430 7362
rect 22482 7310 23156 7362
rect 21980 7308 23156 7310
rect 21868 6466 21924 6478
rect 21868 6414 21870 6466
rect 21922 6414 21924 6466
rect 21868 5908 21924 6414
rect 22316 6466 22372 7308
rect 22428 7298 22484 7308
rect 23436 6692 23492 10892
rect 23884 9938 23940 11116
rect 24108 11106 24164 11116
rect 24220 10836 24276 10846
rect 24220 10742 24276 10780
rect 23884 9886 23886 9938
rect 23938 9886 23940 9938
rect 23884 9874 23940 9886
rect 23548 6692 23604 6702
rect 22316 6414 22318 6466
rect 22370 6414 22372 6466
rect 22204 5908 22260 5918
rect 21868 5906 22260 5908
rect 21868 5854 22206 5906
rect 22258 5854 22260 5906
rect 21868 5852 22260 5854
rect 20636 5182 20638 5234
rect 20690 5182 20692 5234
rect 20636 5170 20692 5182
rect 21308 5794 21812 5796
rect 21308 5742 21758 5794
rect 21810 5742 21812 5794
rect 21308 5740 21812 5742
rect 21308 5234 21364 5740
rect 21756 5730 21812 5740
rect 22204 5572 22260 5852
rect 22204 5506 22260 5516
rect 22316 5908 22372 6414
rect 21532 5348 21588 5358
rect 21532 5254 21588 5292
rect 22316 5348 22372 5852
rect 23212 6690 23604 6692
rect 23212 6638 23550 6690
rect 23602 6638 23604 6690
rect 23212 6636 23604 6638
rect 23212 5908 23268 6636
rect 23548 6626 23604 6636
rect 23212 5794 23268 5852
rect 24220 5908 24276 5918
rect 24220 5814 24276 5852
rect 24444 5906 24500 12684
rect 25116 12292 25172 13468
rect 25228 13188 25284 13198
rect 25228 13074 25284 13132
rect 25228 13022 25230 13074
rect 25282 13022 25284 13074
rect 25228 13010 25284 13022
rect 25116 12226 25172 12236
rect 25228 12180 25284 12190
rect 24668 10612 24724 10622
rect 24668 10518 24724 10556
rect 25228 10500 25284 12124
rect 25788 11508 25844 14588
rect 25900 14642 25956 14702
rect 25900 14590 25902 14642
rect 25954 14590 25956 14642
rect 25900 14578 25956 14590
rect 25900 11508 25956 11518
rect 26236 11508 26292 15484
rect 26460 15428 26516 15438
rect 26460 15334 26516 15372
rect 26348 15202 26404 15214
rect 26348 15150 26350 15202
rect 26402 15150 26404 15202
rect 26348 15148 26404 15150
rect 26572 15148 26628 26460
rect 27132 26404 27188 26414
rect 27020 25394 27076 25406
rect 27020 25342 27022 25394
rect 27074 25342 27076 25394
rect 26684 25284 26740 25294
rect 26684 25190 26740 25228
rect 27020 25284 27076 25342
rect 27020 25218 27076 25228
rect 26796 25172 26852 25182
rect 26684 20580 26740 20590
rect 26684 20020 26740 20524
rect 26684 19954 26740 19964
rect 26684 19236 26740 19246
rect 26684 19142 26740 19180
rect 26684 17442 26740 17454
rect 26684 17390 26686 17442
rect 26738 17390 26740 17442
rect 26684 16996 26740 17390
rect 26684 16930 26740 16940
rect 26796 16772 26852 25116
rect 27020 24724 27076 24734
rect 27020 24630 27076 24668
rect 27132 22482 27188 26348
rect 27804 25732 27860 25742
rect 27356 25284 27412 25294
rect 27804 25284 27860 25676
rect 27356 25282 27748 25284
rect 27356 25230 27358 25282
rect 27410 25230 27748 25282
rect 27356 25228 27748 25230
rect 27356 25218 27412 25228
rect 27692 24836 27748 25228
rect 27804 25190 27860 25228
rect 27804 24836 27860 24846
rect 27692 24834 27860 24836
rect 27692 24782 27806 24834
rect 27858 24782 27860 24834
rect 27692 24780 27860 24782
rect 27804 24770 27860 24780
rect 27916 23826 27972 23838
rect 27916 23774 27918 23826
rect 27970 23774 27972 23826
rect 27580 23716 27636 23726
rect 27356 23714 27636 23716
rect 27356 23662 27582 23714
rect 27634 23662 27636 23714
rect 27356 23660 27636 23662
rect 27356 23266 27412 23660
rect 27580 23650 27636 23660
rect 27916 23380 27972 23774
rect 27916 23314 27972 23324
rect 27356 23214 27358 23266
rect 27410 23214 27412 23266
rect 27356 23202 27412 23214
rect 28028 23268 28084 27468
rect 28028 23156 28084 23212
rect 27132 22430 27134 22482
rect 27186 22430 27188 22482
rect 27020 20916 27076 20926
rect 27132 20916 27188 22430
rect 27692 23154 28084 23156
rect 27692 23102 28030 23154
rect 28082 23102 28084 23154
rect 27692 23100 28084 23102
rect 27692 22482 27748 23100
rect 28028 23090 28084 23100
rect 27692 22430 27694 22482
rect 27746 22430 27748 22482
rect 27692 22418 27748 22430
rect 27020 20914 27188 20916
rect 27020 20862 27022 20914
rect 27074 20862 27188 20914
rect 27020 20860 27188 20862
rect 27020 20850 27076 20860
rect 27244 20802 27300 20814
rect 28140 20804 28196 27692
rect 29260 27524 29316 28028
rect 29260 27458 29316 27468
rect 29820 27188 29876 29372
rect 30044 28868 30100 28878
rect 30044 28754 30100 28812
rect 30044 28702 30046 28754
rect 30098 28702 30100 28754
rect 30044 28690 30100 28702
rect 30156 28084 30212 29708
rect 30380 29538 30436 29932
rect 30380 29486 30382 29538
rect 30434 29486 30436 29538
rect 30380 29474 30436 29486
rect 30380 28868 30436 28878
rect 30492 28868 30548 30046
rect 30380 28866 30548 28868
rect 30380 28814 30382 28866
rect 30434 28814 30548 28866
rect 30380 28812 30548 28814
rect 30380 28802 30436 28812
rect 30156 28018 30212 28028
rect 30268 27746 30324 27758
rect 30268 27694 30270 27746
rect 30322 27694 30324 27746
rect 30268 27636 30324 27694
rect 30492 27636 30548 27646
rect 30268 27634 30548 27636
rect 30268 27582 30494 27634
rect 30546 27582 30548 27634
rect 30268 27580 30548 27582
rect 30492 27570 30548 27580
rect 29932 27298 29988 27310
rect 29932 27246 29934 27298
rect 29986 27246 29988 27298
rect 29932 27188 29988 27246
rect 29820 27186 29988 27188
rect 29820 27134 29934 27186
rect 29986 27134 29988 27186
rect 29820 27132 29988 27134
rect 29932 27122 29988 27132
rect 30380 26964 30436 27002
rect 30380 26898 30436 26908
rect 30156 25282 30212 25294
rect 30156 25230 30158 25282
rect 30210 25230 30212 25282
rect 30156 24948 30212 25230
rect 30492 25284 30548 25294
rect 29820 24892 30212 24948
rect 30268 25172 30324 25182
rect 29708 24724 29764 24734
rect 29820 24724 29876 24892
rect 30268 24836 30324 25116
rect 29764 24668 29876 24724
rect 29932 24834 30324 24836
rect 29932 24782 30270 24834
rect 30322 24782 30324 24834
rect 29932 24780 30324 24782
rect 29708 23940 29764 24668
rect 29932 24610 29988 24780
rect 30268 24770 30324 24780
rect 29932 24558 29934 24610
rect 29986 24558 29988 24610
rect 29932 24546 29988 24558
rect 30492 24498 30548 25228
rect 30492 24446 30494 24498
rect 30546 24446 30548 24498
rect 30492 24276 30548 24446
rect 30268 24220 30548 24276
rect 29708 23846 29764 23884
rect 29820 24052 29876 24062
rect 29148 23492 29204 23502
rect 28588 23268 28644 23278
rect 28588 23174 28644 23212
rect 27244 20750 27246 20802
rect 27298 20750 27300 20802
rect 27244 20580 27300 20750
rect 28028 20748 28196 20804
rect 27244 20514 27300 20524
rect 27580 20580 27636 20590
rect 27580 20578 27860 20580
rect 27580 20526 27582 20578
rect 27634 20526 27860 20578
rect 27580 20524 27860 20526
rect 27580 20514 27636 20524
rect 27804 20130 27860 20524
rect 27804 20078 27806 20130
rect 27858 20078 27860 20130
rect 27804 20066 27860 20078
rect 27132 19236 27188 19246
rect 27132 19010 27188 19180
rect 27132 18958 27134 19010
rect 27186 18958 27188 19010
rect 27132 18452 27188 18958
rect 27692 18452 27748 18462
rect 27132 18450 27748 18452
rect 27132 18398 27694 18450
rect 27746 18398 27748 18450
rect 27132 18396 27748 18398
rect 27692 17780 27748 18396
rect 26908 17108 26964 17118
rect 26908 17014 26964 17052
rect 27692 16996 27748 17724
rect 27692 16930 27748 16940
rect 26796 16706 26852 16716
rect 27804 15988 27860 15998
rect 27356 15986 27860 15988
rect 27356 15934 27806 15986
rect 27858 15934 27860 15986
rect 27356 15932 27860 15934
rect 27356 15538 27412 15932
rect 27804 15922 27860 15932
rect 28028 15876 28084 20748
rect 28140 20132 28196 20142
rect 28140 20130 28420 20132
rect 28140 20078 28142 20130
rect 28194 20078 28420 20130
rect 28140 20076 28420 20078
rect 28140 20066 28196 20076
rect 28364 18562 28420 20076
rect 29148 19348 29204 23436
rect 29260 23380 29316 23390
rect 29260 23286 29316 23324
rect 29820 23154 29876 23996
rect 29820 23102 29822 23154
rect 29874 23102 29876 23154
rect 29820 23090 29876 23102
rect 29596 22930 29652 22942
rect 29596 22878 29598 22930
rect 29650 22878 29652 22930
rect 29260 22148 29316 22158
rect 29596 22148 29652 22878
rect 29260 22146 29652 22148
rect 29260 22094 29262 22146
rect 29314 22094 29652 22146
rect 29260 22092 29652 22094
rect 29260 20580 29316 22092
rect 29596 21476 29652 21486
rect 29596 21382 29652 21420
rect 29260 20514 29316 20524
rect 29708 19460 29764 19470
rect 29260 19348 29316 19358
rect 29148 19292 29260 19348
rect 29260 19254 29316 19292
rect 29708 19346 29764 19404
rect 29708 19294 29710 19346
rect 29762 19294 29764 19346
rect 29708 19282 29764 19294
rect 28364 18510 28366 18562
rect 28418 18510 28420 18562
rect 28364 18498 28420 18510
rect 28028 15810 28084 15820
rect 28588 17780 28644 17790
rect 28588 16098 28644 17724
rect 29260 17780 29316 17790
rect 29260 17106 29316 17724
rect 30044 17780 30100 17790
rect 30044 17686 30100 17724
rect 30268 17108 30324 24220
rect 30492 23828 30548 23838
rect 30492 23734 30548 23772
rect 30604 23548 30660 33964
rect 30940 33954 30996 33964
rect 31164 33460 31220 34412
rect 31276 34242 31332 36204
rect 31612 35700 31668 37102
rect 31836 36482 31892 36494
rect 31836 36430 31838 36482
rect 31890 36430 31892 36482
rect 31836 36260 31892 36430
rect 31836 36194 31892 36204
rect 31612 35644 32004 35700
rect 31836 35476 31892 35486
rect 31388 35474 31892 35476
rect 31388 35422 31838 35474
rect 31890 35422 31892 35474
rect 31388 35420 31892 35422
rect 31388 34914 31444 35420
rect 31836 35410 31892 35420
rect 31948 35252 32004 35644
rect 31836 35196 32004 35252
rect 31836 35028 31892 35196
rect 31388 34862 31390 34914
rect 31442 34862 31444 34914
rect 31388 34850 31444 34862
rect 31724 34972 31892 35028
rect 31612 34804 31668 34814
rect 31612 34710 31668 34748
rect 31276 34190 31278 34242
rect 31330 34190 31332 34242
rect 31276 34178 31332 34190
rect 31500 34132 31556 34142
rect 31500 34038 31556 34076
rect 31500 33572 31556 33582
rect 31276 33460 31332 33470
rect 31164 33458 31332 33460
rect 31164 33406 31278 33458
rect 31330 33406 31332 33458
rect 31164 33404 31332 33406
rect 31276 33394 31332 33404
rect 31500 33348 31556 33516
rect 30940 33124 30996 33134
rect 31500 33124 31556 33292
rect 30940 33122 31556 33124
rect 30940 33070 30942 33122
rect 30994 33070 31556 33122
rect 30940 33068 31556 33070
rect 30940 32340 30996 33068
rect 30940 32274 30996 32284
rect 30716 30884 30772 30894
rect 31276 30884 31332 30894
rect 30716 29652 30772 30828
rect 31164 30882 31332 30884
rect 31164 30830 31278 30882
rect 31330 30830 31332 30882
rect 31164 30828 31332 30830
rect 31164 30436 31220 30828
rect 31276 30818 31332 30828
rect 31612 30884 31668 30894
rect 31724 30884 31780 34972
rect 31948 34914 32004 34926
rect 31948 34862 31950 34914
rect 32002 34862 32004 34914
rect 31948 34580 32004 34862
rect 31948 34514 32004 34524
rect 31948 34356 32004 34366
rect 31948 34262 32004 34300
rect 31836 33122 31892 33134
rect 31836 33070 31838 33122
rect 31890 33070 31892 33122
rect 31836 32676 31892 33070
rect 31836 32610 31892 32620
rect 31948 31220 32004 31230
rect 32060 31220 32116 38612
rect 33292 38610 33348 38622
rect 33292 38558 33294 38610
rect 33346 38558 33348 38610
rect 33292 38276 33348 38558
rect 32284 38220 33348 38276
rect 33628 38612 34020 38668
rect 32172 35588 32228 35598
rect 32172 35474 32228 35532
rect 32172 35422 32174 35474
rect 32226 35422 32228 35474
rect 32172 33572 32228 35422
rect 32172 33506 32228 33516
rect 31948 31218 32116 31220
rect 31948 31166 31950 31218
rect 32002 31166 32116 31218
rect 31948 31164 32116 31166
rect 31948 31154 32004 31164
rect 31668 30828 31780 30884
rect 31612 30818 31668 30828
rect 31836 30436 31892 30446
rect 31164 30434 31892 30436
rect 31164 30382 31838 30434
rect 31890 30382 31892 30434
rect 31164 30380 31892 30382
rect 30828 30100 30884 30110
rect 30828 30006 30884 30044
rect 30716 29586 30772 29596
rect 31052 29986 31108 29998
rect 31052 29934 31054 29986
rect 31106 29934 31108 29986
rect 30716 28868 30772 28878
rect 30716 28774 30772 28812
rect 30940 28756 30996 28766
rect 31052 28756 31108 29934
rect 31164 28868 31220 30380
rect 31836 30370 31892 30380
rect 31612 30212 31668 30222
rect 31612 30118 31668 30156
rect 32060 30100 32116 31164
rect 32172 33234 32228 33246
rect 32172 33182 32174 33234
rect 32226 33182 32228 33234
rect 32172 30210 32228 33182
rect 32172 30158 32174 30210
rect 32226 30158 32228 30210
rect 32172 30146 32228 30158
rect 31276 29986 31332 29998
rect 31276 29934 31278 29986
rect 31330 29934 31332 29986
rect 31276 29652 31332 29934
rect 31388 29988 31444 29998
rect 31388 29986 31892 29988
rect 31388 29934 31390 29986
rect 31442 29934 31892 29986
rect 31388 29932 31892 29934
rect 31388 29922 31444 29932
rect 31276 29586 31332 29596
rect 31164 28802 31220 28812
rect 30940 28754 31108 28756
rect 30940 28702 30942 28754
rect 30994 28702 31108 28754
rect 30940 28700 31108 28702
rect 31836 28754 31892 29932
rect 32060 28868 32116 30044
rect 32060 28812 32228 28868
rect 31836 28702 31838 28754
rect 31890 28702 31892 28754
rect 30716 28084 30772 28094
rect 30716 27990 30772 28028
rect 30828 27636 30884 27646
rect 30940 27636 30996 28700
rect 31836 28690 31892 28702
rect 32060 28644 32116 28654
rect 31948 28642 32116 28644
rect 31948 28590 32062 28642
rect 32114 28590 32116 28642
rect 31948 28588 32116 28590
rect 31948 28532 32004 28588
rect 32060 28578 32116 28588
rect 31612 28476 32004 28532
rect 31500 27748 31556 27758
rect 30828 27634 30996 27636
rect 30828 27582 30830 27634
rect 30882 27582 30996 27634
rect 30828 27580 30996 27582
rect 31388 27692 31500 27748
rect 30828 27570 30884 27580
rect 30716 27298 30772 27310
rect 30716 27246 30718 27298
rect 30770 27246 30772 27298
rect 30716 27076 30772 27246
rect 30828 27076 30884 27086
rect 30716 27074 30884 27076
rect 30716 27022 30830 27074
rect 30882 27022 30884 27074
rect 30716 27020 30884 27022
rect 30828 27010 30884 27020
rect 31388 26964 31444 27692
rect 31500 27654 31556 27692
rect 31500 27300 31556 27310
rect 31612 27300 31668 28476
rect 31500 27298 31668 27300
rect 31500 27246 31502 27298
rect 31554 27246 31668 27298
rect 31500 27244 31668 27246
rect 32060 27972 32116 27982
rect 32172 27972 32228 28812
rect 32284 28644 32340 38220
rect 33404 38050 33460 38062
rect 33404 37998 33406 38050
rect 33458 37998 33460 38050
rect 32620 37938 32676 37950
rect 32620 37886 32622 37938
rect 32674 37886 32676 37938
rect 32396 35812 32452 35822
rect 32396 35698 32452 35756
rect 32396 35646 32398 35698
rect 32450 35646 32452 35698
rect 32396 35634 32452 35646
rect 32508 33236 32564 33246
rect 32620 33236 32676 37886
rect 33404 37828 33460 37998
rect 33404 37762 33460 37772
rect 32844 36260 32900 36270
rect 32844 35476 32900 36204
rect 32956 35588 33012 35598
rect 33180 35588 33236 35598
rect 33012 35586 33236 35588
rect 33012 35534 33182 35586
rect 33234 35534 33236 35586
rect 33012 35532 33236 35534
rect 32956 35522 33012 35532
rect 33180 35522 33236 35532
rect 32844 35410 32900 35420
rect 32732 34804 32788 34814
rect 32732 34710 32788 34748
rect 33404 34356 33460 34366
rect 33404 34262 33460 34300
rect 33068 33572 33124 33582
rect 33068 33478 33124 33516
rect 33292 33348 33348 33358
rect 32508 33234 32676 33236
rect 32508 33182 32510 33234
rect 32562 33182 32676 33234
rect 32508 33180 32676 33182
rect 32732 33346 33348 33348
rect 32732 33294 33294 33346
rect 33346 33294 33348 33346
rect 32732 33292 33348 33294
rect 33628 33348 33684 38612
rect 33852 37828 33908 37838
rect 33852 37044 33908 37772
rect 33852 36978 33908 36988
rect 35084 35922 35140 40124
rect 35532 40114 35588 40124
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35868 39956 35924 41022
rect 35196 39946 35460 39956
rect 35532 39900 35924 39956
rect 35196 39732 35252 39742
rect 35196 39506 35252 39676
rect 35308 39620 35364 39630
rect 35308 39526 35364 39564
rect 35196 39454 35198 39506
rect 35250 39454 35252 39506
rect 35196 39442 35252 39454
rect 35532 39396 35588 39900
rect 35756 39732 35812 39742
rect 35756 39638 35812 39676
rect 35868 39618 35924 39900
rect 35868 39566 35870 39618
rect 35922 39566 35924 39618
rect 35868 39554 35924 39566
rect 36092 40628 36148 40638
rect 36092 39618 36148 40572
rect 36092 39566 36094 39618
rect 36146 39566 36148 39618
rect 36092 39554 36148 39566
rect 36204 40180 36260 40190
rect 36204 39618 36260 40124
rect 36204 39566 36206 39618
rect 36258 39566 36260 39618
rect 35308 39340 35588 39396
rect 35756 39394 35812 39406
rect 35756 39342 35758 39394
rect 35810 39342 35812 39394
rect 35308 38722 35364 39340
rect 35308 38670 35310 38722
rect 35362 38670 35364 38722
rect 35308 38658 35364 38670
rect 35532 39172 35588 39182
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 35532 38162 35588 39116
rect 35532 38110 35534 38162
rect 35586 38110 35588 38162
rect 35532 38098 35588 38110
rect 35756 37268 35812 39342
rect 35532 37212 35812 37268
rect 35308 37156 35364 37166
rect 35308 37062 35364 37100
rect 35532 37044 35588 37212
rect 35868 37156 35924 37166
rect 36204 37156 36260 39566
rect 36428 39620 36484 39630
rect 36428 38668 36484 39564
rect 36428 38612 36596 38668
rect 36428 38052 36484 38062
rect 36428 37958 36484 37996
rect 35924 37100 36260 37156
rect 36428 37156 36484 37166
rect 35868 37090 35924 37100
rect 35532 36988 35700 37044
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35084 35870 35086 35922
rect 35138 35870 35140 35922
rect 33740 35252 33796 35262
rect 33740 34804 33796 35196
rect 34860 35026 34916 35038
rect 34860 34974 34862 35026
rect 34914 34974 34916 35026
rect 33740 34354 33796 34748
rect 33740 34302 33742 34354
rect 33794 34302 33796 34354
rect 33740 34290 33796 34302
rect 34076 34916 34132 34926
rect 34076 34356 34132 34860
rect 34076 34262 34132 34300
rect 34524 34692 34580 34702
rect 34524 34354 34580 34636
rect 34524 34302 34526 34354
rect 34578 34302 34580 34354
rect 34524 34290 34580 34302
rect 33852 34130 33908 34142
rect 33852 34078 33854 34130
rect 33906 34078 33908 34130
rect 33740 33348 33796 33358
rect 33628 33346 33796 33348
rect 33628 33294 33742 33346
rect 33794 33294 33796 33346
rect 33628 33292 33796 33294
rect 32508 33170 32564 33180
rect 32396 30884 32452 30894
rect 32396 30790 32452 30828
rect 32732 30660 32788 33292
rect 33292 33282 33348 33292
rect 33740 33282 33796 33292
rect 33068 32676 33124 32686
rect 33068 32582 33124 32620
rect 33404 32676 33460 32686
rect 33404 32674 33572 32676
rect 33404 32622 33406 32674
rect 33458 32622 33572 32674
rect 33404 32620 33572 32622
rect 33404 32610 33460 32620
rect 33516 31780 33572 32620
rect 33852 32004 33908 34078
rect 34300 34130 34356 34142
rect 34300 34078 34302 34130
rect 34354 34078 34356 34130
rect 33964 34018 34020 34030
rect 33964 33966 33966 34018
rect 34018 33966 34020 34018
rect 33964 33234 34020 33966
rect 34300 33460 34356 34078
rect 34300 33394 34356 33404
rect 34748 34130 34804 34142
rect 34748 34078 34750 34130
rect 34802 34078 34804 34130
rect 33964 33182 33966 33234
rect 34018 33182 34020 33234
rect 33964 33170 34020 33182
rect 34076 33346 34132 33358
rect 34076 33294 34078 33346
rect 34130 33294 34132 33346
rect 33852 31938 33908 31948
rect 33516 31724 33908 31780
rect 33852 31106 33908 31724
rect 33852 31054 33854 31106
rect 33906 31054 33908 31106
rect 33852 31042 33908 31054
rect 33180 30994 33236 31006
rect 33180 30942 33182 30994
rect 33234 30942 33236 30994
rect 32396 30604 32788 30660
rect 32956 30884 33012 30894
rect 33180 30884 33236 30942
rect 33516 30884 33572 30894
rect 33180 30828 33516 30884
rect 32396 28866 32452 30604
rect 32732 30212 32788 30222
rect 32620 30156 32732 30212
rect 32508 30100 32564 30110
rect 32508 30006 32564 30044
rect 32508 29316 32564 29326
rect 32620 29316 32676 30156
rect 32732 30118 32788 30156
rect 32956 30098 33012 30828
rect 32956 30046 32958 30098
rect 33010 30046 33012 30098
rect 32956 30034 33012 30046
rect 33068 29986 33124 29998
rect 33068 29934 33070 29986
rect 33122 29934 33124 29986
rect 33068 29426 33124 29934
rect 33068 29374 33070 29426
rect 33122 29374 33124 29426
rect 33068 29362 33124 29374
rect 32508 29314 32676 29316
rect 32508 29262 32510 29314
rect 32562 29262 32676 29314
rect 32508 29260 32676 29262
rect 32508 29250 32564 29260
rect 33292 29204 33348 29214
rect 32396 28814 32398 28866
rect 32450 28814 32452 28866
rect 32396 28802 32452 28814
rect 32620 29202 33348 29204
rect 32620 29150 33294 29202
rect 33346 29150 33348 29202
rect 32620 29148 33348 29150
rect 32284 28588 32452 28644
rect 32060 27970 32228 27972
rect 32060 27918 32062 27970
rect 32114 27918 32228 27970
rect 32060 27916 32228 27918
rect 31500 27234 31556 27244
rect 31836 27188 31892 27198
rect 32060 27188 32116 27916
rect 31836 27186 32116 27188
rect 31836 27134 31838 27186
rect 31890 27134 32116 27186
rect 31836 27132 32116 27134
rect 31836 27122 31892 27132
rect 32060 27074 32116 27132
rect 32060 27022 32062 27074
rect 32114 27022 32116 27074
rect 31444 26908 31780 26964
rect 31388 26898 31444 26908
rect 31164 26850 31220 26862
rect 31164 26798 31166 26850
rect 31218 26798 31220 26850
rect 31052 25284 31108 25294
rect 31052 25190 31108 25228
rect 31164 25172 31220 26798
rect 31724 26514 31780 26908
rect 31724 26462 31726 26514
rect 31778 26462 31780 26514
rect 31724 26450 31780 26462
rect 32060 26514 32116 27022
rect 32284 27858 32340 27870
rect 32284 27806 32286 27858
rect 32338 27806 32340 27858
rect 32284 26908 32340 27806
rect 32396 27186 32452 28588
rect 32620 28082 32676 29148
rect 33292 29138 33348 29148
rect 33404 28980 33460 30828
rect 33516 30818 33572 30828
rect 33628 29652 33684 29662
rect 33852 29652 33908 29662
rect 33628 29650 33852 29652
rect 33628 29598 33630 29650
rect 33682 29598 33852 29650
rect 33628 29596 33852 29598
rect 33628 29586 33684 29596
rect 33852 29586 33908 29596
rect 32620 28030 32622 28082
rect 32674 28030 32676 28082
rect 32620 28018 32676 28030
rect 32844 28924 33460 28980
rect 32844 28754 32900 28924
rect 32844 28702 32846 28754
rect 32898 28702 32900 28754
rect 32844 28084 32900 28702
rect 32844 28018 32900 28028
rect 32508 27970 32564 27982
rect 32508 27918 32510 27970
rect 32562 27918 32564 27970
rect 32508 27748 32564 27918
rect 32564 27692 32676 27748
rect 32508 27682 32564 27692
rect 32396 27134 32398 27186
rect 32450 27134 32452 27186
rect 32396 27122 32452 27134
rect 32060 26462 32062 26514
rect 32114 26462 32116 26514
rect 32060 26450 32116 26462
rect 32172 26852 32340 26908
rect 32620 26962 32676 27692
rect 32620 26910 32622 26962
rect 32674 26910 32676 26962
rect 32620 26898 32676 26910
rect 34076 26908 34132 33294
rect 34748 29652 34804 34078
rect 34860 33460 34916 34974
rect 35084 34916 35140 35870
rect 35532 36708 35588 36718
rect 35532 35586 35588 36652
rect 35532 35534 35534 35586
rect 35586 35534 35588 35586
rect 35532 35474 35588 35534
rect 35532 35422 35534 35474
rect 35586 35422 35588 35474
rect 35532 35410 35588 35422
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35644 35252 35700 36988
rect 36204 36484 36260 36494
rect 36204 36482 36372 36484
rect 36204 36430 36206 36482
rect 36258 36430 36372 36482
rect 36204 36428 36372 36430
rect 36204 36418 36260 36428
rect 35756 36260 35812 36270
rect 35756 36258 35924 36260
rect 35756 36206 35758 36258
rect 35810 36206 35924 36258
rect 35756 36204 35924 36206
rect 35756 36194 35812 36204
rect 35644 35186 35700 35196
rect 35756 35812 35812 35822
rect 35084 34850 35140 34860
rect 35420 35028 35476 35038
rect 35196 34244 35252 34254
rect 35196 34150 35252 34188
rect 35420 34242 35476 34972
rect 35644 35028 35700 35066
rect 35644 34962 35700 34972
rect 35532 34804 35588 34814
rect 35532 34710 35588 34748
rect 35644 34692 35700 34702
rect 35756 34692 35812 35756
rect 35868 35588 35924 36204
rect 36316 35924 36372 36428
rect 36428 36370 36484 37100
rect 36428 36318 36430 36370
rect 36482 36318 36484 36370
rect 36428 36306 36484 36318
rect 36428 35924 36484 35934
rect 36316 35922 36484 35924
rect 36316 35870 36430 35922
rect 36482 35870 36484 35922
rect 36316 35868 36484 35870
rect 36428 35858 36484 35868
rect 36092 35588 36148 35598
rect 35868 35532 36092 35588
rect 35980 35364 36036 35374
rect 35868 34916 35924 34926
rect 35868 34822 35924 34860
rect 35980 34914 36036 35308
rect 35980 34862 35982 34914
rect 36034 34862 36036 34914
rect 35644 34690 35812 34692
rect 35644 34638 35646 34690
rect 35698 34638 35812 34690
rect 35644 34636 35812 34638
rect 35644 34356 35700 34636
rect 35644 34290 35700 34300
rect 35420 34190 35422 34242
rect 35474 34190 35476 34242
rect 35420 34178 35476 34190
rect 35980 34132 36036 34862
rect 35644 34076 36036 34132
rect 35532 34020 35588 34030
rect 35532 33926 35588 33964
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 34860 33394 34916 33404
rect 35308 33460 35364 33470
rect 35308 33366 35364 33404
rect 34972 33348 35028 33358
rect 35532 33348 35588 33358
rect 35028 33292 35140 33348
rect 34972 33254 35028 33292
rect 35084 32340 35140 33292
rect 35532 33254 35588 33292
rect 35308 32452 35364 32462
rect 35644 32452 35700 34076
rect 36092 33348 36148 35532
rect 36204 35474 36260 35486
rect 36204 35422 36206 35474
rect 36258 35422 36260 35474
rect 36204 34356 36260 35422
rect 36204 34290 36260 34300
rect 36428 35476 36484 35486
rect 36204 34020 36260 34030
rect 36260 33964 36372 34020
rect 36204 33954 36260 33964
rect 36092 33282 36148 33292
rect 35868 33236 35924 33246
rect 35868 33142 35924 33180
rect 35308 32450 35700 32452
rect 35308 32398 35310 32450
rect 35362 32398 35700 32450
rect 35308 32396 35700 32398
rect 35308 32386 35364 32396
rect 35084 32004 35140 32284
rect 35868 32340 35924 32350
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35644 32004 35700 32014
rect 35084 31948 35476 32004
rect 35420 31890 35476 31948
rect 35420 31838 35422 31890
rect 35474 31838 35476 31890
rect 35420 31826 35476 31838
rect 35644 31892 35700 31948
rect 35868 32002 35924 32284
rect 35868 31950 35870 32002
rect 35922 31950 35924 32002
rect 35868 31938 35924 31950
rect 35644 31890 35812 31892
rect 35644 31838 35646 31890
rect 35698 31838 35812 31890
rect 35644 31836 35812 31838
rect 35644 31826 35700 31836
rect 35756 31556 35812 31836
rect 36204 31668 36260 31678
rect 36204 31574 36260 31612
rect 35756 31500 36036 31556
rect 35980 30882 36036 31500
rect 35980 30830 35982 30882
rect 36034 30830 36036 30882
rect 35980 30818 36036 30830
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 34748 29586 34804 29596
rect 35308 29316 35364 29326
rect 35308 29222 35364 29260
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 35308 27300 35364 27310
rect 31164 25106 31220 25116
rect 31500 25284 31556 25294
rect 31164 24946 31220 24958
rect 31164 24894 31166 24946
rect 31218 24894 31220 24946
rect 30828 24612 30884 24622
rect 30828 24518 30884 24556
rect 31164 23828 31220 24894
rect 31388 24722 31444 24734
rect 31388 24670 31390 24722
rect 31442 24670 31444 24722
rect 31388 24612 31444 24670
rect 31500 24724 31556 25228
rect 32172 25172 32228 26852
rect 31500 24658 31556 24668
rect 31836 25116 32228 25172
rect 32396 26850 32452 26862
rect 32396 26798 32398 26850
rect 32450 26798 32452 26850
rect 31836 24834 31892 25116
rect 32396 24836 32452 26798
rect 33964 26852 34132 26908
rect 34972 26964 35028 27002
rect 35196 26964 35252 26974
rect 34972 26962 35252 26964
rect 34972 26910 34974 26962
rect 35026 26910 35198 26962
rect 35250 26910 35252 26962
rect 34972 26908 35252 26910
rect 31836 24782 31838 24834
rect 31890 24782 31892 24834
rect 31388 24546 31444 24556
rect 31836 24388 31892 24782
rect 32172 24780 32452 24836
rect 33404 24836 33460 24846
rect 32060 24724 32116 24734
rect 32060 24630 32116 24668
rect 31836 24322 31892 24332
rect 32172 24052 32228 24780
rect 33404 24742 33460 24780
rect 33068 24722 33124 24734
rect 33068 24670 33070 24722
rect 33122 24670 33124 24722
rect 32396 24612 32452 24622
rect 33068 24612 33124 24670
rect 32396 24610 33124 24612
rect 32396 24558 32398 24610
rect 32450 24558 33124 24610
rect 32396 24556 33124 24558
rect 32396 24546 32452 24556
rect 32172 23986 32228 23996
rect 32620 24388 32676 24398
rect 32620 24050 32676 24332
rect 32620 23998 32622 24050
rect 32674 23998 32676 24050
rect 32620 23986 32676 23998
rect 32956 24052 33012 24062
rect 32956 23958 33012 23996
rect 31164 23762 31220 23772
rect 33180 23940 33236 23950
rect 30604 23492 30884 23548
rect 30828 22932 30884 23492
rect 33180 23380 33236 23884
rect 33628 23380 33684 23390
rect 30716 22876 30884 22932
rect 32732 23378 33684 23380
rect 32732 23326 33182 23378
rect 33234 23326 33630 23378
rect 33682 23326 33684 23378
rect 32732 23324 33684 23326
rect 30492 19460 30548 19470
rect 30380 19234 30436 19246
rect 30380 19182 30382 19234
rect 30434 19182 30436 19234
rect 30380 18340 30436 19182
rect 30492 19234 30548 19404
rect 30716 19346 30772 22876
rect 32732 22484 32788 23324
rect 33180 23314 33236 23324
rect 33628 23314 33684 23324
rect 32508 22482 32788 22484
rect 32508 22430 32734 22482
rect 32786 22430 32788 22482
rect 32508 22428 32788 22430
rect 32508 21588 32564 22428
rect 32732 22418 32788 22428
rect 33740 22930 33796 22942
rect 33740 22878 33742 22930
rect 33794 22878 33796 22930
rect 32508 21494 32564 21532
rect 31724 21476 31780 21486
rect 31500 21474 31780 21476
rect 31500 21422 31726 21474
rect 31778 21422 31780 21474
rect 31500 21420 31780 21422
rect 31500 20690 31556 21420
rect 31724 21410 31780 21420
rect 33628 21476 33684 21486
rect 33740 21476 33796 22878
rect 33628 21474 33796 21476
rect 33628 21422 33630 21474
rect 33682 21422 33796 21474
rect 33628 21420 33796 21422
rect 31836 21364 31892 21374
rect 31836 20802 31892 21308
rect 33068 21364 33124 21374
rect 33068 21270 33124 21308
rect 33404 21362 33460 21374
rect 33404 21310 33406 21362
rect 33458 21310 33460 21362
rect 31836 20750 31838 20802
rect 31890 20750 31892 20802
rect 31836 20738 31892 20750
rect 31500 20638 31502 20690
rect 31554 20638 31556 20690
rect 31500 20626 31556 20638
rect 32732 20580 32788 20590
rect 32732 20486 32788 20524
rect 33404 20580 33460 21310
rect 33404 20514 33460 20524
rect 33292 19906 33348 19918
rect 33292 19854 33294 19906
rect 33346 19854 33348 19906
rect 32844 19460 32900 19470
rect 30716 19294 30718 19346
rect 30770 19294 30772 19346
rect 30716 19282 30772 19294
rect 30828 19348 30884 19358
rect 30492 19182 30494 19234
rect 30546 19182 30548 19234
rect 30492 19170 30548 19182
rect 30828 19234 30884 19292
rect 32396 19348 32452 19358
rect 32396 19254 32452 19292
rect 32844 19346 32900 19404
rect 32844 19294 32846 19346
rect 32898 19294 32900 19346
rect 32844 19282 32900 19294
rect 33292 19348 33348 19854
rect 33628 19908 33684 21420
rect 33628 19842 33684 19852
rect 33740 20020 33796 20030
rect 33740 19906 33796 19964
rect 33740 19854 33742 19906
rect 33794 19854 33796 19906
rect 33292 19282 33348 19292
rect 33628 19460 33684 19470
rect 33740 19460 33796 19854
rect 33684 19404 33796 19460
rect 30828 19182 30830 19234
rect 30882 19182 30884 19234
rect 30828 19170 30884 19182
rect 33628 19234 33684 19404
rect 33964 19346 34020 26852
rect 34972 24722 35028 26908
rect 35196 26898 35252 26908
rect 35308 26178 35364 27244
rect 36204 27188 36260 27198
rect 36204 27094 36260 27132
rect 35308 26126 35310 26178
rect 35362 26126 35364 26178
rect 35308 26114 35364 26126
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35420 25396 35476 25406
rect 35420 25302 35476 25340
rect 35868 25396 35924 25406
rect 35756 25282 35812 25294
rect 35756 25230 35758 25282
rect 35810 25230 35812 25282
rect 34972 24670 34974 24722
rect 35026 24670 35028 24722
rect 34636 24612 34692 24622
rect 34972 24612 35028 24670
rect 34636 24610 35028 24612
rect 34636 24558 34638 24610
rect 34690 24558 35028 24610
rect 34636 24556 35028 24558
rect 35084 24836 35140 24846
rect 34636 23940 34692 24556
rect 35084 24050 35140 24780
rect 35756 24834 35812 25230
rect 35756 24782 35758 24834
rect 35810 24782 35812 24834
rect 35756 24770 35812 24782
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35084 23998 35086 24050
rect 35138 23998 35140 24050
rect 35084 23986 35140 23998
rect 34636 23874 34692 23884
rect 35756 23940 35812 23950
rect 35756 23846 35812 23884
rect 34972 23492 35028 23502
rect 34860 23436 34972 23492
rect 34748 23380 34804 23390
rect 34076 23378 34804 23380
rect 34076 23326 34750 23378
rect 34802 23326 34804 23378
rect 34076 23324 34804 23326
rect 34076 23042 34132 23324
rect 34748 23314 34804 23324
rect 34860 23378 34916 23436
rect 34972 23426 35028 23436
rect 34860 23326 34862 23378
rect 34914 23326 34916 23378
rect 34860 23314 34916 23326
rect 34076 22990 34078 23042
rect 34130 22990 34132 23042
rect 34076 20020 34132 22990
rect 34524 23154 34580 23166
rect 34524 23102 34526 23154
rect 34578 23102 34580 23154
rect 34076 19954 34132 19964
rect 34188 22932 34244 22942
rect 34188 22146 34244 22876
rect 34300 22932 34356 22942
rect 34524 22932 34580 23102
rect 34300 22930 34580 22932
rect 34300 22878 34302 22930
rect 34354 22878 34580 22930
rect 34300 22876 34580 22878
rect 34972 23156 35028 23166
rect 34300 22866 34356 22876
rect 34188 22094 34190 22146
rect 34242 22094 34244 22146
rect 34188 20244 34244 22094
rect 34524 21588 34580 21598
rect 34580 21532 34804 21588
rect 34524 21494 34580 21532
rect 34748 21252 34804 21532
rect 34860 21476 34916 21486
rect 34972 21476 35028 23100
rect 35196 23154 35252 23166
rect 35196 23102 35198 23154
rect 35250 23102 35252 23154
rect 35196 22932 35252 23102
rect 35532 23156 35588 23166
rect 35532 23062 35588 23100
rect 35756 22932 35812 22942
rect 35196 22866 35252 22876
rect 35644 22930 35812 22932
rect 35644 22878 35758 22930
rect 35810 22878 35812 22930
rect 35644 22876 35812 22878
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 35196 22148 35252 22158
rect 35196 22146 35364 22148
rect 35196 22094 35198 22146
rect 35250 22094 35364 22146
rect 35196 22092 35364 22094
rect 35196 22082 35252 22092
rect 34860 21474 35028 21476
rect 34860 21422 34862 21474
rect 34914 21422 35028 21474
rect 34860 21420 35028 21422
rect 34860 21410 34916 21420
rect 35308 21364 35364 22092
rect 35644 21364 35700 22876
rect 35756 22866 35812 22876
rect 35308 21308 35700 21364
rect 34748 21196 35028 21252
rect 34972 20914 35028 21196
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 34972 20862 34974 20914
rect 35026 20862 35028 20914
rect 34972 20850 35028 20862
rect 33964 19294 33966 19346
rect 34018 19294 34020 19346
rect 33964 19282 34020 19294
rect 34076 19348 34132 19358
rect 34188 19348 34244 20188
rect 34860 20580 34916 20590
rect 34636 20132 34692 20142
rect 34636 20038 34692 20076
rect 34132 19292 34244 19348
rect 34412 20018 34468 20030
rect 34412 19966 34414 20018
rect 34466 19966 34468 20018
rect 33628 19182 33630 19234
rect 33682 19182 33684 19234
rect 33628 19170 33684 19182
rect 34076 19234 34132 19292
rect 34076 19182 34078 19234
rect 34130 19182 34132 19234
rect 34076 19170 34132 19182
rect 33404 19124 33460 19134
rect 33292 19122 33460 19124
rect 33292 19070 33406 19122
rect 33458 19070 33460 19122
rect 33292 19068 33460 19070
rect 34412 19124 34468 19966
rect 34524 20020 34580 20030
rect 34524 19926 34580 19964
rect 34748 20020 34804 20030
rect 34748 19926 34804 19964
rect 34860 19796 34916 20524
rect 34972 20244 35028 20254
rect 34972 20018 35028 20188
rect 34972 19966 34974 20018
rect 35026 19966 35028 20018
rect 34972 19954 35028 19966
rect 35532 20020 35588 20030
rect 35308 19908 35364 19918
rect 35308 19814 35364 19852
rect 34748 19740 34916 19796
rect 34636 19124 34692 19134
rect 34412 19122 34692 19124
rect 34412 19070 34638 19122
rect 34690 19070 34692 19122
rect 34412 19068 34692 19070
rect 30716 19012 30772 19022
rect 30716 19010 30996 19012
rect 30716 18958 30718 19010
rect 30770 18958 30996 19010
rect 30716 18956 30996 18958
rect 30716 18946 30772 18956
rect 30492 18340 30548 18350
rect 30380 18284 30492 18340
rect 30492 18246 30548 18284
rect 30828 18340 30884 18350
rect 30828 18246 30884 18284
rect 30492 17780 30548 17790
rect 30492 17666 30548 17724
rect 30492 17614 30494 17666
rect 30546 17614 30548 17666
rect 30492 17602 30548 17614
rect 29260 17054 29262 17106
rect 29314 17054 29316 17106
rect 29260 17042 29316 17054
rect 30156 17052 30268 17108
rect 28588 16046 28590 16098
rect 28642 16046 28644 16098
rect 27356 15486 27358 15538
rect 27410 15486 27412 15538
rect 27356 15474 27412 15486
rect 26348 15092 26628 15148
rect 26684 15314 26740 15326
rect 26684 15262 26686 15314
rect 26738 15262 26740 15314
rect 26684 15148 26740 15262
rect 27132 15314 27188 15326
rect 27132 15262 27134 15314
rect 27186 15262 27188 15314
rect 27132 15148 27188 15262
rect 26684 15092 26852 15148
rect 27132 15092 27412 15148
rect 26460 14980 26516 14990
rect 25788 11506 26068 11508
rect 25788 11454 25902 11506
rect 25954 11454 26068 11506
rect 25788 11452 26068 11454
rect 25900 11442 25956 11452
rect 25340 10836 25396 10846
rect 25340 10742 25396 10780
rect 25452 10836 25508 10846
rect 25452 10834 25956 10836
rect 25452 10782 25454 10834
rect 25506 10782 25956 10834
rect 25452 10780 25956 10782
rect 25452 10770 25508 10780
rect 25676 10612 25732 10622
rect 25676 10518 25732 10556
rect 25788 10610 25844 10622
rect 25788 10558 25790 10610
rect 25842 10558 25844 10610
rect 25340 10500 25396 10510
rect 25228 10498 25396 10500
rect 25228 10446 25342 10498
rect 25394 10446 25396 10498
rect 25228 10444 25396 10446
rect 25340 10434 25396 10444
rect 25452 9042 25508 9054
rect 25788 9044 25844 10558
rect 25900 9940 25956 10780
rect 26012 10612 26068 11452
rect 26236 11442 26292 11452
rect 26348 14754 26404 14766
rect 26348 14702 26350 14754
rect 26402 14702 26404 14754
rect 26348 11506 26404 14702
rect 26460 14642 26516 14924
rect 26460 14590 26462 14642
rect 26514 14590 26516 14642
rect 26460 14578 26516 14590
rect 26796 14530 26852 15092
rect 26796 14478 26798 14530
rect 26850 14478 26852 14530
rect 26796 12066 26852 14478
rect 26796 12014 26798 12066
rect 26850 12014 26852 12066
rect 26796 12002 26852 12014
rect 27020 14980 27076 14990
rect 27020 14530 27076 14924
rect 27356 14754 27412 15092
rect 27356 14702 27358 14754
rect 27410 14702 27412 14754
rect 27356 14690 27412 14702
rect 27020 14478 27022 14530
rect 27074 14478 27076 14530
rect 26348 11454 26350 11506
rect 26402 11454 26404 11506
rect 26012 10546 26068 10556
rect 26348 10836 26404 11454
rect 27020 11508 27076 14478
rect 28588 12180 28644 16046
rect 28700 16772 28756 16782
rect 28700 16100 28756 16716
rect 28812 16770 28868 16782
rect 28812 16718 28814 16770
rect 28866 16718 28868 16770
rect 28812 16658 28868 16718
rect 28812 16606 28814 16658
rect 28866 16606 28868 16658
rect 28812 16594 28868 16606
rect 29372 16660 29428 16670
rect 29372 16658 29540 16660
rect 29372 16606 29374 16658
rect 29426 16606 29540 16658
rect 29372 16604 29540 16606
rect 29372 16594 29428 16604
rect 28700 15538 28756 16044
rect 29484 16322 29540 16604
rect 29484 16270 29486 16322
rect 29538 16270 29540 16322
rect 28700 15486 28702 15538
rect 28754 15486 28756 15538
rect 28700 15474 28756 15486
rect 29148 15874 29204 15886
rect 29148 15822 29150 15874
rect 29202 15822 29204 15874
rect 29036 15314 29092 15326
rect 29036 15262 29038 15314
rect 29090 15262 29092 15314
rect 29036 13636 29092 15262
rect 29148 15148 29204 15822
rect 29148 15092 29316 15148
rect 29260 14530 29316 15092
rect 29484 14980 29540 16270
rect 29708 16100 29764 16110
rect 29708 16006 29764 16044
rect 29484 14914 29540 14924
rect 29708 15202 29764 15214
rect 29708 15150 29710 15202
rect 29762 15150 29764 15202
rect 29260 14478 29262 14530
rect 29314 14478 29316 14530
rect 29260 14466 29316 14478
rect 29596 14420 29652 14430
rect 29708 14420 29764 15150
rect 29596 14418 29764 14420
rect 29596 14366 29598 14418
rect 29650 14366 29764 14418
rect 29596 14364 29764 14366
rect 29596 14354 29652 14364
rect 29036 13570 29092 13580
rect 30044 13636 30100 13646
rect 28588 12114 28644 12124
rect 29708 12180 29764 12190
rect 28028 12068 28084 12078
rect 27132 11508 27188 11518
rect 27020 11506 27860 11508
rect 27020 11454 27134 11506
rect 27186 11454 27860 11506
rect 27020 11452 27860 11454
rect 27132 11442 27188 11452
rect 26348 10612 26404 10780
rect 26796 11284 26852 11294
rect 27692 11284 27748 11294
rect 26796 10834 26852 11228
rect 26796 10782 26798 10834
rect 26850 10782 26852 10834
rect 26796 10770 26852 10782
rect 27468 11282 27748 11284
rect 27468 11230 27694 11282
rect 27746 11230 27748 11282
rect 27468 11228 27748 11230
rect 27468 10834 27524 11228
rect 27692 11218 27748 11228
rect 27468 10782 27470 10834
rect 27522 10782 27524 10834
rect 27468 10770 27524 10782
rect 26460 10612 26516 10622
rect 26348 10610 26516 10612
rect 26348 10558 26462 10610
rect 26514 10558 26516 10610
rect 26348 10556 26516 10558
rect 26348 10052 26404 10556
rect 26460 10546 26516 10556
rect 26684 10610 26740 10622
rect 26908 10612 26964 10622
rect 26684 10558 26686 10610
rect 26738 10558 26740 10610
rect 26012 9940 26068 9950
rect 25900 9938 26068 9940
rect 25900 9886 26014 9938
rect 26066 9886 26068 9938
rect 25900 9884 26068 9886
rect 26012 9604 26068 9884
rect 26348 9826 26404 9996
rect 26460 9940 26516 9950
rect 26460 9846 26516 9884
rect 26684 9940 26740 10558
rect 26684 9874 26740 9884
rect 26796 10556 26908 10612
rect 26348 9774 26350 9826
rect 26402 9774 26404 9826
rect 26348 9762 26404 9774
rect 26796 9826 26852 10556
rect 26908 10518 26964 10556
rect 27132 10612 27188 10622
rect 27468 10612 27524 10622
rect 27132 10610 27300 10612
rect 27132 10558 27134 10610
rect 27186 10558 27300 10610
rect 27132 10556 27300 10558
rect 27132 10546 27188 10556
rect 27244 10050 27300 10556
rect 27244 9998 27246 10050
rect 27298 9998 27300 10050
rect 27244 9986 27300 9998
rect 27468 9938 27524 10556
rect 27468 9886 27470 9938
rect 27522 9886 27524 9938
rect 27468 9874 27524 9886
rect 27804 10386 27860 11452
rect 28028 11282 28084 12012
rect 28924 12068 28980 12078
rect 28924 11974 28980 12012
rect 29708 11956 29764 12124
rect 29932 11956 29988 11966
rect 29708 11954 29988 11956
rect 29708 11902 29934 11954
rect 29986 11902 29988 11954
rect 29708 11900 29988 11902
rect 28028 11230 28030 11282
rect 28082 11230 28084 11282
rect 28028 11218 28084 11230
rect 29932 11170 29988 11900
rect 29932 11118 29934 11170
rect 29986 11118 29988 11170
rect 27804 10334 27806 10386
rect 27858 10334 27860 10386
rect 26796 9774 26798 9826
rect 26850 9774 26852 9826
rect 26796 9762 26852 9774
rect 27020 9714 27076 9726
rect 27020 9662 27022 9714
rect 27074 9662 27076 9714
rect 26012 9548 26292 9604
rect 25452 8990 25454 9042
rect 25506 8990 25508 9042
rect 25452 8484 25508 8990
rect 25452 8418 25508 8428
rect 25676 8988 25844 9044
rect 25564 8260 25620 8270
rect 25564 8166 25620 8204
rect 25116 8036 25172 8046
rect 24444 5854 24446 5906
rect 24498 5854 24500 5906
rect 24444 5842 24500 5854
rect 24892 6466 24948 6478
rect 24892 6414 24894 6466
rect 24946 6414 24948 6466
rect 24892 5908 24948 6414
rect 24892 5842 24948 5852
rect 23212 5742 23214 5794
rect 23266 5742 23268 5794
rect 23212 5730 23268 5742
rect 23884 5684 23940 5694
rect 23548 5682 23940 5684
rect 23548 5630 23886 5682
rect 23938 5630 23940 5682
rect 23548 5628 23940 5630
rect 22316 5282 22372 5292
rect 23100 5460 23156 5470
rect 21308 5182 21310 5234
rect 21362 5182 21364 5234
rect 21308 5170 21364 5182
rect 23100 5234 23156 5404
rect 23100 5182 23102 5234
rect 23154 5182 23156 5234
rect 23100 5170 23156 5182
rect 23324 5236 23380 5246
rect 21868 5124 21924 5134
rect 22428 5124 22484 5134
rect 21868 5122 22484 5124
rect 21868 5070 21870 5122
rect 21922 5070 22430 5122
rect 22482 5070 22484 5122
rect 21868 5068 22484 5070
rect 21868 5058 21924 5068
rect 22428 5058 22484 5068
rect 20076 4900 20132 4938
rect 22204 4900 22260 4910
rect 20076 4834 20132 4844
rect 22092 4898 22260 4900
rect 22092 4846 22206 4898
rect 22258 4846 22260 4898
rect 22092 4844 22260 4846
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 19628 4510 19630 4562
rect 19682 4510 19684 4562
rect 19628 4498 19684 4510
rect 22092 4450 22148 4844
rect 22204 4834 22260 4844
rect 23324 4564 23380 5180
rect 23548 5122 23604 5628
rect 23884 5618 23940 5628
rect 25116 5460 25172 7980
rect 25564 6692 25620 6702
rect 25564 5908 25620 6636
rect 25676 5908 25732 8988
rect 26124 8932 26180 8942
rect 25788 8930 26180 8932
rect 25788 8878 26126 8930
rect 26178 8878 26180 8930
rect 25788 8876 26180 8878
rect 25788 8146 25844 8876
rect 26124 8866 26180 8876
rect 26124 8372 26180 8382
rect 26236 8372 26292 9548
rect 26124 8370 26292 8372
rect 26124 8318 26126 8370
rect 26178 8318 26292 8370
rect 26124 8316 26292 8318
rect 26572 9602 26628 9614
rect 26572 9550 26574 9602
rect 26626 9550 26628 9602
rect 26124 8306 26180 8316
rect 25788 8094 25790 8146
rect 25842 8094 25844 8146
rect 25788 8082 25844 8094
rect 26348 8258 26404 8270
rect 26348 8206 26350 8258
rect 26402 8206 26404 8258
rect 26348 8036 26404 8206
rect 26348 7970 26404 7980
rect 26572 7364 26628 9550
rect 27020 8484 27076 9662
rect 27020 8428 27636 8484
rect 27020 8260 27076 8270
rect 27020 8166 27076 8204
rect 26684 8034 26740 8046
rect 26684 7982 26686 8034
rect 26738 7982 26740 8034
rect 26684 7474 26740 7982
rect 27132 7812 27188 8428
rect 27580 8370 27636 8428
rect 27580 8318 27582 8370
rect 27634 8318 27636 8370
rect 27580 8306 27636 8318
rect 27020 7756 27188 7812
rect 27244 8260 27300 8270
rect 26908 7588 26964 7598
rect 26908 7494 26964 7532
rect 26684 7422 26686 7474
rect 26738 7422 26740 7474
rect 26684 7410 26740 7422
rect 26572 7298 26628 7308
rect 25788 5908 25844 5918
rect 25676 5906 26068 5908
rect 25676 5854 25790 5906
rect 25842 5854 26068 5906
rect 25676 5852 26068 5854
rect 25564 5814 25620 5852
rect 25788 5842 25844 5852
rect 25116 5394 25172 5404
rect 25228 5682 25284 5694
rect 25228 5630 25230 5682
rect 25282 5630 25284 5682
rect 23548 5070 23550 5122
rect 23602 5070 23604 5122
rect 23548 5058 23604 5070
rect 24220 5236 24276 5246
rect 24220 5122 24276 5180
rect 24220 5070 24222 5122
rect 24274 5070 24276 5122
rect 24220 5058 24276 5070
rect 24444 5124 24500 5134
rect 22092 4398 22094 4450
rect 22146 4398 22148 4450
rect 22092 4386 22148 4398
rect 23212 4562 23380 4564
rect 23212 4510 23326 4562
rect 23378 4510 23380 4562
rect 23212 4508 23380 4510
rect 19404 4286 19406 4338
rect 19458 4286 19460 4338
rect 19404 4274 19460 4286
rect 22876 4340 22932 4350
rect 23212 4340 23268 4508
rect 23324 4498 23380 4508
rect 23772 4898 23828 4910
rect 23772 4846 23774 4898
rect 23826 4846 23828 4898
rect 22876 4338 23268 4340
rect 22876 4286 22878 4338
rect 22930 4286 23268 4338
rect 22876 4284 23268 4286
rect 22876 4274 22932 4284
rect 19964 4228 20020 4238
rect 19516 4226 20020 4228
rect 19516 4174 19966 4226
rect 20018 4174 20020 4226
rect 19516 4172 20020 4174
rect 19516 4116 19572 4172
rect 19964 4162 20020 4172
rect 19292 4060 19572 4116
rect 17724 3836 18116 3892
rect 16044 3556 16100 3566
rect 15484 3502 15486 3554
rect 15538 3502 15540 3554
rect 15036 3444 15092 3454
rect 14476 2482 14532 2492
rect 14588 3332 14868 3388
rect 14924 3442 15092 3444
rect 14924 3390 15038 3442
rect 15090 3390 15092 3442
rect 14924 3388 15092 3390
rect 13692 1596 13860 1652
rect 12348 1484 12852 1540
rect 12796 400 12852 1484
rect 13692 400 13748 1596
rect 14588 400 14644 3332
rect 14812 2772 14868 2782
rect 14924 2772 14980 3388
rect 15036 3378 15092 3388
rect 14812 2770 14980 2772
rect 14812 2718 14814 2770
rect 14866 2718 14980 2770
rect 14812 2716 14980 2718
rect 15148 3332 15204 3342
rect 14812 2706 14868 2716
rect 14924 1876 14980 1886
rect 15148 1876 15204 3276
rect 15260 2884 15316 2894
rect 15260 2790 15316 2828
rect 14924 1874 15204 1876
rect 14924 1822 14926 1874
rect 14978 1822 15204 1874
rect 14924 1820 15204 1822
rect 14924 1810 14980 1820
rect 15484 400 15540 3502
rect 15708 3554 16100 3556
rect 15708 3502 16046 3554
rect 16098 3502 16100 3554
rect 15708 3500 16100 3502
rect 15708 3442 15764 3500
rect 16044 3490 16100 3500
rect 15708 3390 15710 3442
rect 15762 3390 15764 3442
rect 15708 3378 15764 3390
rect 17164 3442 17220 3454
rect 17164 3390 17166 3442
rect 17218 3390 17220 3442
rect 16156 3332 16212 3342
rect 16156 3238 16212 3276
rect 16380 2996 16436 3006
rect 16268 2940 16380 2996
rect 17164 2996 17220 3390
rect 17388 2996 17444 3006
rect 17164 2994 17444 2996
rect 17164 2942 17390 2994
rect 17442 2942 17444 2994
rect 17164 2940 17444 2942
rect 16268 1986 16324 2940
rect 16380 2930 16436 2940
rect 17388 2930 17444 2940
rect 16268 1934 16270 1986
rect 16322 1934 16324 1986
rect 16268 1922 16324 1934
rect 16380 2772 16436 2782
rect 16380 400 16436 2716
rect 17612 2772 17668 2782
rect 17612 2678 17668 2716
rect 17612 1988 17668 1998
rect 17724 1988 17780 3836
rect 18172 3556 18228 3566
rect 18172 3554 18564 3556
rect 18172 3502 18174 3554
rect 18226 3502 18564 3554
rect 18172 3500 18564 3502
rect 18172 3490 18228 3500
rect 17388 1986 17780 1988
rect 17388 1934 17614 1986
rect 17666 1934 17780 1986
rect 17388 1932 17780 1934
rect 17836 3444 17892 3454
rect 17276 1764 17332 1774
rect 17276 1670 17332 1708
rect 17388 1540 17444 1932
rect 17612 1922 17668 1932
rect 17836 1874 17892 3388
rect 18172 2772 18228 2782
rect 18172 2678 18228 2716
rect 18508 2660 18564 3500
rect 23212 3554 23268 4284
rect 23772 3668 23828 4846
rect 24444 4338 24500 5068
rect 25228 5124 25284 5630
rect 25228 5058 25284 5068
rect 24892 5012 24948 5022
rect 24668 5010 24948 5012
rect 24668 4958 24894 5010
rect 24946 4958 24948 5010
rect 24668 4956 24948 4958
rect 24668 4562 24724 4956
rect 24892 4946 24948 4956
rect 24668 4510 24670 4562
rect 24722 4510 24724 4562
rect 24668 4498 24724 4510
rect 25228 4452 25284 4462
rect 25228 4358 25284 4396
rect 25564 4450 25620 4462
rect 25564 4398 25566 4450
rect 25618 4398 25620 4450
rect 24444 4286 24446 4338
rect 24498 4286 24500 4338
rect 24444 4274 24500 4286
rect 23884 3668 23940 3678
rect 23772 3666 23940 3668
rect 23772 3614 23886 3666
rect 23938 3614 23940 3666
rect 23772 3612 23940 3614
rect 23884 3602 23940 3612
rect 23212 3502 23214 3554
rect 23266 3502 23268 3554
rect 23212 3490 23268 3502
rect 18620 3444 18676 3482
rect 18620 3378 18676 3388
rect 20860 3332 20916 3342
rect 22652 3332 22708 3342
rect 25564 3332 25620 4398
rect 20860 3330 21140 3332
rect 20860 3278 20862 3330
rect 20914 3278 21140 3330
rect 20860 3276 21140 3278
rect 20860 3266 20916 3276
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 19852 2996 19908 3006
rect 19852 2902 19908 2940
rect 20300 2884 20356 2894
rect 20188 2882 20356 2884
rect 20188 2830 20302 2882
rect 20354 2830 20356 2882
rect 20188 2828 20356 2830
rect 19740 2770 19796 2782
rect 19740 2718 19742 2770
rect 19794 2718 19796 2770
rect 18508 2604 18788 2660
rect 18396 1876 18452 1886
rect 17836 1822 17838 1874
rect 17890 1822 17892 1874
rect 17836 1810 17892 1822
rect 18172 1874 18452 1876
rect 18172 1822 18398 1874
rect 18450 1822 18452 1874
rect 18172 1820 18452 1822
rect 17276 1484 17444 1540
rect 18172 1764 18228 1820
rect 18396 1810 18452 1820
rect 18732 1874 18788 2604
rect 18732 1822 18734 1874
rect 18786 1822 18788 1874
rect 18732 1810 18788 1822
rect 19068 2658 19124 2670
rect 19516 2660 19572 2670
rect 19068 2606 19070 2658
rect 19122 2606 19124 2658
rect 19068 1876 19124 2606
rect 19404 2658 19572 2660
rect 19404 2606 19518 2658
rect 19570 2606 19572 2658
rect 19404 2604 19572 2606
rect 19180 1876 19236 1886
rect 19068 1874 19236 1876
rect 19068 1822 19182 1874
rect 19234 1822 19236 1874
rect 19068 1820 19236 1822
rect 17276 400 17332 1484
rect 18172 400 18228 1708
rect 19068 400 19124 1820
rect 19180 1810 19236 1820
rect 19404 1652 19460 2604
rect 19516 2594 19572 2604
rect 19516 1876 19572 1886
rect 19740 1876 19796 2718
rect 19516 1874 19796 1876
rect 19516 1822 19518 1874
rect 19570 1822 19796 1874
rect 19516 1820 19796 1822
rect 19852 1874 19908 1886
rect 19852 1822 19854 1874
rect 19906 1822 19908 1874
rect 19516 1810 19572 1820
rect 19852 1764 19908 1822
rect 20188 1874 20244 2828
rect 20300 2818 20356 2828
rect 21084 1988 21140 3276
rect 22652 3330 22932 3332
rect 22652 3278 22654 3330
rect 22706 3278 22932 3330
rect 22652 3276 22932 3278
rect 22652 3266 22708 3276
rect 20188 1822 20190 1874
rect 20242 1822 20244 1874
rect 20188 1810 20244 1822
rect 20860 1986 21140 1988
rect 20860 1934 21086 1986
rect 21138 1934 21140 1986
rect 20860 1932 21140 1934
rect 19628 1708 19908 1764
rect 19628 1652 19684 1708
rect 19404 1596 19684 1652
rect 19628 1428 19684 1596
rect 19836 1596 20100 1606
rect 19892 1540 19940 1596
rect 19996 1540 20044 1596
rect 19836 1530 20100 1540
rect 19628 1372 20020 1428
rect 19964 400 20020 1372
rect 20860 400 20916 1932
rect 21084 1922 21140 1932
rect 21420 2884 21476 2894
rect 21420 1874 21476 2828
rect 22316 2884 22372 2894
rect 22316 2790 22372 2828
rect 21868 2772 21924 2782
rect 21868 2770 22260 2772
rect 21868 2718 21870 2770
rect 21922 2718 22260 2770
rect 21868 2716 22260 2718
rect 21868 2706 21924 2716
rect 21980 1988 22036 1998
rect 21420 1822 21422 1874
rect 21474 1822 21476 1874
rect 21420 1810 21476 1822
rect 21756 1932 21980 1988
rect 21756 400 21812 1932
rect 21980 1894 22036 1932
rect 22204 1876 22260 2716
rect 22876 1988 22932 3276
rect 25564 3266 25620 3276
rect 25900 4338 25956 4350
rect 25900 4286 25902 4338
rect 25954 4286 25956 4338
rect 25900 2994 25956 4286
rect 26012 3666 26068 5852
rect 26572 5236 26628 5246
rect 26012 3614 26014 3666
rect 26066 3614 26068 3666
rect 26012 3602 26068 3614
rect 26460 4226 26516 4238
rect 26460 4174 26462 4226
rect 26514 4174 26516 4226
rect 26460 3108 26516 4174
rect 26572 3666 26628 5180
rect 27020 5234 27076 7756
rect 27244 7474 27300 8204
rect 27244 7422 27246 7474
rect 27298 7422 27300 7474
rect 27244 5460 27300 7422
rect 27356 8258 27412 8270
rect 27356 8206 27358 8258
rect 27410 8206 27412 8258
rect 27356 8036 27412 8206
rect 27804 8036 27860 10334
rect 28028 10498 28084 10510
rect 28028 10446 28030 10498
rect 28082 10446 28084 10498
rect 27916 10052 27972 10062
rect 27916 9938 27972 9996
rect 27916 9886 27918 9938
rect 27970 9886 27972 9938
rect 27916 9874 27972 9886
rect 28028 10050 28084 10446
rect 28028 9998 28030 10050
rect 28082 9998 28084 10050
rect 28028 8932 28084 9998
rect 29148 9940 29204 9950
rect 28364 9602 28420 9614
rect 28364 9550 28366 9602
rect 28418 9550 28420 9602
rect 28252 8932 28308 8942
rect 28028 8930 28308 8932
rect 28028 8878 28254 8930
rect 28306 8878 28308 8930
rect 28028 8876 28308 8878
rect 28364 8932 28420 9550
rect 28700 8932 28756 8942
rect 28364 8930 28756 8932
rect 28364 8878 28702 8930
rect 28754 8878 28756 8930
rect 28364 8876 28756 8878
rect 28252 8866 28308 8876
rect 28700 8484 28756 8876
rect 29148 8930 29204 9884
rect 29708 9826 29764 9838
rect 29708 9774 29710 9826
rect 29762 9774 29764 9826
rect 29708 9716 29764 9774
rect 29708 9650 29764 9660
rect 29148 8878 29150 8930
rect 29202 8878 29204 8930
rect 29148 8866 29204 8878
rect 28700 8418 28756 8428
rect 29932 8484 29988 11118
rect 29932 8390 29988 8428
rect 30044 9938 30100 13580
rect 30156 13188 30212 17052
rect 30268 17042 30324 17052
rect 30716 16212 30772 16222
rect 30604 14980 30660 14990
rect 30604 14644 30660 14924
rect 30604 14550 30660 14588
rect 30156 13122 30212 13132
rect 30268 13076 30324 13086
rect 30716 13076 30772 16156
rect 30940 15316 30996 18956
rect 31388 19010 31444 19022
rect 31388 18958 31390 19010
rect 31442 18958 31444 19010
rect 31052 18788 31108 18798
rect 31388 18788 31444 18958
rect 31108 18732 31444 18788
rect 31052 18450 31108 18732
rect 31052 18398 31054 18450
rect 31106 18398 31108 18450
rect 31052 16212 31108 18398
rect 31724 18562 31780 18574
rect 31724 18510 31726 18562
rect 31778 18510 31780 18562
rect 31388 18340 31444 18350
rect 31388 18246 31444 18284
rect 31724 18004 31780 18510
rect 32060 18450 32116 18462
rect 32060 18398 32062 18450
rect 32114 18398 32116 18450
rect 32060 18340 32116 18398
rect 32060 18274 32116 18284
rect 32508 18338 32564 18350
rect 32508 18286 32510 18338
rect 32562 18286 32564 18338
rect 31164 17948 31780 18004
rect 31164 17778 31220 17948
rect 31164 17726 31166 17778
rect 31218 17726 31220 17778
rect 31164 17714 31220 17726
rect 32508 17780 32564 18286
rect 32508 17714 32564 17724
rect 33292 17780 33348 19068
rect 33404 19058 33460 19068
rect 33852 19010 33908 19022
rect 33852 18958 33854 19010
rect 33906 18958 33908 19010
rect 33740 18562 33796 18574
rect 33740 18510 33742 18562
rect 33794 18510 33796 18562
rect 33516 18450 33572 18462
rect 33516 18398 33518 18450
rect 33570 18398 33572 18450
rect 33516 17892 33572 18398
rect 33628 17892 33684 17902
rect 33516 17890 33684 17892
rect 33516 17838 33630 17890
rect 33682 17838 33684 17890
rect 33516 17836 33684 17838
rect 33628 17826 33684 17836
rect 33292 17686 33348 17724
rect 33180 17668 33236 17678
rect 32508 17108 32564 17118
rect 31052 16146 31108 16156
rect 32284 17052 32508 17108
rect 32284 15538 32340 17052
rect 32508 17014 32564 17052
rect 33180 17108 33236 17612
rect 33180 16882 33236 17052
rect 33740 16996 33796 18510
rect 33852 17220 33908 18958
rect 34300 18788 34356 18798
rect 34300 18674 34356 18732
rect 34300 18622 34302 18674
rect 34354 18622 34356 18674
rect 34300 18610 34356 18622
rect 34636 18452 34692 19068
rect 34636 18386 34692 18396
rect 34188 17780 34244 17790
rect 34188 17686 34244 17724
rect 33964 17666 34020 17678
rect 33964 17614 33966 17666
rect 34018 17614 34020 17666
rect 33964 17556 34020 17614
rect 34636 17556 34692 17566
rect 34748 17556 34804 19740
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 34860 19460 34916 19470
rect 34860 19234 34916 19404
rect 35532 19348 35588 19964
rect 34860 19182 34862 19234
rect 34914 19182 34916 19234
rect 34860 18788 34916 19182
rect 35308 19346 35588 19348
rect 35308 19294 35534 19346
rect 35586 19294 35588 19346
rect 35308 19292 35588 19294
rect 35196 19012 35252 19022
rect 35196 18918 35252 18956
rect 34860 18722 34916 18732
rect 34972 18564 35028 18574
rect 34972 18338 35028 18508
rect 34972 18286 34974 18338
rect 35026 18286 35028 18338
rect 34972 17892 35028 18286
rect 35308 18338 35364 19292
rect 35532 19282 35588 19292
rect 35644 19236 35700 21308
rect 35868 21028 35924 25340
rect 36092 25394 36148 25406
rect 36092 25342 36094 25394
rect 36146 25342 36148 25394
rect 36092 23378 36148 25342
rect 36092 23326 36094 23378
rect 36146 23326 36148 23378
rect 36092 23314 36148 23326
rect 35756 20972 35924 21028
rect 36092 21476 36148 21486
rect 35756 19460 35812 20972
rect 35868 20804 35924 20814
rect 35868 20802 36036 20804
rect 35868 20750 35870 20802
rect 35922 20750 36036 20802
rect 35868 20748 36036 20750
rect 35868 20738 35924 20748
rect 35980 19460 36036 20748
rect 36092 20690 36148 21420
rect 36092 20638 36094 20690
rect 36146 20638 36148 20690
rect 36092 20626 36148 20638
rect 36316 20132 36372 33964
rect 36428 33348 36484 35420
rect 36428 33282 36484 33292
rect 36428 30884 36484 30894
rect 36428 30790 36484 30828
rect 36540 23492 36596 38612
rect 36652 26908 36708 41132
rect 36764 35588 36820 45500
rect 36764 35494 36820 35532
rect 36876 42980 36932 42990
rect 36876 34244 36932 42924
rect 36988 42644 37044 42654
rect 36988 42550 37044 42588
rect 37324 42530 37380 42542
rect 37324 42478 37326 42530
rect 37378 42478 37380 42530
rect 37324 42084 37380 42478
rect 37436 42084 37492 42094
rect 37324 42082 37492 42084
rect 37324 42030 37438 42082
rect 37490 42030 37492 42082
rect 37324 42028 37492 42030
rect 37436 42018 37492 42028
rect 37436 41412 37492 41422
rect 37436 41318 37492 41356
rect 37100 41300 37156 41310
rect 37100 41206 37156 41244
rect 37772 40290 37828 40302
rect 37772 40238 37774 40290
rect 37826 40238 37828 40290
rect 37212 39620 37268 39630
rect 37772 39620 37828 40238
rect 37212 39618 37828 39620
rect 37212 39566 37214 39618
rect 37266 39566 37828 39618
rect 37212 39564 37828 39566
rect 37884 39730 37940 50316
rect 38220 48802 38276 48814
rect 38220 48750 38222 48802
rect 38274 48750 38276 48802
rect 38108 48244 38164 48254
rect 38220 48244 38276 48750
rect 38108 48242 38276 48244
rect 38108 48190 38110 48242
rect 38162 48190 38276 48242
rect 38108 48188 38276 48190
rect 37996 47234 38052 47246
rect 37996 47182 37998 47234
rect 38050 47182 38052 47234
rect 37996 47012 38052 47182
rect 37996 46946 38052 46956
rect 38108 46674 38164 48188
rect 38108 46622 38110 46674
rect 38162 46622 38164 46674
rect 38108 45668 38164 46622
rect 38220 45668 38276 45678
rect 38164 45666 38276 45668
rect 38164 45614 38222 45666
rect 38274 45614 38276 45666
rect 38164 45612 38276 45614
rect 38108 45602 38164 45612
rect 38220 45602 38276 45612
rect 38220 42868 38276 42878
rect 38220 41972 38276 42812
rect 37884 39678 37886 39730
rect 37938 39678 37940 39730
rect 36988 37940 37044 37950
rect 36988 37846 37044 37884
rect 37212 37716 37268 39564
rect 37436 38722 37492 38734
rect 37436 38670 37438 38722
rect 37490 38670 37492 38722
rect 37324 37940 37380 37950
rect 37436 37940 37492 38670
rect 37884 38668 37940 39678
rect 37772 38612 37940 38668
rect 38108 41970 38276 41972
rect 38108 41918 38222 41970
rect 38274 41918 38276 41970
rect 38108 41916 38276 41918
rect 38108 38834 38164 41916
rect 38220 41906 38276 41916
rect 38220 41748 38276 41758
rect 38220 41188 38276 41692
rect 38220 41186 38388 41188
rect 38220 41134 38222 41186
rect 38274 41134 38388 41186
rect 38220 41132 38388 41134
rect 38220 41122 38276 41132
rect 38332 40626 38388 41132
rect 38332 40574 38334 40626
rect 38386 40574 38388 40626
rect 38332 40562 38388 40574
rect 38108 38782 38110 38834
rect 38162 38782 38164 38834
rect 38108 38668 38164 38782
rect 38108 38612 38276 38668
rect 37772 38052 37828 38612
rect 37772 37958 37828 37996
rect 38220 38162 38276 38612
rect 38220 38110 38222 38162
rect 38274 38110 38276 38162
rect 37324 37938 37492 37940
rect 37324 37886 37326 37938
rect 37378 37886 37492 37938
rect 37324 37884 37492 37886
rect 37548 37940 37604 37950
rect 37324 37874 37380 37884
rect 37212 37660 37380 37716
rect 36988 36482 37044 36494
rect 36988 36430 36990 36482
rect 37042 36430 37044 36482
rect 36988 35812 37044 36430
rect 36988 35746 37044 35756
rect 37212 36482 37268 36494
rect 37212 36430 37214 36482
rect 37266 36430 37268 36482
rect 36988 35586 37044 35598
rect 36988 35534 36990 35586
rect 37042 35534 37044 35586
rect 36988 35364 37044 35534
rect 37212 35588 37268 36430
rect 37212 35522 37268 35532
rect 36988 35298 37044 35308
rect 36876 34178 36932 34188
rect 36876 33348 36932 33358
rect 37324 33348 37380 37660
rect 37436 37156 37492 37166
rect 37436 37062 37492 37100
rect 37548 36706 37604 37884
rect 37548 36654 37550 36706
rect 37602 36654 37604 36706
rect 37548 36642 37604 36654
rect 38220 37266 38276 38110
rect 38220 37214 38222 37266
rect 38274 37214 38276 37266
rect 38220 36594 38276 37214
rect 38220 36542 38222 36594
rect 38274 36542 38276 36594
rect 38220 36530 38276 36542
rect 36876 28082 36932 33292
rect 37212 33292 37380 33348
rect 38220 34356 38276 34366
rect 36988 33236 37044 33246
rect 36988 33142 37044 33180
rect 36988 31668 37044 31678
rect 36988 31574 37044 31612
rect 36876 28030 36878 28082
rect 36930 28030 36932 28082
rect 36876 28018 36932 28030
rect 36988 27858 37044 27870
rect 36988 27806 36990 27858
rect 37042 27806 37044 27858
rect 36988 27300 37044 27806
rect 36988 27234 37044 27244
rect 36988 26962 37044 26974
rect 36988 26910 36990 26962
rect 37042 26910 37044 26962
rect 36652 26852 36820 26908
rect 36764 25396 36820 26852
rect 36988 25730 37044 26910
rect 36988 25678 36990 25730
rect 37042 25678 37044 25730
rect 36988 25666 37044 25678
rect 36764 25330 36820 25340
rect 36540 23426 36596 23436
rect 36988 21476 37044 21486
rect 36988 21382 37044 21420
rect 36316 20066 36372 20076
rect 36092 19460 36148 19470
rect 35980 19458 36148 19460
rect 35980 19406 36094 19458
rect 36146 19406 36148 19458
rect 35980 19404 36148 19406
rect 35756 19394 35812 19404
rect 36092 19394 36148 19404
rect 35756 19236 35812 19246
rect 35644 19234 35812 19236
rect 35644 19182 35758 19234
rect 35810 19182 35812 19234
rect 35644 19180 35812 19182
rect 35756 18564 35812 19180
rect 36988 19122 37044 19134
rect 36988 19070 36990 19122
rect 37042 19070 37044 19122
rect 36988 19012 37044 19070
rect 36988 18946 37044 18956
rect 35756 18498 35812 18508
rect 35308 18286 35310 18338
rect 35362 18286 35364 18338
rect 35308 18274 35364 18286
rect 35980 18452 36036 18462
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 34972 17836 35252 17892
rect 35084 17668 35140 17678
rect 35084 17574 35140 17612
rect 33964 17554 34804 17556
rect 33964 17502 34638 17554
rect 34690 17502 34804 17554
rect 33964 17500 34804 17502
rect 34636 17490 34692 17500
rect 35196 17220 35252 17836
rect 33852 17164 35028 17220
rect 33852 16996 33908 17006
rect 33740 16994 33908 16996
rect 33740 16942 33854 16994
rect 33906 16942 33908 16994
rect 33740 16940 33908 16942
rect 33852 16930 33908 16940
rect 33180 16830 33182 16882
rect 33234 16830 33236 16882
rect 33180 16818 33236 16830
rect 34972 16210 35028 17164
rect 34972 16158 34974 16210
rect 35026 16158 35028 16210
rect 32284 15486 32286 15538
rect 32338 15486 32340 15538
rect 30940 14642 30996 15260
rect 31836 15316 31892 15326
rect 31836 15202 31892 15260
rect 31836 15150 31838 15202
rect 31890 15150 31892 15202
rect 31836 15138 31892 15150
rect 30940 14590 30942 14642
rect 30994 14590 30996 14642
rect 30940 14578 30996 14590
rect 31164 14644 31220 14654
rect 31164 14550 31220 14588
rect 31948 14532 32004 14542
rect 32284 14532 32340 15486
rect 34636 16100 34692 16110
rect 34636 15874 34692 16044
rect 34636 15822 34638 15874
rect 34690 15822 34692 15874
rect 34636 15204 34692 15822
rect 34972 15148 35028 16158
rect 35084 17164 35252 17220
rect 35084 16100 35140 17164
rect 35980 16770 36036 18396
rect 36652 18340 36708 18350
rect 36652 17106 36708 18284
rect 36652 17054 36654 17106
rect 36706 17054 36708 17106
rect 36652 17042 36708 17054
rect 36316 16884 36372 16894
rect 35980 16718 35982 16770
rect 36034 16718 36036 16770
rect 35980 16706 36036 16718
rect 36092 16882 36372 16884
rect 36092 16830 36318 16882
rect 36370 16830 36372 16882
rect 36092 16828 36372 16830
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 36092 16436 36148 16828
rect 36316 16818 36372 16828
rect 35196 16426 35460 16436
rect 35532 16380 36148 16436
rect 35532 16322 35588 16380
rect 35532 16270 35534 16322
rect 35586 16270 35588 16322
rect 35532 16258 35588 16270
rect 35196 16100 35252 16110
rect 35084 16044 35196 16100
rect 35196 16006 35252 16044
rect 34636 15138 34692 15148
rect 34748 15092 35028 15148
rect 34748 14642 34804 15092
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 34748 14590 34750 14642
rect 34802 14590 34804 14642
rect 34748 14578 34804 14590
rect 31948 14530 32340 14532
rect 31948 14478 31950 14530
rect 32002 14478 32340 14530
rect 31948 14476 32340 14478
rect 31500 14308 31556 14318
rect 31500 14214 31556 14252
rect 31500 13636 31556 13646
rect 31500 13542 31556 13580
rect 31948 13636 32004 14476
rect 32620 14420 32676 14430
rect 32620 14418 33124 14420
rect 32620 14366 32622 14418
rect 32674 14366 33124 14418
rect 32620 14364 33124 14366
rect 32620 14354 32676 14364
rect 33068 13970 33124 14364
rect 33068 13918 33070 13970
rect 33122 13918 33124 13970
rect 33068 13906 33124 13918
rect 33292 14308 33348 14318
rect 33292 13746 33348 14252
rect 33292 13694 33294 13746
rect 33346 13694 33348 13746
rect 33292 13682 33348 13694
rect 31948 13570 32004 13580
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 31164 13188 31220 13198
rect 31164 13094 31220 13132
rect 30268 13074 30772 13076
rect 30268 13022 30270 13074
rect 30322 13022 30772 13074
rect 30268 13020 30772 13022
rect 30268 13010 30324 13020
rect 30716 12962 30772 13020
rect 30716 12910 30718 12962
rect 30770 12910 30772 12962
rect 30716 12898 30772 12910
rect 30156 12066 30212 12078
rect 30156 12014 30158 12066
rect 30210 12014 30212 12066
rect 30156 11954 30212 12014
rect 30156 11902 30158 11954
rect 30210 11902 30212 11954
rect 30156 11890 30212 11902
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 30268 11508 30324 11518
rect 30268 11414 30324 11452
rect 33068 11394 33124 11406
rect 33068 11342 33070 11394
rect 33122 11342 33124 11394
rect 31388 11284 31444 11294
rect 31388 10834 31444 11228
rect 32396 11284 32452 11294
rect 32396 11190 32452 11228
rect 31388 10782 31390 10834
rect 31442 10782 31444 10834
rect 31388 10770 31444 10782
rect 31164 10610 31220 10622
rect 31164 10558 31166 10610
rect 31218 10558 31220 10610
rect 31164 10050 31220 10558
rect 31164 9998 31166 10050
rect 31218 9998 31220 10050
rect 31164 9986 31220 9998
rect 30044 9886 30046 9938
rect 30098 9886 30100 9938
rect 29596 8260 29652 8270
rect 30044 8260 30100 9886
rect 31724 9940 31780 9950
rect 31724 9846 31780 9884
rect 31500 9828 31556 9838
rect 31388 9772 31500 9828
rect 30828 9716 30884 9726
rect 30828 9622 30884 9660
rect 31276 8932 31332 8942
rect 31052 8930 31332 8932
rect 31052 8878 31278 8930
rect 31330 8878 31332 8930
rect 31052 8876 31332 8878
rect 30156 8484 30212 8494
rect 30156 8372 30212 8428
rect 30156 8316 30436 8372
rect 29596 8258 30100 8260
rect 29596 8206 29598 8258
rect 29650 8206 30100 8258
rect 29596 8204 30100 8206
rect 29596 8194 29652 8204
rect 28028 8036 28084 8046
rect 27356 8034 28084 8036
rect 27356 7982 28030 8034
rect 28082 7982 28084 8034
rect 27356 7980 28084 7982
rect 27356 6692 27412 7980
rect 28028 7970 28084 7980
rect 30044 7700 30100 8204
rect 30044 7634 30100 7644
rect 27692 7588 27748 7598
rect 28028 7588 28084 7598
rect 27748 7586 28084 7588
rect 27748 7534 28030 7586
rect 28082 7534 28084 7586
rect 27748 7532 28084 7534
rect 27692 7522 27748 7532
rect 28028 7522 28084 7532
rect 30156 7364 30212 7374
rect 30156 7270 30212 7308
rect 27356 6626 27412 6636
rect 30380 6690 30436 8316
rect 30940 8036 30996 8046
rect 30604 8034 30996 8036
rect 30604 7982 30942 8034
rect 30994 7982 30996 8034
rect 30604 7980 30996 7982
rect 30604 7474 30660 7980
rect 30940 7970 30996 7980
rect 31052 7812 31108 8876
rect 31276 8866 31332 8876
rect 31276 8260 31332 8270
rect 31388 8260 31444 9772
rect 31500 9734 31556 9772
rect 32172 9828 32228 9838
rect 32172 9734 32228 9772
rect 31948 9044 32004 9054
rect 32508 9044 32564 9054
rect 33068 9044 33124 11342
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 31948 9042 33124 9044
rect 31948 8990 31950 9042
rect 32002 8990 32510 9042
rect 32562 8990 33124 9042
rect 31948 8988 33124 8990
rect 37212 9716 37268 33292
rect 37324 33124 37380 33134
rect 37324 33122 37492 33124
rect 37324 33070 37326 33122
rect 37378 33070 37492 33122
rect 37324 33068 37492 33070
rect 37324 33058 37380 33068
rect 37436 32674 37492 33068
rect 37436 32622 37438 32674
rect 37490 32622 37492 32674
rect 37436 32610 37492 32622
rect 38220 32562 38276 34300
rect 38220 32510 38222 32562
rect 38274 32510 38276 32562
rect 37324 31554 37380 31566
rect 37324 31502 37326 31554
rect 37378 31502 37380 31554
rect 37324 29540 37380 31502
rect 38220 31554 38276 32510
rect 38220 31502 38222 31554
rect 38274 31502 38276 31554
rect 38220 30884 38276 31502
rect 37436 29540 37492 29550
rect 37324 29538 37492 29540
rect 37324 29486 37438 29538
rect 37490 29486 37492 29538
rect 37324 29484 37492 29486
rect 37436 29474 37492 29484
rect 38220 29426 38276 30828
rect 38220 29374 38222 29426
rect 38274 29374 38276 29426
rect 38220 28418 38276 29374
rect 38220 28366 38222 28418
rect 38274 28366 38276 28418
rect 38220 27188 38276 28366
rect 38220 26962 38276 27132
rect 38220 26910 38222 26962
rect 38274 26910 38276 26962
rect 37324 26852 37380 26862
rect 37324 26850 37492 26852
rect 37324 26798 37326 26850
rect 37378 26798 37492 26850
rect 37324 26796 37492 26798
rect 37324 26786 37380 26796
rect 37436 26402 37492 26796
rect 37436 26350 37438 26402
rect 37490 26350 37492 26402
rect 37436 26338 37492 26350
rect 38220 26290 38276 26910
rect 38220 26238 38222 26290
rect 38274 26238 38276 26290
rect 38220 26226 38276 26238
rect 37324 25620 37380 25630
rect 37324 25618 37940 25620
rect 37324 25566 37326 25618
rect 37378 25566 37940 25618
rect 37324 25564 37940 25566
rect 37324 25554 37380 25564
rect 37548 25396 37604 25406
rect 37548 25302 37604 25340
rect 37884 25394 37940 25564
rect 37884 25342 37886 25394
rect 37938 25342 37940 25394
rect 37884 25330 37940 25342
rect 38220 25394 38276 25406
rect 38220 25342 38222 25394
rect 38274 25342 38276 25394
rect 38220 25172 38276 25342
rect 37884 24948 37940 24958
rect 37884 24610 37940 24892
rect 37884 24558 37886 24610
rect 37938 24558 37940 24610
rect 37884 24546 37940 24558
rect 38220 24052 38276 25116
rect 38332 24052 38388 24062
rect 38220 24050 38388 24052
rect 38220 23998 38334 24050
rect 38386 23998 38388 24050
rect 38220 23996 38388 23998
rect 38332 23986 38388 23996
rect 37772 21588 37828 21598
rect 37828 21532 38164 21588
rect 37772 21494 37828 21532
rect 38108 20018 38164 21532
rect 38108 19966 38110 20018
rect 38162 19966 38164 20018
rect 37436 19908 37492 19918
rect 37324 19906 37492 19908
rect 37324 19854 37438 19906
rect 37490 19854 37492 19906
rect 37324 19852 37492 19854
rect 37324 19122 37380 19852
rect 37436 19842 37492 19852
rect 37324 19070 37326 19122
rect 37378 19070 37380 19122
rect 37324 19058 37380 19070
rect 38108 18450 38164 19966
rect 38108 18398 38110 18450
rect 38162 18398 38164 18450
rect 37436 18340 37492 18350
rect 37436 18246 37492 18284
rect 38108 17668 38164 18398
rect 38108 17602 38164 17612
rect 31948 8484 32004 8988
rect 32508 8978 32564 8988
rect 37212 8930 37268 9660
rect 37212 8878 37214 8930
rect 37266 8878 37268 8930
rect 37212 8866 37268 8878
rect 38220 9042 38276 9054
rect 38220 8990 38222 9042
rect 38274 8990 38276 9042
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 38220 8596 38276 8990
rect 38332 8596 38388 8606
rect 38220 8540 38332 8596
rect 31948 8418 32004 8428
rect 38332 8370 38388 8540
rect 38332 8318 38334 8370
rect 38386 8318 38388 8370
rect 38332 8306 38388 8318
rect 31276 8258 31444 8260
rect 31276 8206 31278 8258
rect 31330 8206 31444 8258
rect 31276 8204 31444 8206
rect 31500 8258 31556 8270
rect 31500 8206 31502 8258
rect 31554 8206 31556 8258
rect 31276 8036 31332 8204
rect 31276 7970 31332 7980
rect 30828 7756 31108 7812
rect 30828 7698 30884 7756
rect 30828 7646 30830 7698
rect 30882 7646 30884 7698
rect 30828 7634 30884 7646
rect 31388 7700 31444 7710
rect 31388 7606 31444 7644
rect 30604 7422 30606 7474
rect 30658 7422 30660 7474
rect 30604 7410 30660 7422
rect 31500 7364 31556 8206
rect 31948 8036 32004 8046
rect 31948 7942 32004 7980
rect 31500 7298 31556 7308
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 30380 6638 30382 6690
rect 30434 6638 30436 6690
rect 30380 6626 30436 6638
rect 35196 5516 35460 5526
rect 27356 5460 27412 5470
rect 27244 5404 27356 5460
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 27356 5394 27412 5404
rect 27020 5182 27022 5234
rect 27074 5182 27076 5234
rect 27020 5170 27076 5182
rect 27692 5236 27748 5246
rect 27692 5124 27748 5180
rect 27468 5068 27748 5124
rect 27468 5010 27524 5068
rect 27468 4958 27470 5010
rect 27522 4958 27524 5010
rect 27468 4946 27524 4958
rect 34412 4338 34468 4350
rect 34412 4286 34414 4338
rect 34466 4286 34468 4338
rect 26572 3614 26574 3666
rect 26626 3614 26628 3666
rect 26572 3602 26628 3614
rect 33964 4114 34020 4126
rect 33964 4062 33966 4114
rect 34018 4062 34020 4114
rect 27468 3554 27524 3566
rect 27468 3502 27470 3554
rect 27522 3502 27524 3554
rect 25900 2942 25902 2994
rect 25954 2942 25956 2994
rect 25900 2930 25956 2942
rect 26236 3052 26516 3108
rect 26908 3442 26964 3454
rect 26908 3390 26910 3442
rect 26962 3390 26964 3442
rect 25340 2882 25396 2894
rect 25788 2884 25844 2894
rect 26236 2884 26292 3052
rect 25340 2830 25342 2882
rect 25394 2830 25396 2882
rect 22652 1986 22932 1988
rect 22652 1934 22878 1986
rect 22930 1934 22932 1986
rect 22652 1932 22932 1934
rect 22316 1876 22372 1886
rect 22204 1874 22372 1876
rect 22204 1822 22318 1874
rect 22370 1822 22372 1874
rect 22204 1820 22372 1822
rect 22316 1810 22372 1820
rect 22652 400 22708 1932
rect 22876 1922 22932 1932
rect 23212 2772 23268 2782
rect 23212 1874 23268 2716
rect 25228 2772 25284 2782
rect 25228 2678 25284 2716
rect 24332 2658 24388 2670
rect 24332 2606 24334 2658
rect 24386 2606 24388 2658
rect 23660 1988 23716 1998
rect 23660 1894 23716 1932
rect 23212 1822 23214 1874
rect 23266 1822 23268 1874
rect 23212 1810 23268 1822
rect 24332 1540 24388 2606
rect 24780 2658 24836 2670
rect 24780 2606 24782 2658
rect 24834 2606 24836 2658
rect 24556 1874 24612 1886
rect 24556 1822 24558 1874
rect 24610 1822 24612 1874
rect 24556 1540 24612 1822
rect 24780 1652 24836 2606
rect 25340 2324 25396 2830
rect 24892 2268 25396 2324
rect 25564 2828 25788 2884
rect 24892 1874 24948 2268
rect 25228 1876 25284 1886
rect 24892 1822 24894 1874
rect 24946 1822 24948 1874
rect 24892 1810 24948 1822
rect 25116 1874 25284 1876
rect 25116 1822 25230 1874
rect 25282 1822 25284 1874
rect 25116 1820 25284 1822
rect 25116 1652 25172 1820
rect 25228 1810 25284 1820
rect 25564 1874 25620 2828
rect 25788 2818 25844 2828
rect 26124 2828 26292 2884
rect 26796 2884 26852 2894
rect 25564 1822 25566 1874
rect 25618 1822 25620 1874
rect 25564 1810 25620 1822
rect 26012 1988 26068 1998
rect 26124 1988 26180 2828
rect 26796 2790 26852 2828
rect 26012 1986 26180 1988
rect 26012 1934 26014 1986
rect 26066 1934 26180 1986
rect 26012 1932 26180 1934
rect 26348 2770 26404 2782
rect 26348 2718 26350 2770
rect 26402 2718 26404 2770
rect 24780 1596 25172 1652
rect 24220 1484 24612 1540
rect 23548 476 23828 532
rect 23548 400 23604 476
rect 3808 0 3920 400
rect 4704 0 4816 400
rect 5600 0 5712 400
rect 6496 0 6608 400
rect 7392 0 7504 400
rect 8288 0 8400 400
rect 9184 0 9296 400
rect 10080 0 10192 400
rect 10976 0 11088 400
rect 11872 0 11984 400
rect 12768 0 12880 400
rect 13664 0 13776 400
rect 14560 0 14672 400
rect 15456 0 15568 400
rect 16352 0 16464 400
rect 17248 0 17360 400
rect 18144 0 18256 400
rect 19040 0 19152 400
rect 19936 0 20048 400
rect 20832 0 20944 400
rect 21728 0 21840 400
rect 22624 0 22736 400
rect 23520 0 23632 400
rect 23772 308 23828 476
rect 24220 308 24276 1484
rect 24444 476 24724 532
rect 24444 400 24500 476
rect 23772 252 24276 308
rect 24416 0 24528 400
rect 24668 308 24724 476
rect 25116 308 25172 1596
rect 25340 476 25732 532
rect 25340 400 25396 476
rect 24668 252 25172 308
rect 25312 0 25424 400
rect 25676 308 25732 476
rect 26012 308 26068 1932
rect 26236 1876 26292 1886
rect 26348 1876 26404 2718
rect 26236 1874 26404 1876
rect 26236 1822 26238 1874
rect 26290 1822 26404 1874
rect 26236 1820 26404 1822
rect 26572 2660 26628 2670
rect 26572 1874 26628 2604
rect 26908 2100 26964 3390
rect 27020 3332 27076 3342
rect 27020 3238 27076 3276
rect 27356 2660 27412 2670
rect 27356 2566 27412 2604
rect 26908 2044 27412 2100
rect 26572 1822 26574 1874
rect 26626 1822 26628 1874
rect 26236 1810 26292 1820
rect 26572 1540 26628 1822
rect 27356 1874 27412 2044
rect 27356 1822 27358 1874
rect 27410 1822 27412 1874
rect 27356 1810 27412 1822
rect 26908 1764 26964 1774
rect 26908 1762 27300 1764
rect 26908 1710 26910 1762
rect 26962 1710 27300 1762
rect 26908 1708 27300 1710
rect 26908 1698 26964 1708
rect 27244 1652 27300 1708
rect 27468 1652 27524 3502
rect 27916 3554 27972 3566
rect 27916 3502 27918 3554
rect 27970 3502 27972 3554
rect 27804 2658 27860 2670
rect 27804 2606 27806 2658
rect 27858 2606 27860 2658
rect 27244 1596 27524 1652
rect 27580 1988 27636 1998
rect 27804 1988 27860 2606
rect 27580 1986 27860 1988
rect 27580 1934 27582 1986
rect 27634 1934 27860 1986
rect 27580 1932 27860 1934
rect 26236 1484 26628 1540
rect 26236 400 26292 1484
rect 27580 1428 27636 1932
rect 27916 1764 27972 3502
rect 31052 3554 31108 3566
rect 31052 3502 31054 3554
rect 31106 3502 31108 3554
rect 28476 3442 28532 3454
rect 28476 3390 28478 3442
rect 28530 3390 28532 3442
rect 28364 2658 28420 2670
rect 28364 2606 28366 2658
rect 28418 2606 28420 2658
rect 28364 1876 28420 2606
rect 27916 1698 27972 1708
rect 28028 1874 28420 1876
rect 28028 1822 28366 1874
rect 28418 1822 28420 1874
rect 28028 1820 28420 1822
rect 28476 1876 28532 3390
rect 31052 2884 31108 3502
rect 33180 3554 33236 3566
rect 33180 3502 33182 3554
rect 33234 3502 33236 3554
rect 30604 2828 31108 2884
rect 31164 3442 31220 3454
rect 31164 3390 31166 3442
rect 31218 3390 31220 3442
rect 28924 2658 28980 2670
rect 28924 2606 28926 2658
rect 28978 2606 28980 2658
rect 28700 1876 28756 1886
rect 28476 1874 28756 1876
rect 28476 1822 28702 1874
rect 28754 1822 28756 1874
rect 28476 1820 28756 1822
rect 27132 1372 27636 1428
rect 27132 400 27188 1372
rect 28028 400 28084 1820
rect 28364 1810 28420 1820
rect 28700 1810 28756 1820
rect 28924 1540 28980 2606
rect 29820 2658 29876 2670
rect 29820 2606 29822 2658
rect 29874 2606 29876 2658
rect 29372 1986 29428 1998
rect 29372 1934 29374 1986
rect 29426 1934 29428 1986
rect 29148 1764 29204 1774
rect 29148 1670 29204 1708
rect 29372 1540 29428 1934
rect 28924 1484 29428 1540
rect 29820 1876 29876 2606
rect 30044 1876 30100 1886
rect 29820 1874 30100 1876
rect 29820 1822 30046 1874
rect 30098 1822 30100 1874
rect 29820 1820 30100 1822
rect 28924 400 28980 1484
rect 29820 400 29876 1820
rect 30044 1810 30100 1820
rect 30380 1876 30436 1886
rect 30604 1876 30660 2828
rect 30380 1874 30660 1876
rect 30380 1822 30382 1874
rect 30434 1822 30660 1874
rect 30380 1820 30660 1822
rect 30716 2658 30772 2670
rect 30716 2606 30718 2658
rect 30770 2606 30772 2658
rect 30716 1876 30772 2606
rect 30940 1876 30996 1886
rect 30716 1874 30996 1876
rect 30716 1822 30942 1874
rect 30994 1822 30996 1874
rect 30716 1820 30996 1822
rect 31164 1876 31220 3390
rect 32508 3444 32564 3454
rect 31948 2658 32004 2670
rect 31948 2606 31950 2658
rect 32002 2606 32004 2658
rect 31948 1988 32004 2606
rect 32172 1988 32228 1998
rect 31948 1986 32228 1988
rect 31948 1934 32174 1986
rect 32226 1934 32228 1986
rect 31948 1932 32228 1934
rect 31276 1876 31332 1886
rect 31164 1874 31332 1876
rect 31164 1822 31278 1874
rect 31330 1822 31332 1874
rect 31164 1820 31332 1822
rect 30380 1810 30436 1820
rect 30716 400 30772 1820
rect 30940 1810 30996 1820
rect 31276 1810 31332 1820
rect 31948 1764 32004 1932
rect 32172 1922 32228 1932
rect 32508 1874 32564 3388
rect 33180 3388 33236 3502
rect 33628 3444 33684 3482
rect 33068 3330 33124 3342
rect 33180 3332 33348 3388
rect 33628 3378 33684 3388
rect 33068 3278 33070 3330
rect 33122 3278 33124 3330
rect 33068 2770 33124 3278
rect 33068 2718 33070 2770
rect 33122 2718 33124 2770
rect 33068 2706 33124 2718
rect 32508 1822 32510 1874
rect 32562 1822 32564 1874
rect 32508 1810 32564 1822
rect 32620 2658 32676 2670
rect 32620 2606 32622 2658
rect 32674 2606 32676 2658
rect 31612 1708 32004 1764
rect 31612 400 31668 1708
rect 32620 1540 32676 2606
rect 33180 2548 33236 2558
rect 33180 2454 33236 2492
rect 32844 1874 32900 1886
rect 32844 1822 32846 1874
rect 32898 1822 32900 1874
rect 32844 1540 32900 1822
rect 33180 1876 33236 1886
rect 33292 1876 33348 3332
rect 33964 2882 34020 4062
rect 34412 2996 34468 4286
rect 34748 4338 34804 4350
rect 34748 4286 34750 4338
rect 34802 4286 34804 4338
rect 34412 2930 34468 2940
rect 34524 4226 34580 4238
rect 34524 4174 34526 4226
rect 34578 4174 34580 4226
rect 33964 2830 33966 2882
rect 34018 2830 34020 2882
rect 33964 2818 34020 2830
rect 33740 1988 33796 1998
rect 33180 1874 33348 1876
rect 33180 1822 33182 1874
rect 33234 1822 33348 1874
rect 33180 1820 33348 1822
rect 33404 1932 33740 1988
rect 33180 1810 33236 1820
rect 32508 1484 32900 1540
rect 32508 400 32564 1484
rect 33404 400 33460 1932
rect 33740 1894 33796 1932
rect 34524 1874 34580 4174
rect 34748 3108 34804 4286
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 34748 3042 34804 3052
rect 36652 3108 36708 3118
rect 35980 2996 36036 3006
rect 34748 2772 34804 2782
rect 34524 1822 34526 1874
rect 34578 1822 34580 1874
rect 34524 1810 34580 1822
rect 34636 2770 34804 2772
rect 34636 2718 34750 2770
rect 34802 2718 34804 2770
rect 34636 2716 34804 2718
rect 33964 1764 34020 1774
rect 33964 1762 34468 1764
rect 33964 1710 33966 1762
rect 34018 1710 34468 1762
rect 33964 1708 34468 1710
rect 33964 1698 34020 1708
rect 34412 1652 34468 1708
rect 34636 1652 34692 2716
rect 34748 2706 34804 2716
rect 34412 1596 34692 1652
rect 34860 2660 34916 2670
rect 34860 1986 34916 2604
rect 35196 2380 35460 2390
rect 35252 2324 35300 2380
rect 35356 2324 35404 2380
rect 35196 2314 35460 2324
rect 34860 1934 34862 1986
rect 34914 1934 34916 1986
rect 34300 476 34580 532
rect 34300 400 34356 476
rect 25676 252 26068 308
rect 26208 0 26320 400
rect 27104 0 27216 400
rect 28000 0 28112 400
rect 28896 0 29008 400
rect 29792 0 29904 400
rect 30688 0 30800 400
rect 31584 0 31696 400
rect 32480 0 32592 400
rect 33376 0 33488 400
rect 34272 0 34384 400
rect 34524 308 34580 476
rect 34860 308 34916 1934
rect 35308 1988 35364 1998
rect 35308 1894 35364 1932
rect 35196 1876 35252 1886
rect 35196 400 35252 1820
rect 35980 1874 36036 2940
rect 36092 2660 36148 2670
rect 36092 2566 36148 2604
rect 36540 2658 36596 2670
rect 36540 2606 36542 2658
rect 36594 2606 36596 2658
rect 35980 1822 35982 1874
rect 36034 1822 36036 1874
rect 35980 1810 36036 1822
rect 36204 1988 36260 1998
rect 36540 1988 36596 2606
rect 36204 1986 36596 1988
rect 36204 1934 36206 1986
rect 36258 1934 36596 1986
rect 36204 1932 36596 1934
rect 36204 1876 36260 1932
rect 36204 1810 36260 1820
rect 36652 1874 36708 3052
rect 36652 1822 36654 1874
rect 36706 1822 36708 1874
rect 36652 1810 36708 1822
rect 36876 1986 36932 1998
rect 36876 1934 36878 1986
rect 36930 1934 36932 1986
rect 36092 1764 36148 1774
rect 36092 400 36148 1708
rect 36876 1764 36932 1934
rect 36876 1698 36932 1708
rect 37436 1764 37492 1774
rect 37436 1670 37492 1708
rect 34524 252 34916 308
rect 35168 0 35280 400
rect 36064 0 36176 400
<< via2 >>
rect 4476 98026 4532 98028
rect 4476 97974 4478 98026
rect 4478 97974 4530 98026
rect 4530 97974 4532 98026
rect 4476 97972 4532 97974
rect 4580 98026 4636 98028
rect 4580 97974 4582 98026
rect 4582 97974 4634 98026
rect 4634 97974 4636 98026
rect 4580 97972 4636 97974
rect 4684 98026 4740 98028
rect 4684 97974 4686 98026
rect 4686 97974 4738 98026
rect 4738 97974 4740 98026
rect 4684 97972 4740 97974
rect 13020 97522 13076 97524
rect 13020 97470 13022 97522
rect 13022 97470 13074 97522
rect 13074 97470 13076 97522
rect 13020 97468 13076 97470
rect 13692 97356 13748 97412
rect 14476 97468 14532 97524
rect 6188 96572 6244 96628
rect 4476 96458 4532 96460
rect 4476 96406 4478 96458
rect 4478 96406 4530 96458
rect 4530 96406 4532 96458
rect 4476 96404 4532 96406
rect 4580 96458 4636 96460
rect 4580 96406 4582 96458
rect 4582 96406 4634 96458
rect 4634 96406 4636 96458
rect 4580 96404 4636 96406
rect 4684 96458 4740 96460
rect 4684 96406 4686 96458
rect 4686 96406 4738 96458
rect 4738 96406 4740 96458
rect 4684 96404 4740 96406
rect 1708 94386 1764 94388
rect 1708 94334 1710 94386
rect 1710 94334 1762 94386
rect 1762 94334 1764 94386
rect 1708 94332 1764 94334
rect 6860 96626 6916 96628
rect 6860 96574 6862 96626
rect 6862 96574 6914 96626
rect 6914 96574 6916 96626
rect 6860 96572 6916 96574
rect 7644 96572 7700 96628
rect 2940 93660 2996 93716
rect 2044 93490 2100 93492
rect 2044 93438 2046 93490
rect 2046 93438 2098 93490
rect 2098 93438 2100 93490
rect 2044 93436 2100 93438
rect 4476 94890 4532 94892
rect 4476 94838 4478 94890
rect 4478 94838 4530 94890
rect 4530 94838 4532 94890
rect 4476 94836 4532 94838
rect 4580 94890 4636 94892
rect 4580 94838 4582 94890
rect 4582 94838 4634 94890
rect 4634 94838 4636 94890
rect 4580 94836 4636 94838
rect 4684 94890 4740 94892
rect 4684 94838 4686 94890
rect 4686 94838 4738 94890
rect 4738 94838 4740 94890
rect 4684 94836 4740 94838
rect 4172 93714 4228 93716
rect 4172 93662 4174 93714
rect 4174 93662 4226 93714
rect 4226 93662 4228 93714
rect 4172 93660 4228 93662
rect 3388 93436 3444 93492
rect 4476 93322 4532 93324
rect 4476 93270 4478 93322
rect 4478 93270 4530 93322
rect 4530 93270 4532 93322
rect 4476 93268 4532 93270
rect 4580 93322 4636 93324
rect 4580 93270 4582 93322
rect 4582 93270 4634 93322
rect 4634 93270 4636 93322
rect 4580 93268 4636 93270
rect 4684 93322 4740 93324
rect 4684 93270 4686 93322
rect 4686 93270 4738 93322
rect 4738 93270 4740 93322
rect 4684 93268 4740 93270
rect 6748 96066 6804 96068
rect 6748 96014 6750 96066
rect 6750 96014 6802 96066
rect 6802 96014 6804 96066
rect 6748 96012 6804 96014
rect 8876 96012 8932 96068
rect 9324 96066 9380 96068
rect 9324 96014 9326 96066
rect 9326 96014 9378 96066
rect 9378 96014 9380 96066
rect 9324 96012 9380 96014
rect 8652 95788 8708 95844
rect 9660 95788 9716 95844
rect 10332 95788 10388 95844
rect 11676 95842 11732 95844
rect 11676 95790 11678 95842
rect 11678 95790 11730 95842
rect 11730 95790 11732 95842
rect 11676 95788 11732 95790
rect 13580 95676 13636 95732
rect 12348 95506 12404 95508
rect 12348 95454 12350 95506
rect 12350 95454 12402 95506
rect 12402 95454 12404 95506
rect 12348 95452 12404 95454
rect 13916 95452 13972 95508
rect 15708 97410 15764 97412
rect 15708 97358 15710 97410
rect 15710 97358 15762 97410
rect 15762 97358 15764 97410
rect 15708 97356 15764 97358
rect 16156 97356 16212 97412
rect 14476 95452 14532 95508
rect 14700 95676 14756 95732
rect 16940 97410 16996 97412
rect 16940 97358 16942 97410
rect 16942 97358 16994 97410
rect 16994 97358 16996 97410
rect 16940 97356 16996 97358
rect 19836 97242 19892 97244
rect 19836 97190 19838 97242
rect 19838 97190 19890 97242
rect 19890 97190 19892 97242
rect 19836 97188 19892 97190
rect 19940 97242 19996 97244
rect 19940 97190 19942 97242
rect 19942 97190 19994 97242
rect 19994 97190 19996 97242
rect 19940 97188 19996 97190
rect 20044 97242 20100 97244
rect 20044 97190 20046 97242
rect 20046 97190 20098 97242
rect 20098 97190 20100 97242
rect 20044 97188 20100 97190
rect 16268 95676 16324 95732
rect 14700 94668 14756 94724
rect 15148 95506 15204 95508
rect 15148 95454 15150 95506
rect 15150 95454 15202 95506
rect 15202 95454 15204 95506
rect 15148 95452 15204 95454
rect 6748 93714 6804 93716
rect 6748 93662 6750 93714
rect 6750 93662 6802 93714
rect 6802 93662 6804 93714
rect 6748 93660 6804 93662
rect 6524 92540 6580 92596
rect 3836 92146 3892 92148
rect 3836 92094 3838 92146
rect 3838 92094 3890 92146
rect 3890 92094 3892 92146
rect 3836 92092 3892 92094
rect 4956 92092 5012 92148
rect 4476 91754 4532 91756
rect 4476 91702 4478 91754
rect 4478 91702 4530 91754
rect 4530 91702 4532 91754
rect 4476 91700 4532 91702
rect 4580 91754 4636 91756
rect 4580 91702 4582 91754
rect 4582 91702 4634 91754
rect 4634 91702 4636 91754
rect 4580 91700 4636 91702
rect 4684 91754 4740 91756
rect 4684 91702 4686 91754
rect 4686 91702 4738 91754
rect 4738 91702 4740 91754
rect 4684 91700 4740 91702
rect 6972 92540 7028 92596
rect 10332 93660 10388 93716
rect 7308 92428 7364 92484
rect 7756 92428 7812 92484
rect 9660 92818 9716 92820
rect 9660 92766 9662 92818
rect 9662 92766 9714 92818
rect 9714 92766 9716 92818
rect 9660 92764 9716 92766
rect 12012 93714 12068 93716
rect 12012 93662 12014 93714
rect 12014 93662 12066 93714
rect 12066 93662 12068 93714
rect 12012 93660 12068 93662
rect 13356 93714 13412 93716
rect 13356 93662 13358 93714
rect 13358 93662 13410 93714
rect 13410 93662 13412 93714
rect 13356 93660 13412 93662
rect 14140 93660 14196 93716
rect 12684 93602 12740 93604
rect 12684 93550 12686 93602
rect 12686 93550 12738 93602
rect 12738 93550 12740 93602
rect 12684 93548 12740 93550
rect 10780 92764 10836 92820
rect 9660 92428 9716 92484
rect 10780 92540 10836 92596
rect 10220 92258 10276 92260
rect 10220 92206 10222 92258
rect 10222 92206 10274 92258
rect 10274 92206 10276 92258
rect 10220 92204 10276 92206
rect 12572 92764 12628 92820
rect 12348 92146 12404 92148
rect 12348 92094 12350 92146
rect 12350 92094 12402 92146
rect 12402 92094 12404 92146
rect 12348 92092 12404 92094
rect 11564 91362 11620 91364
rect 11564 91310 11566 91362
rect 11566 91310 11618 91362
rect 11618 91310 11620 91362
rect 11564 91308 11620 91310
rect 12012 91362 12068 91364
rect 12012 91310 12014 91362
rect 12014 91310 12066 91362
rect 12066 91310 12068 91362
rect 12012 91308 12068 91310
rect 4476 90186 4532 90188
rect 4476 90134 4478 90186
rect 4478 90134 4530 90186
rect 4530 90134 4532 90186
rect 4476 90132 4532 90134
rect 4580 90186 4636 90188
rect 4580 90134 4582 90186
rect 4582 90134 4634 90186
rect 4634 90134 4636 90186
rect 4580 90132 4636 90134
rect 4684 90186 4740 90188
rect 4684 90134 4686 90186
rect 4686 90134 4738 90186
rect 4738 90134 4740 90186
rect 4684 90132 4740 90134
rect 3164 89740 3220 89796
rect 4284 89794 4340 89796
rect 4284 89742 4286 89794
rect 4286 89742 4338 89794
rect 4338 89742 4340 89794
rect 4284 89740 4340 89742
rect 11676 90636 11732 90692
rect 13804 92818 13860 92820
rect 13804 92766 13806 92818
rect 13806 92766 13858 92818
rect 13858 92766 13860 92818
rect 13804 92764 13860 92766
rect 14588 93548 14644 93604
rect 14252 92988 14308 93044
rect 13580 92316 13636 92372
rect 12908 92204 12964 92260
rect 12348 90636 12404 90692
rect 4476 88618 4532 88620
rect 4476 88566 4478 88618
rect 4478 88566 4530 88618
rect 4530 88566 4532 88618
rect 4476 88564 4532 88566
rect 4580 88618 4636 88620
rect 4580 88566 4582 88618
rect 4582 88566 4634 88618
rect 4634 88566 4636 88618
rect 4580 88564 4636 88566
rect 4684 88618 4740 88620
rect 4684 88566 4686 88618
rect 4686 88566 4738 88618
rect 4738 88566 4740 88618
rect 4684 88564 4740 88566
rect 6860 89010 6916 89012
rect 6860 88958 6862 89010
rect 6862 88958 6914 89010
rect 6914 88958 6916 89010
rect 6860 88956 6916 88958
rect 7980 88956 8036 89012
rect 7980 88172 8036 88228
rect 7756 87948 7812 88004
rect 8428 87948 8484 88004
rect 4476 87050 4532 87052
rect 4476 86998 4478 87050
rect 4478 86998 4530 87050
rect 4530 86998 4532 87050
rect 4476 86996 4532 86998
rect 4580 87050 4636 87052
rect 4580 86998 4582 87050
rect 4582 86998 4634 87050
rect 4634 86998 4636 87050
rect 4580 86996 4636 86998
rect 4684 87050 4740 87052
rect 4684 86998 4686 87050
rect 4686 86998 4738 87050
rect 4738 86998 4740 87050
rect 4684 86996 4740 86998
rect 4284 86492 4340 86548
rect 6972 87164 7028 87220
rect 13580 91362 13636 91364
rect 13580 91310 13582 91362
rect 13582 91310 13634 91362
rect 13634 91310 13636 91362
rect 13580 91308 13636 91310
rect 16828 95394 16884 95396
rect 16828 95342 16830 95394
rect 16830 95342 16882 95394
rect 16882 95342 16884 95394
rect 16828 95340 16884 95342
rect 17500 95340 17556 95396
rect 15596 94668 15652 94724
rect 17500 94444 17556 94500
rect 17276 93996 17332 94052
rect 15932 93660 15988 93716
rect 16604 93714 16660 93716
rect 16604 93662 16606 93714
rect 16606 93662 16658 93714
rect 16658 93662 16660 93714
rect 16604 93660 16660 93662
rect 14364 92316 14420 92372
rect 14700 92258 14756 92260
rect 14700 92206 14702 92258
rect 14702 92206 14754 92258
rect 14754 92206 14756 92258
rect 14700 92204 14756 92206
rect 15148 92258 15204 92260
rect 15148 92206 15150 92258
rect 15150 92206 15202 92258
rect 15202 92206 15204 92258
rect 15148 92204 15204 92206
rect 17052 93660 17108 93716
rect 17724 93996 17780 94052
rect 19516 95676 19572 95732
rect 19836 95674 19892 95676
rect 19836 95622 19838 95674
rect 19838 95622 19890 95674
rect 19890 95622 19892 95674
rect 19836 95620 19892 95622
rect 19940 95674 19996 95676
rect 19940 95622 19942 95674
rect 19942 95622 19994 95674
rect 19994 95622 19996 95674
rect 19940 95620 19996 95622
rect 20044 95674 20100 95676
rect 20044 95622 20046 95674
rect 20046 95622 20098 95674
rect 20098 95622 20100 95674
rect 20044 95620 20100 95622
rect 20636 95228 20692 95284
rect 18508 94498 18564 94500
rect 18508 94446 18510 94498
rect 18510 94446 18562 94498
rect 18562 94446 18564 94498
rect 18508 94444 18564 94446
rect 18396 93714 18452 93716
rect 18396 93662 18398 93714
rect 18398 93662 18450 93714
rect 18450 93662 18452 93714
rect 18396 93660 18452 93662
rect 19292 93660 19348 93716
rect 17724 93324 17780 93380
rect 20300 94332 20356 94388
rect 19836 94106 19892 94108
rect 19836 94054 19838 94106
rect 19838 94054 19890 94106
rect 19890 94054 19892 94106
rect 19836 94052 19892 94054
rect 19940 94106 19996 94108
rect 19940 94054 19942 94106
rect 19942 94054 19994 94106
rect 19994 94054 19996 94106
rect 19940 94052 19996 94054
rect 20044 94106 20100 94108
rect 20044 94054 20046 94106
rect 20046 94054 20098 94106
rect 20098 94054 20100 94106
rect 20044 94052 20100 94054
rect 20636 93938 20692 93940
rect 20636 93886 20638 93938
rect 20638 93886 20690 93938
rect 20690 93886 20692 93938
rect 20636 93884 20692 93886
rect 20076 93324 20132 93380
rect 17276 93042 17332 93044
rect 17276 92990 17278 93042
rect 17278 92990 17330 93042
rect 17330 92990 17332 93042
rect 17276 92988 17332 92990
rect 18620 93042 18676 93044
rect 18620 92990 18622 93042
rect 18622 92990 18674 93042
rect 18674 92990 18676 93042
rect 18620 92988 18676 92990
rect 17948 92652 18004 92708
rect 19404 92652 19460 92708
rect 19836 92538 19892 92540
rect 19836 92486 19838 92538
rect 19838 92486 19890 92538
rect 19890 92486 19892 92538
rect 19836 92484 19892 92486
rect 19940 92538 19996 92540
rect 19940 92486 19942 92538
rect 19942 92486 19994 92538
rect 19994 92486 19996 92538
rect 19940 92484 19996 92486
rect 20044 92538 20100 92540
rect 20044 92486 20046 92538
rect 20046 92486 20098 92538
rect 20098 92486 20100 92538
rect 20044 92484 20100 92486
rect 16828 92204 16884 92260
rect 20748 93324 20804 93380
rect 19836 90970 19892 90972
rect 19836 90918 19838 90970
rect 19838 90918 19890 90970
rect 19890 90918 19892 90970
rect 19836 90916 19892 90918
rect 19940 90970 19996 90972
rect 19940 90918 19942 90970
rect 19942 90918 19994 90970
rect 19994 90918 19996 90970
rect 19940 90916 19996 90918
rect 20044 90970 20100 90972
rect 20044 90918 20046 90970
rect 20046 90918 20098 90970
rect 20098 90918 20100 90970
rect 20044 90916 20100 90918
rect 13356 89010 13412 89012
rect 13356 88958 13358 89010
rect 13358 88958 13410 89010
rect 13410 88958 13412 89010
rect 13356 88956 13412 88958
rect 9324 88060 9380 88116
rect 9660 88226 9716 88228
rect 9660 88174 9662 88226
rect 9662 88174 9714 88226
rect 9714 88174 9716 88226
rect 9660 88172 9716 88174
rect 9548 87836 9604 87892
rect 9100 87164 9156 87220
rect 10556 88060 10612 88116
rect 10556 87500 10612 87556
rect 10668 87948 10724 88004
rect 9324 86658 9380 86660
rect 9324 86606 9326 86658
rect 9326 86606 9378 86658
rect 9378 86606 9380 86658
rect 9324 86604 9380 86606
rect 10108 86658 10164 86660
rect 10108 86606 10110 86658
rect 10110 86606 10162 86658
rect 10162 86606 10164 86658
rect 10108 86604 10164 86606
rect 12236 88002 12292 88004
rect 12236 87950 12238 88002
rect 12238 87950 12290 88002
rect 12290 87950 12292 88002
rect 12236 87948 12292 87950
rect 12012 87836 12068 87892
rect 12460 87724 12516 87780
rect 10892 86546 10948 86548
rect 10892 86494 10894 86546
rect 10894 86494 10946 86546
rect 10946 86494 10948 86546
rect 10892 86492 10948 86494
rect 5404 85874 5460 85876
rect 5404 85822 5406 85874
rect 5406 85822 5458 85874
rect 5458 85822 5460 85874
rect 5404 85820 5460 85822
rect 4476 85482 4532 85484
rect 4476 85430 4478 85482
rect 4478 85430 4530 85482
rect 4530 85430 4532 85482
rect 4476 85428 4532 85430
rect 4580 85482 4636 85484
rect 4580 85430 4582 85482
rect 4582 85430 4634 85482
rect 4634 85430 4636 85482
rect 4580 85428 4636 85430
rect 4684 85482 4740 85484
rect 4684 85430 4686 85482
rect 4686 85430 4738 85482
rect 4738 85430 4740 85482
rect 4684 85428 4740 85430
rect 11564 86044 11620 86100
rect 12124 86098 12180 86100
rect 12124 86046 12126 86098
rect 12126 86046 12178 86098
rect 12178 86046 12180 86098
rect 12124 86044 12180 86046
rect 13804 88002 13860 88004
rect 13804 87950 13806 88002
rect 13806 87950 13858 88002
rect 13858 87950 13860 88002
rect 13804 87948 13860 87950
rect 13580 87554 13636 87556
rect 13580 87502 13582 87554
rect 13582 87502 13634 87554
rect 13634 87502 13636 87554
rect 13580 87500 13636 87502
rect 13020 87442 13076 87444
rect 13020 87390 13022 87442
rect 13022 87390 13074 87442
rect 13074 87390 13076 87442
rect 13020 87388 13076 87390
rect 12796 86044 12852 86100
rect 19964 89794 20020 89796
rect 19964 89742 19966 89794
rect 19966 89742 20018 89794
rect 20018 89742 20020 89794
rect 19964 89740 20020 89742
rect 14252 89068 14308 89124
rect 17500 89516 17556 89572
rect 15932 89068 15988 89124
rect 16716 89122 16772 89124
rect 16716 89070 16718 89122
rect 16718 89070 16770 89122
rect 16770 89070 16772 89122
rect 16716 89068 16772 89070
rect 16044 88956 16100 89012
rect 14252 88002 14308 88004
rect 14252 87950 14254 88002
rect 14254 87950 14306 88002
rect 14306 87950 14308 88002
rect 14252 87948 14308 87950
rect 14140 87724 14196 87780
rect 15260 87666 15316 87668
rect 15260 87614 15262 87666
rect 15262 87614 15314 87666
rect 15314 87614 15316 87666
rect 15260 87612 15316 87614
rect 13916 87442 13972 87444
rect 13916 87390 13918 87442
rect 13918 87390 13970 87442
rect 13970 87390 13972 87442
rect 13916 87388 13972 87390
rect 15708 87666 15764 87668
rect 15708 87614 15710 87666
rect 15710 87614 15762 87666
rect 15762 87614 15764 87666
rect 15708 87612 15764 87614
rect 15596 87442 15652 87444
rect 15596 87390 15598 87442
rect 15598 87390 15650 87442
rect 15650 87390 15652 87442
rect 15596 87388 15652 87390
rect 14140 86492 14196 86548
rect 6972 85874 7028 85876
rect 6972 85822 6974 85874
rect 6974 85822 7026 85874
rect 7026 85822 7028 85874
rect 6972 85820 7028 85822
rect 12908 84866 12964 84868
rect 12908 84814 12910 84866
rect 12910 84814 12962 84866
rect 12962 84814 12964 84866
rect 12908 84812 12964 84814
rect 4956 84476 5012 84532
rect 4476 83914 4532 83916
rect 4476 83862 4478 83914
rect 4478 83862 4530 83914
rect 4530 83862 4532 83914
rect 4476 83860 4532 83862
rect 4580 83914 4636 83916
rect 4580 83862 4582 83914
rect 4582 83862 4634 83914
rect 4634 83862 4636 83914
rect 4580 83860 4636 83862
rect 4684 83914 4740 83916
rect 4684 83862 4686 83914
rect 4686 83862 4738 83914
rect 4738 83862 4740 83914
rect 4684 83860 4740 83862
rect 3276 83356 3332 83412
rect 4396 83356 4452 83412
rect 4956 82572 5012 82628
rect 6076 82626 6132 82628
rect 6076 82574 6078 82626
rect 6078 82574 6130 82626
rect 6130 82574 6132 82626
rect 6076 82572 6132 82574
rect 7196 82460 7252 82516
rect 4476 82346 4532 82348
rect 4476 82294 4478 82346
rect 4478 82294 4530 82346
rect 4530 82294 4532 82346
rect 4476 82292 4532 82294
rect 4580 82346 4636 82348
rect 4580 82294 4582 82346
rect 4582 82294 4634 82346
rect 4634 82294 4636 82346
rect 4580 82292 4636 82294
rect 4684 82346 4740 82348
rect 4684 82294 4686 82346
rect 4686 82294 4738 82346
rect 4738 82294 4740 82346
rect 4684 82292 4740 82294
rect 6636 81954 6692 81956
rect 6636 81902 6638 81954
rect 6638 81902 6690 81954
rect 6690 81902 6692 81954
rect 6636 81900 6692 81902
rect 4844 81228 4900 81284
rect 5852 81730 5908 81732
rect 5852 81678 5854 81730
rect 5854 81678 5906 81730
rect 5906 81678 5908 81730
rect 5852 81676 5908 81678
rect 8428 82908 8484 82964
rect 7980 82460 8036 82516
rect 12572 84194 12628 84196
rect 12572 84142 12574 84194
rect 12574 84142 12626 84194
rect 12626 84142 12628 84194
rect 12572 84140 12628 84142
rect 8764 82460 8820 82516
rect 7196 81676 7252 81732
rect 6524 81340 6580 81396
rect 4476 80778 4532 80780
rect 4476 80726 4478 80778
rect 4478 80726 4530 80778
rect 4530 80726 4532 80778
rect 4476 80724 4532 80726
rect 4580 80778 4636 80780
rect 4580 80726 4582 80778
rect 4582 80726 4634 80778
rect 4634 80726 4636 80778
rect 4580 80724 4636 80726
rect 4684 80778 4740 80780
rect 4684 80726 4686 80778
rect 4686 80726 4738 80778
rect 4738 80726 4740 80778
rect 4684 80724 4740 80726
rect 4476 79210 4532 79212
rect 4476 79158 4478 79210
rect 4478 79158 4530 79210
rect 4530 79158 4532 79210
rect 4476 79156 4532 79158
rect 4580 79210 4636 79212
rect 4580 79158 4582 79210
rect 4582 79158 4634 79210
rect 4634 79158 4636 79210
rect 4580 79156 4636 79158
rect 4684 79210 4740 79212
rect 4684 79158 4686 79210
rect 4686 79158 4738 79210
rect 4738 79158 4740 79210
rect 4684 79156 4740 79158
rect 3612 78428 3668 78484
rect 2156 74226 2212 74228
rect 2156 74174 2158 74226
rect 2158 74174 2210 74226
rect 2210 74174 2212 74226
rect 2156 74172 2212 74174
rect 4476 77642 4532 77644
rect 4476 77590 4478 77642
rect 4478 77590 4530 77642
rect 4530 77590 4532 77642
rect 4476 77588 4532 77590
rect 4580 77642 4636 77644
rect 4580 77590 4582 77642
rect 4582 77590 4634 77642
rect 4634 77590 4636 77642
rect 4580 77588 4636 77590
rect 4684 77642 4740 77644
rect 4684 77590 4686 77642
rect 4686 77590 4738 77642
rect 4738 77590 4740 77642
rect 4684 77588 4740 77590
rect 4476 76074 4532 76076
rect 4476 76022 4478 76074
rect 4478 76022 4530 76074
rect 4530 76022 4532 76074
rect 4476 76020 4532 76022
rect 4580 76074 4636 76076
rect 4580 76022 4582 76074
rect 4582 76022 4634 76074
rect 4634 76022 4636 76074
rect 4580 76020 4636 76022
rect 4684 76074 4740 76076
rect 4684 76022 4686 76074
rect 4686 76022 4738 76074
rect 4738 76022 4740 76074
rect 4684 76020 4740 76022
rect 4844 75740 4900 75796
rect 4284 75628 4340 75684
rect 4172 74732 4228 74788
rect 4396 74786 4452 74788
rect 4396 74734 4398 74786
rect 4398 74734 4450 74786
rect 4450 74734 4452 74786
rect 4396 74732 4452 74734
rect 4844 74620 4900 74676
rect 4476 74506 4532 74508
rect 4476 74454 4478 74506
rect 4478 74454 4530 74506
rect 4530 74454 4532 74506
rect 4476 74452 4532 74454
rect 4580 74506 4636 74508
rect 4580 74454 4582 74506
rect 4582 74454 4634 74506
rect 4634 74454 4636 74506
rect 4580 74452 4636 74454
rect 4684 74506 4740 74508
rect 4684 74454 4686 74506
rect 4686 74454 4738 74506
rect 4738 74454 4740 74506
rect 4684 74452 4740 74454
rect 4172 74060 4228 74116
rect 3724 73948 3780 74004
rect 1708 62188 1764 62244
rect 2940 62188 2996 62244
rect 3388 60508 3444 60564
rect 1820 59164 1876 59220
rect 3052 55356 3108 55412
rect 3388 55916 3444 55972
rect 4476 72938 4532 72940
rect 4476 72886 4478 72938
rect 4478 72886 4530 72938
rect 4530 72886 4532 72938
rect 4476 72884 4532 72886
rect 4580 72938 4636 72940
rect 4580 72886 4582 72938
rect 4582 72886 4634 72938
rect 4634 72886 4636 72938
rect 4580 72884 4636 72886
rect 4684 72938 4740 72940
rect 4684 72886 4686 72938
rect 4686 72886 4738 72938
rect 4738 72886 4740 72938
rect 4684 72884 4740 72886
rect 4476 71370 4532 71372
rect 4476 71318 4478 71370
rect 4478 71318 4530 71370
rect 4530 71318 4532 71370
rect 4476 71316 4532 71318
rect 4580 71370 4636 71372
rect 4580 71318 4582 71370
rect 4582 71318 4634 71370
rect 4634 71318 4636 71370
rect 4580 71316 4636 71318
rect 4684 71370 4740 71372
rect 4684 71318 4686 71370
rect 4686 71318 4738 71370
rect 4738 71318 4740 71370
rect 4684 71316 4740 71318
rect 3836 68460 3892 68516
rect 3612 66332 3668 66388
rect 3724 65996 3780 66052
rect 3164 54684 3220 54740
rect 3836 65212 3892 65268
rect 3948 61628 4004 61684
rect 4476 69802 4532 69804
rect 4476 69750 4478 69802
rect 4478 69750 4530 69802
rect 4530 69750 4532 69802
rect 4476 69748 4532 69750
rect 4580 69802 4636 69804
rect 4580 69750 4582 69802
rect 4582 69750 4634 69802
rect 4634 69750 4636 69802
rect 4580 69748 4636 69750
rect 4684 69802 4740 69804
rect 4684 69750 4686 69802
rect 4686 69750 4738 69802
rect 4738 69750 4740 69802
rect 4684 69748 4740 69750
rect 4508 68626 4564 68628
rect 4508 68574 4510 68626
rect 4510 68574 4562 68626
rect 4562 68574 4564 68626
rect 4508 68572 4564 68574
rect 4476 68234 4532 68236
rect 4476 68182 4478 68234
rect 4478 68182 4530 68234
rect 4530 68182 4532 68234
rect 4476 68180 4532 68182
rect 4580 68234 4636 68236
rect 4580 68182 4582 68234
rect 4582 68182 4634 68234
rect 4634 68182 4636 68234
rect 4580 68180 4636 68182
rect 4684 68234 4740 68236
rect 4684 68182 4686 68234
rect 4686 68182 4738 68234
rect 4738 68182 4740 68234
rect 4684 68180 4740 68182
rect 4476 66666 4532 66668
rect 4476 66614 4478 66666
rect 4478 66614 4530 66666
rect 4530 66614 4532 66666
rect 4476 66612 4532 66614
rect 4580 66666 4636 66668
rect 4580 66614 4582 66666
rect 4582 66614 4634 66666
rect 4634 66614 4636 66666
rect 4580 66612 4636 66614
rect 4684 66666 4740 66668
rect 4684 66614 4686 66666
rect 4686 66614 4738 66666
rect 4738 66614 4740 66666
rect 4684 66612 4740 66614
rect 4396 66332 4452 66388
rect 4284 66050 4340 66052
rect 4284 65998 4286 66050
rect 4286 65998 4338 66050
rect 4338 65998 4340 66050
rect 4284 65996 4340 65998
rect 4508 65212 4564 65268
rect 4476 65098 4532 65100
rect 4476 65046 4478 65098
rect 4478 65046 4530 65098
rect 4530 65046 4532 65098
rect 4476 65044 4532 65046
rect 4580 65098 4636 65100
rect 4580 65046 4582 65098
rect 4582 65046 4634 65098
rect 4634 65046 4636 65098
rect 4580 65044 4636 65046
rect 4684 65098 4740 65100
rect 4684 65046 4686 65098
rect 4686 65046 4738 65098
rect 4738 65046 4740 65098
rect 4684 65044 4740 65046
rect 4172 64540 4228 64596
rect 4844 64594 4900 64596
rect 4844 64542 4846 64594
rect 4846 64542 4898 64594
rect 4898 64542 4900 64594
rect 4844 64540 4900 64542
rect 4620 63756 4676 63812
rect 4476 63530 4532 63532
rect 4476 63478 4478 63530
rect 4478 63478 4530 63530
rect 4530 63478 4532 63530
rect 4476 63476 4532 63478
rect 4580 63530 4636 63532
rect 4580 63478 4582 63530
rect 4582 63478 4634 63530
rect 4634 63478 4636 63530
rect 4580 63476 4636 63478
rect 4684 63530 4740 63532
rect 4684 63478 4686 63530
rect 4686 63478 4738 63530
rect 4738 63478 4740 63530
rect 4684 63476 4740 63478
rect 4172 61346 4228 61348
rect 4172 61294 4174 61346
rect 4174 61294 4226 61346
rect 4226 61294 4228 61346
rect 4172 61292 4228 61294
rect 4476 61962 4532 61964
rect 4476 61910 4478 61962
rect 4478 61910 4530 61962
rect 4530 61910 4532 61962
rect 4476 61908 4532 61910
rect 4580 61962 4636 61964
rect 4580 61910 4582 61962
rect 4582 61910 4634 61962
rect 4634 61910 4636 61962
rect 4580 61908 4636 61910
rect 4684 61962 4740 61964
rect 4684 61910 4686 61962
rect 4686 61910 4738 61962
rect 4738 61910 4740 61962
rect 4684 61908 4740 61910
rect 4284 60844 4340 60900
rect 3724 60562 3780 60564
rect 3724 60510 3726 60562
rect 3726 60510 3778 60562
rect 3778 60510 3780 60562
rect 3724 60508 3780 60510
rect 4396 61628 4452 61684
rect 3612 55410 3668 55412
rect 3612 55358 3614 55410
rect 3614 55358 3666 55410
rect 3666 55358 3668 55410
rect 3612 55356 3668 55358
rect 3500 54908 3556 54964
rect 3612 54738 3668 54740
rect 3612 54686 3614 54738
rect 3614 54686 3666 54738
rect 3666 54686 3668 54738
rect 3612 54684 3668 54686
rect 3836 59052 3892 59108
rect 4508 61292 4564 61348
rect 4508 60562 4564 60564
rect 4508 60510 4510 60562
rect 4510 60510 4562 60562
rect 4562 60510 4564 60562
rect 4508 60508 4564 60510
rect 4476 60394 4532 60396
rect 4476 60342 4478 60394
rect 4478 60342 4530 60394
rect 4530 60342 4532 60394
rect 4476 60340 4532 60342
rect 4580 60394 4636 60396
rect 4580 60342 4582 60394
rect 4582 60342 4634 60394
rect 4634 60342 4636 60394
rect 4580 60340 4636 60342
rect 4684 60394 4740 60396
rect 4684 60342 4686 60394
rect 4686 60342 4738 60394
rect 4738 60342 4740 60394
rect 4684 60340 4740 60342
rect 4844 59948 4900 60004
rect 4620 59724 4676 59780
rect 4476 58826 4532 58828
rect 4476 58774 4478 58826
rect 4478 58774 4530 58826
rect 4530 58774 4532 58826
rect 4476 58772 4532 58774
rect 4580 58826 4636 58828
rect 4580 58774 4582 58826
rect 4582 58774 4634 58826
rect 4634 58774 4636 58826
rect 4580 58772 4636 58774
rect 4684 58826 4740 58828
rect 4684 58774 4686 58826
rect 4686 58774 4738 58826
rect 4738 58774 4740 58826
rect 4684 58772 4740 58774
rect 4620 58210 4676 58212
rect 4620 58158 4622 58210
rect 4622 58158 4674 58210
rect 4674 58158 4676 58210
rect 4620 58156 4676 58158
rect 4476 57258 4532 57260
rect 4476 57206 4478 57258
rect 4478 57206 4530 57258
rect 4530 57206 4532 57258
rect 4476 57204 4532 57206
rect 4580 57258 4636 57260
rect 4580 57206 4582 57258
rect 4582 57206 4634 57258
rect 4634 57206 4636 57258
rect 4580 57204 4636 57206
rect 4684 57258 4740 57260
rect 4684 57206 4686 57258
rect 4686 57206 4738 57258
rect 4738 57206 4740 57258
rect 4684 57204 4740 57206
rect 4476 55690 4532 55692
rect 4476 55638 4478 55690
rect 4478 55638 4530 55690
rect 4530 55638 4532 55690
rect 4476 55636 4532 55638
rect 4580 55690 4636 55692
rect 4580 55638 4582 55690
rect 4582 55638 4634 55690
rect 4634 55638 4636 55690
rect 4580 55636 4636 55638
rect 4684 55690 4740 55692
rect 4684 55638 4686 55690
rect 4686 55638 4738 55690
rect 4738 55638 4740 55690
rect 4684 55636 4740 55638
rect 2044 52162 2100 52164
rect 2044 52110 2046 52162
rect 2046 52110 2098 52162
rect 2098 52110 2100 52162
rect 2044 52108 2100 52110
rect 2716 52050 2772 52052
rect 2716 51998 2718 52050
rect 2718 51998 2770 52050
rect 2770 51998 2772 52050
rect 2716 51996 2772 51998
rect 3500 52668 3556 52724
rect 2940 48300 2996 48356
rect 2268 47068 2324 47124
rect 3276 45612 3332 45668
rect 2268 44322 2324 44324
rect 2268 44270 2270 44322
rect 2270 44270 2322 44322
rect 2322 44270 2324 44322
rect 2268 44268 2324 44270
rect 3164 40348 3220 40404
rect 1932 38668 1988 38724
rect 3276 37772 3332 37828
rect 3724 53618 3780 53620
rect 3724 53566 3726 53618
rect 3726 53566 3778 53618
rect 3778 53566 3780 53618
rect 3724 53564 3780 53566
rect 3948 54402 4004 54404
rect 3948 54350 3950 54402
rect 3950 54350 4002 54402
rect 4002 54350 4004 54402
rect 3948 54348 4004 54350
rect 3948 54012 4004 54068
rect 3836 51996 3892 52052
rect 3724 48354 3780 48356
rect 3724 48302 3726 48354
rect 3726 48302 3778 48354
rect 3778 48302 3780 48354
rect 3724 48300 3780 48302
rect 3612 45666 3668 45668
rect 3612 45614 3614 45666
rect 3614 45614 3666 45666
rect 3666 45614 3668 45666
rect 3612 45612 3668 45614
rect 3500 45052 3556 45108
rect 3612 44322 3668 44324
rect 3612 44270 3614 44322
rect 3614 44270 3666 44322
rect 3666 44270 3668 44322
rect 3612 44268 3668 44270
rect 3612 40460 3668 40516
rect 3612 35644 3668 35700
rect 3724 39340 3780 39396
rect 3164 35196 3220 35252
rect 3612 35196 3668 35252
rect 2492 32396 2548 32452
rect 4620 54402 4676 54404
rect 4620 54350 4622 54402
rect 4622 54350 4674 54402
rect 4674 54350 4676 54402
rect 4620 54348 4676 54350
rect 4476 54122 4532 54124
rect 4476 54070 4478 54122
rect 4478 54070 4530 54122
rect 4530 54070 4532 54122
rect 4476 54068 4532 54070
rect 4580 54122 4636 54124
rect 4580 54070 4582 54122
rect 4582 54070 4634 54122
rect 4634 54070 4636 54122
rect 4580 54068 4636 54070
rect 4684 54122 4740 54124
rect 4684 54070 4686 54122
rect 4686 54070 4738 54122
rect 4738 54070 4740 54122
rect 4684 54068 4740 54070
rect 4844 53842 4900 53844
rect 4844 53790 4846 53842
rect 4846 53790 4898 53842
rect 4898 53790 4900 53842
rect 4844 53788 4900 53790
rect 4060 53004 4116 53060
rect 5628 81228 5684 81284
rect 7084 81394 7140 81396
rect 7084 81342 7086 81394
rect 7086 81342 7138 81394
rect 7138 81342 7140 81394
rect 7084 81340 7140 81342
rect 5964 79436 6020 79492
rect 5964 78876 6020 78932
rect 6860 78764 6916 78820
rect 6524 78706 6580 78708
rect 6524 78654 6526 78706
rect 6526 78654 6578 78706
rect 6578 78654 6580 78706
rect 6524 78652 6580 78654
rect 6076 78428 6132 78484
rect 7084 78876 7140 78932
rect 8988 81340 9044 81396
rect 7420 81116 7476 81172
rect 9660 82908 9716 82964
rect 10220 82850 10276 82852
rect 10220 82798 10222 82850
rect 10222 82798 10274 82850
rect 10274 82798 10276 82850
rect 10220 82796 10276 82798
rect 9772 82572 9828 82628
rect 9660 81842 9716 81844
rect 9660 81790 9662 81842
rect 9662 81790 9714 81842
rect 9714 81790 9716 81842
rect 9660 81788 9716 81790
rect 9884 81394 9940 81396
rect 9884 81342 9886 81394
rect 9886 81342 9938 81394
rect 9938 81342 9940 81394
rect 9884 81340 9940 81342
rect 6860 77420 6916 77476
rect 7308 78540 7364 78596
rect 7308 77420 7364 77476
rect 6972 77308 7028 77364
rect 5964 75964 6020 76020
rect 6860 75852 6916 75908
rect 6300 75682 6356 75684
rect 6300 75630 6302 75682
rect 6302 75630 6354 75682
rect 6354 75630 6356 75682
rect 6300 75628 6356 75630
rect 5292 74284 5348 74340
rect 6524 74786 6580 74788
rect 6524 74734 6526 74786
rect 6526 74734 6578 74786
rect 6578 74734 6580 74786
rect 6524 74732 6580 74734
rect 5852 74002 5908 74004
rect 5852 73950 5854 74002
rect 5854 73950 5906 74002
rect 5906 73950 5908 74002
rect 5852 73948 5908 73950
rect 5740 73836 5796 73892
rect 6188 73836 6244 73892
rect 6748 74060 6804 74116
rect 6636 73836 6692 73892
rect 5068 68796 5124 68852
rect 5292 69132 5348 69188
rect 6748 70028 6804 70084
rect 5964 69132 6020 69188
rect 5516 68908 5572 68964
rect 6076 68908 6132 68964
rect 5068 66946 5124 66948
rect 5068 66894 5070 66946
rect 5070 66894 5122 66946
rect 5122 66894 5124 66946
rect 5068 66892 5124 66894
rect 5068 66386 5124 66388
rect 5068 66334 5070 66386
rect 5070 66334 5122 66386
rect 5122 66334 5124 66386
rect 5068 66332 5124 66334
rect 5292 64428 5348 64484
rect 5068 62242 5124 62244
rect 5068 62190 5070 62242
rect 5070 62190 5122 62242
rect 5122 62190 5124 62242
rect 5068 62188 5124 62190
rect 5628 68572 5684 68628
rect 6636 69186 6692 69188
rect 6636 69134 6638 69186
rect 6638 69134 6690 69186
rect 6690 69134 6692 69186
rect 6636 69132 6692 69134
rect 7084 74396 7140 74452
rect 7308 75964 7364 76020
rect 7308 74844 7364 74900
rect 7196 74338 7252 74340
rect 7196 74286 7198 74338
rect 7198 74286 7250 74338
rect 7250 74286 7252 74338
rect 7196 74284 7252 74286
rect 7196 73948 7252 74004
rect 8988 79436 9044 79492
rect 9772 81170 9828 81172
rect 9772 81118 9774 81170
rect 9774 81118 9826 81170
rect 9826 81118 9828 81170
rect 9772 81116 9828 81118
rect 10668 82460 10724 82516
rect 11004 82460 11060 82516
rect 10444 82348 10500 82404
rect 10220 81282 10276 81284
rect 10220 81230 10222 81282
rect 10222 81230 10274 81282
rect 10274 81230 10276 81282
rect 10220 81228 10276 81230
rect 9996 81004 10052 81060
rect 10892 81842 10948 81844
rect 10892 81790 10894 81842
rect 10894 81790 10946 81842
rect 10946 81790 10948 81842
rect 10892 81788 10948 81790
rect 10780 81340 10836 81396
rect 11564 82348 11620 82404
rect 12012 82348 12068 82404
rect 12684 83244 12740 83300
rect 10668 81058 10724 81060
rect 10668 81006 10670 81058
rect 10670 81006 10722 81058
rect 10722 81006 10724 81058
rect 10668 81004 10724 81006
rect 10556 79602 10612 79604
rect 10556 79550 10558 79602
rect 10558 79550 10610 79602
rect 10610 79550 10612 79602
rect 10556 79548 10612 79550
rect 9660 79490 9716 79492
rect 9660 79438 9662 79490
rect 9662 79438 9714 79490
rect 9714 79438 9716 79490
rect 9660 79436 9716 79438
rect 7532 78818 7588 78820
rect 7532 78766 7534 78818
rect 7534 78766 7586 78818
rect 7586 78766 7588 78818
rect 7532 78764 7588 78766
rect 10668 78876 10724 78932
rect 10220 78594 10276 78596
rect 10220 78542 10222 78594
rect 10222 78542 10274 78594
rect 10274 78542 10276 78594
rect 10220 78540 10276 78542
rect 11564 79548 11620 79604
rect 8316 76524 8372 76580
rect 7644 76412 7700 76468
rect 7644 75794 7700 75796
rect 7644 75742 7646 75794
rect 7646 75742 7698 75794
rect 7698 75742 7700 75794
rect 7644 75740 7700 75742
rect 7756 74898 7812 74900
rect 7756 74846 7758 74898
rect 7758 74846 7810 74898
rect 7810 74846 7812 74898
rect 7756 74844 7812 74846
rect 8092 74786 8148 74788
rect 8092 74734 8094 74786
rect 8094 74734 8146 74786
rect 8146 74734 8148 74786
rect 8092 74732 8148 74734
rect 7868 74396 7924 74452
rect 7420 72268 7476 72324
rect 10108 77250 10164 77252
rect 10108 77198 10110 77250
rect 10110 77198 10162 77250
rect 10162 77198 10164 77250
rect 10108 77196 10164 77198
rect 9548 76524 9604 76580
rect 9772 76466 9828 76468
rect 9772 76414 9774 76466
rect 9774 76414 9826 76466
rect 9826 76414 9828 76466
rect 9772 76412 9828 76414
rect 8764 76188 8820 76244
rect 8316 74956 8372 75012
rect 10220 76466 10276 76468
rect 10220 76414 10222 76466
rect 10222 76414 10274 76466
rect 10274 76414 10276 76466
rect 10220 76412 10276 76414
rect 10332 76300 10388 76356
rect 8764 75010 8820 75012
rect 8764 74958 8766 75010
rect 8766 74958 8818 75010
rect 8818 74958 8820 75010
rect 8764 74956 8820 74958
rect 8428 74844 8484 74900
rect 7980 73948 8036 74004
rect 11116 78204 11172 78260
rect 11340 77868 11396 77924
rect 10668 76354 10724 76356
rect 10668 76302 10670 76354
rect 10670 76302 10722 76354
rect 10722 76302 10724 76354
rect 10668 76300 10724 76302
rect 11116 76354 11172 76356
rect 11116 76302 11118 76354
rect 11118 76302 11170 76354
rect 11170 76302 11172 76354
rect 11116 76300 11172 76302
rect 11564 78818 11620 78820
rect 11564 78766 11566 78818
rect 11566 78766 11618 78818
rect 11618 78766 11620 78818
rect 11564 78764 11620 78766
rect 12460 78818 12516 78820
rect 12460 78766 12462 78818
rect 12462 78766 12514 78818
rect 12514 78766 12516 78818
rect 12460 78764 12516 78766
rect 13692 85036 13748 85092
rect 14028 85260 14084 85316
rect 15820 86604 15876 86660
rect 14588 85090 14644 85092
rect 14588 85038 14590 85090
rect 14590 85038 14642 85090
rect 14642 85038 14644 85090
rect 14588 85036 14644 85038
rect 13804 84866 13860 84868
rect 13804 84814 13806 84866
rect 13806 84814 13858 84866
rect 13858 84814 13860 84866
rect 13804 84812 13860 84814
rect 13692 84140 13748 84196
rect 13916 84476 13972 84532
rect 13804 83356 13860 83412
rect 13692 81340 13748 81396
rect 13468 80892 13524 80948
rect 13468 78540 13524 78596
rect 13580 79548 13636 79604
rect 12908 77922 12964 77924
rect 12908 77870 12910 77922
rect 12910 77870 12962 77922
rect 12962 77870 12964 77922
rect 12908 77868 12964 77870
rect 15148 85314 15204 85316
rect 15148 85262 15150 85314
rect 15150 85262 15202 85314
rect 15202 85262 15204 85314
rect 15148 85260 15204 85262
rect 15596 85090 15652 85092
rect 15596 85038 15598 85090
rect 15598 85038 15650 85090
rect 15650 85038 15652 85090
rect 15596 85036 15652 85038
rect 14140 82908 14196 82964
rect 14028 82460 14084 82516
rect 14812 83020 14868 83076
rect 15260 83298 15316 83300
rect 15260 83246 15262 83298
rect 15262 83246 15314 83298
rect 15314 83246 15316 83298
rect 15260 83244 15316 83246
rect 15148 82460 15204 82516
rect 15372 83132 15428 83188
rect 14476 81394 14532 81396
rect 14476 81342 14478 81394
rect 14478 81342 14530 81394
rect 14530 81342 14532 81394
rect 14476 81340 14532 81342
rect 14028 80892 14084 80948
rect 16044 87612 16100 87668
rect 16716 88284 16772 88340
rect 16716 87612 16772 87668
rect 15596 83410 15652 83412
rect 15596 83358 15598 83410
rect 15598 83358 15650 83410
rect 15650 83358 15652 83410
rect 15596 83356 15652 83358
rect 15484 82236 15540 82292
rect 14924 81340 14980 81396
rect 14140 79602 14196 79604
rect 14140 79550 14142 79602
rect 14142 79550 14194 79602
rect 14194 79550 14196 79602
rect 14140 79548 14196 79550
rect 12908 77308 12964 77364
rect 12348 77138 12404 77140
rect 12348 77086 12350 77138
rect 12350 77086 12402 77138
rect 12402 77086 12404 77138
rect 12348 77084 12404 77086
rect 10892 74620 10948 74676
rect 13468 76300 13524 76356
rect 6188 68796 6244 68852
rect 6188 68236 6244 68292
rect 7084 68908 7140 68964
rect 5852 66892 5908 66948
rect 6524 65436 6580 65492
rect 5740 62636 5796 62692
rect 6860 68124 6916 68180
rect 7084 65436 7140 65492
rect 6748 64764 6804 64820
rect 6188 63644 6244 63700
rect 6972 63756 7028 63812
rect 5740 62188 5796 62244
rect 6748 62636 6804 62692
rect 5964 61682 6020 61684
rect 5964 61630 5966 61682
rect 5966 61630 6018 61682
rect 6018 61630 6020 61682
rect 5964 61628 6020 61630
rect 6524 61682 6580 61684
rect 6524 61630 6526 61682
rect 6526 61630 6578 61682
rect 6578 61630 6580 61682
rect 6524 61628 6580 61630
rect 5740 60898 5796 60900
rect 5740 60846 5742 60898
rect 5742 60846 5794 60898
rect 5794 60846 5796 60898
rect 5740 60844 5796 60846
rect 6188 60786 6244 60788
rect 6188 60734 6190 60786
rect 6190 60734 6242 60786
rect 6242 60734 6244 60786
rect 6188 60732 6244 60734
rect 5292 60508 5348 60564
rect 5852 60002 5908 60004
rect 5852 59950 5854 60002
rect 5854 59950 5906 60002
rect 5906 59950 5908 60002
rect 5852 59948 5908 59950
rect 5740 59836 5796 59892
rect 5628 59778 5684 59780
rect 5628 59726 5630 59778
rect 5630 59726 5682 59778
rect 5682 59726 5684 59778
rect 5628 59724 5684 59726
rect 5404 59052 5460 59108
rect 5068 58268 5124 58324
rect 6860 60898 6916 60900
rect 6860 60846 6862 60898
rect 6862 60846 6914 60898
rect 6914 60846 6916 60898
rect 6860 60844 6916 60846
rect 7532 71820 7588 71876
rect 7644 68124 7700 68180
rect 7532 64482 7588 64484
rect 7532 64430 7534 64482
rect 7534 64430 7586 64482
rect 7586 64430 7588 64482
rect 7532 64428 7588 64430
rect 8092 72268 8148 72324
rect 8540 71874 8596 71876
rect 8540 71822 8542 71874
rect 8542 71822 8594 71874
rect 8594 71822 8596 71874
rect 8540 71820 8596 71822
rect 8764 70082 8820 70084
rect 8764 70030 8766 70082
rect 8766 70030 8818 70082
rect 8818 70030 8820 70082
rect 8764 70028 8820 70030
rect 9548 70812 9604 70868
rect 9996 70812 10052 70868
rect 9548 70028 9604 70084
rect 9884 70082 9940 70084
rect 9884 70030 9886 70082
rect 9886 70030 9938 70082
rect 9938 70030 9940 70082
rect 9884 70028 9940 70030
rect 8204 64428 8260 64484
rect 8428 63308 8484 63364
rect 7644 61346 7700 61348
rect 7644 61294 7646 61346
rect 7646 61294 7698 61346
rect 7698 61294 7700 61346
rect 7644 61292 7700 61294
rect 6188 58268 6244 58324
rect 5740 58210 5796 58212
rect 5740 58158 5742 58210
rect 5742 58158 5794 58210
rect 5794 58158 5796 58210
rect 5740 58156 5796 58158
rect 5852 57148 5908 57204
rect 4956 53228 5012 53284
rect 5068 53788 5124 53844
rect 4620 53116 4676 53172
rect 4844 53004 4900 53060
rect 4476 52554 4532 52556
rect 4476 52502 4478 52554
rect 4478 52502 4530 52554
rect 4530 52502 4532 52554
rect 4476 52500 4532 52502
rect 4580 52554 4636 52556
rect 4580 52502 4582 52554
rect 4582 52502 4634 52554
rect 4634 52502 4636 52554
rect 4580 52500 4636 52502
rect 4684 52554 4740 52556
rect 4684 52502 4686 52554
rect 4686 52502 4738 52554
rect 4738 52502 4740 52554
rect 4684 52500 4740 52502
rect 5404 53170 5460 53172
rect 5404 53118 5406 53170
rect 5406 53118 5458 53170
rect 5458 53118 5460 53170
rect 5404 53116 5460 53118
rect 5180 52946 5236 52948
rect 5180 52894 5182 52946
rect 5182 52894 5234 52946
rect 5234 52894 5236 52946
rect 5180 52892 5236 52894
rect 6188 57148 6244 57204
rect 6188 55020 6244 55076
rect 6188 53788 6244 53844
rect 6300 53564 6356 53620
rect 6076 52892 6132 52948
rect 5068 52108 5124 52164
rect 4956 51996 5012 52052
rect 4172 51378 4228 51380
rect 4172 51326 4174 51378
rect 4174 51326 4226 51378
rect 4226 51326 4228 51378
rect 4172 51324 4228 51326
rect 4476 50986 4532 50988
rect 4476 50934 4478 50986
rect 4478 50934 4530 50986
rect 4530 50934 4532 50986
rect 4476 50932 4532 50934
rect 4580 50986 4636 50988
rect 4580 50934 4582 50986
rect 4582 50934 4634 50986
rect 4634 50934 4636 50986
rect 4580 50932 4636 50934
rect 4684 50986 4740 50988
rect 4684 50934 4686 50986
rect 4686 50934 4738 50986
rect 4738 50934 4740 50986
rect 4684 50932 4740 50934
rect 4732 49532 4788 49588
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 4172 45276 4228 45332
rect 3948 43596 4004 43652
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 3948 40402 4004 40404
rect 3948 40350 3950 40402
rect 3950 40350 4002 40402
rect 4002 40350 4004 40402
rect 3948 40348 4004 40350
rect 5628 51996 5684 52052
rect 5068 50034 5124 50036
rect 5068 49982 5070 50034
rect 5070 49982 5122 50034
rect 5122 49982 5124 50034
rect 5068 49980 5124 49982
rect 4956 49420 5012 49476
rect 5292 48130 5348 48132
rect 5292 48078 5294 48130
rect 5294 48078 5346 48130
rect 5346 48078 5348 48130
rect 5292 48076 5348 48078
rect 5068 47740 5124 47796
rect 5964 49980 6020 50036
rect 4956 45276 5012 45332
rect 5292 47292 5348 47348
rect 5292 47068 5348 47124
rect 4844 44156 4900 44212
rect 4844 43596 4900 43652
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 5516 43538 5572 43540
rect 5516 43486 5518 43538
rect 5518 43486 5570 43538
rect 5570 43486 5572 43538
rect 5516 43484 5572 43486
rect 5740 47234 5796 47236
rect 5740 47182 5742 47234
rect 5742 47182 5794 47234
rect 5794 47182 5796 47234
rect 5740 47180 5796 47182
rect 4844 42700 4900 42756
rect 5068 42754 5124 42756
rect 5068 42702 5070 42754
rect 5070 42702 5122 42754
rect 5122 42702 5124 42754
rect 5068 42700 5124 42702
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 4956 41580 5012 41636
rect 4508 40572 4564 40628
rect 4284 40460 4340 40516
rect 4956 40514 5012 40516
rect 4956 40462 4958 40514
rect 4958 40462 5010 40514
rect 5010 40462 5012 40514
rect 4956 40460 5012 40462
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 5516 42364 5572 42420
rect 5292 41692 5348 41748
rect 4620 39004 4676 39060
rect 5180 39452 5236 39508
rect 5180 38780 5236 38836
rect 3836 37212 3892 37268
rect 3948 37660 4004 37716
rect 4732 38556 4788 38612
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 4844 38162 4900 38164
rect 4844 38110 4846 38162
rect 4846 38110 4898 38162
rect 4898 38110 4900 38162
rect 4844 38108 4900 38110
rect 4284 37826 4340 37828
rect 4284 37774 4286 37826
rect 4286 37774 4338 37826
rect 4338 37774 4340 37826
rect 4284 37772 4340 37774
rect 4620 37772 4676 37828
rect 4172 36652 4228 36708
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4284 36316 4340 36372
rect 4508 36652 4564 36708
rect 4732 35698 4788 35700
rect 4732 35646 4734 35698
rect 4734 35646 4786 35698
rect 4786 35646 4788 35698
rect 4732 35644 4788 35646
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 5068 37772 5124 37828
rect 5180 37212 5236 37268
rect 4620 34018 4676 34020
rect 4620 33966 4622 34018
rect 4622 33966 4674 34018
rect 4674 33966 4676 34018
rect 4620 33964 4676 33966
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 3948 33068 4004 33124
rect 3948 32396 4004 32452
rect 3836 29596 3892 29652
rect 4844 33122 4900 33124
rect 4844 33070 4846 33122
rect 4846 33070 4898 33122
rect 4898 33070 4900 33122
rect 4844 33068 4900 33070
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 5852 42754 5908 42756
rect 5852 42702 5854 42754
rect 5854 42702 5906 42754
rect 5906 42702 5908 42754
rect 5852 42700 5908 42702
rect 5852 42082 5908 42084
rect 5852 42030 5854 42082
rect 5854 42030 5906 42082
rect 5906 42030 5908 42082
rect 5852 42028 5908 42030
rect 6076 47292 6132 47348
rect 6300 51324 6356 51380
rect 6188 46172 6244 46228
rect 6188 43538 6244 43540
rect 6188 43486 6190 43538
rect 6190 43486 6242 43538
rect 6242 43486 6244 43538
rect 6188 43484 6244 43486
rect 6188 42978 6244 42980
rect 6188 42926 6190 42978
rect 6190 42926 6242 42978
rect 6242 42926 6244 42978
rect 6188 42924 6244 42926
rect 6300 42700 6356 42756
rect 6076 41970 6132 41972
rect 6076 41918 6078 41970
rect 6078 41918 6130 41970
rect 6130 41918 6132 41970
rect 6076 41916 6132 41918
rect 5740 40572 5796 40628
rect 5964 40402 6020 40404
rect 5964 40350 5966 40402
rect 5966 40350 6018 40402
rect 6018 40350 6020 40402
rect 5964 40348 6020 40350
rect 5628 40236 5684 40292
rect 5628 39618 5684 39620
rect 5628 39566 5630 39618
rect 5630 39566 5682 39618
rect 5682 39566 5684 39618
rect 5628 39564 5684 39566
rect 5516 39058 5572 39060
rect 5516 39006 5518 39058
rect 5518 39006 5570 39058
rect 5570 39006 5572 39058
rect 5516 39004 5572 39006
rect 5852 39676 5908 39732
rect 5852 39004 5908 39060
rect 6300 41692 6356 41748
rect 6748 58380 6804 58436
rect 7532 60844 7588 60900
rect 6972 58210 7028 58212
rect 6972 58158 6974 58210
rect 6974 58158 7026 58210
rect 7026 58158 7028 58210
rect 6972 58156 7028 58158
rect 7308 59836 7364 59892
rect 7196 59106 7252 59108
rect 7196 59054 7198 59106
rect 7198 59054 7250 59106
rect 7250 59054 7252 59106
rect 7196 59052 7252 59054
rect 7756 60002 7812 60004
rect 7756 59950 7758 60002
rect 7758 59950 7810 60002
rect 7810 59950 7812 60002
rect 7756 59948 7812 59950
rect 7644 58940 7700 58996
rect 7196 58434 7252 58436
rect 7196 58382 7198 58434
rect 7198 58382 7250 58434
rect 7250 58382 7252 58434
rect 7196 58380 7252 58382
rect 7308 58322 7364 58324
rect 7308 58270 7310 58322
rect 7310 58270 7362 58322
rect 7362 58270 7364 58322
rect 7308 58268 7364 58270
rect 6972 57596 7028 57652
rect 6860 54626 6916 54628
rect 6860 54574 6862 54626
rect 6862 54574 6914 54626
rect 6914 54574 6916 54626
rect 6860 54572 6916 54574
rect 6636 53116 6692 53172
rect 6860 52834 6916 52836
rect 6860 52782 6862 52834
rect 6862 52782 6914 52834
rect 6914 52782 6916 52834
rect 6860 52780 6916 52782
rect 7308 53676 7364 53732
rect 7308 53170 7364 53172
rect 7308 53118 7310 53170
rect 7310 53118 7362 53170
rect 7362 53118 7364 53170
rect 7308 53116 7364 53118
rect 7308 52444 7364 52500
rect 7532 57596 7588 57652
rect 7644 52722 7700 52724
rect 7644 52670 7646 52722
rect 7646 52670 7698 52722
rect 7698 52670 7700 52722
rect 7644 52668 7700 52670
rect 7532 52556 7588 52612
rect 7980 61628 8036 61684
rect 8092 60732 8148 60788
rect 7868 58210 7924 58212
rect 7868 58158 7870 58210
rect 7870 58158 7922 58210
rect 7922 58158 7924 58210
rect 7868 58156 7924 58158
rect 6860 48636 6916 48692
rect 6636 42924 6692 42980
rect 6636 42754 6692 42756
rect 6636 42702 6638 42754
rect 6638 42702 6690 42754
rect 6690 42702 6692 42754
rect 6636 42700 6692 42702
rect 7308 41916 7364 41972
rect 7196 41858 7252 41860
rect 7196 41806 7198 41858
rect 7198 41806 7250 41858
rect 7250 41806 7252 41858
rect 7196 41804 7252 41806
rect 6972 41580 7028 41636
rect 7420 41692 7476 41748
rect 6524 40236 6580 40292
rect 6300 39452 6356 39508
rect 6076 39394 6132 39396
rect 6076 39342 6078 39394
rect 6078 39342 6130 39394
rect 6130 39342 6132 39394
rect 6076 39340 6132 39342
rect 5628 38668 5684 38724
rect 5404 38108 5460 38164
rect 5964 38556 6020 38612
rect 3948 29484 4004 29540
rect 4732 30210 4788 30212
rect 4732 30158 4734 30210
rect 4734 30158 4786 30210
rect 4786 30158 4788 30210
rect 4732 30156 4788 30158
rect 5292 30156 5348 30212
rect 4732 29596 4788 29652
rect 4620 29372 4676 29428
rect 2604 25340 2660 25396
rect 3836 26012 3892 26068
rect 4844 29260 4900 29316
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4172 28642 4228 28644
rect 4172 28590 4174 28642
rect 4174 28590 4226 28642
rect 4226 28590 4228 28642
rect 4172 28588 4228 28590
rect 4620 28588 4676 28644
rect 5292 28700 5348 28756
rect 4844 28588 4900 28644
rect 5628 37266 5684 37268
rect 5628 37214 5630 37266
rect 5630 37214 5682 37266
rect 5682 37214 5684 37266
rect 5628 37212 5684 37214
rect 6076 36652 6132 36708
rect 5852 36482 5908 36484
rect 5852 36430 5854 36482
rect 5854 36430 5906 36482
rect 5906 36430 5908 36482
rect 5852 36428 5908 36430
rect 5628 36370 5684 36372
rect 5628 36318 5630 36370
rect 5630 36318 5682 36370
rect 5682 36318 5684 36370
rect 5628 36316 5684 36318
rect 5516 35698 5572 35700
rect 5516 35646 5518 35698
rect 5518 35646 5570 35698
rect 5570 35646 5572 35698
rect 5516 35644 5572 35646
rect 5516 35308 5572 35364
rect 5964 34914 6020 34916
rect 5964 34862 5966 34914
rect 5966 34862 6018 34914
rect 6018 34862 6020 34914
rect 5964 34860 6020 34862
rect 6188 35644 6244 35700
rect 6412 35756 6468 35812
rect 6748 39730 6804 39732
rect 6748 39678 6750 39730
rect 6750 39678 6802 39730
rect 6802 39678 6804 39730
rect 6748 39676 6804 39678
rect 6972 40796 7028 40852
rect 6972 40348 7028 40404
rect 6860 38946 6916 38948
rect 6860 38894 6862 38946
rect 6862 38894 6914 38946
rect 6914 38894 6916 38946
rect 6860 38892 6916 38894
rect 7196 39452 7252 39508
rect 6748 37154 6804 37156
rect 6748 37102 6750 37154
rect 6750 37102 6802 37154
rect 6802 37102 6804 37154
rect 6748 37100 6804 37102
rect 6748 36876 6804 36932
rect 6748 36428 6804 36484
rect 7420 38162 7476 38164
rect 7420 38110 7422 38162
rect 7422 38110 7474 38162
rect 7474 38110 7476 38162
rect 7420 38108 7476 38110
rect 7980 53618 8036 53620
rect 7980 53566 7982 53618
rect 7982 53566 8034 53618
rect 8034 53566 8036 53618
rect 7980 53564 8036 53566
rect 7980 53116 8036 53172
rect 7644 49420 7700 49476
rect 7980 49196 8036 49252
rect 7756 47180 7812 47236
rect 7644 44828 7700 44884
rect 7644 41580 7700 41636
rect 7532 36540 7588 36596
rect 6300 35196 6356 35252
rect 6636 35644 6692 35700
rect 6524 35196 6580 35252
rect 6188 34130 6244 34132
rect 6188 34078 6190 34130
rect 6190 34078 6242 34130
rect 6242 34078 6244 34130
rect 6188 34076 6244 34078
rect 5852 33964 5908 34020
rect 6188 33346 6244 33348
rect 6188 33294 6190 33346
rect 6190 33294 6242 33346
rect 6242 33294 6244 33346
rect 6188 33292 6244 33294
rect 5740 31724 5796 31780
rect 5516 29426 5572 29428
rect 5516 29374 5518 29426
rect 5518 29374 5570 29426
rect 5570 29374 5572 29426
rect 5516 29372 5572 29374
rect 6524 33852 6580 33908
rect 6412 32396 6468 32452
rect 5740 28476 5796 28532
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 4508 26178 4564 26180
rect 4508 26126 4510 26178
rect 4510 26126 4562 26178
rect 4562 26126 4564 26178
rect 4508 26124 4564 26126
rect 5180 26124 5236 26180
rect 4844 26066 4900 26068
rect 4844 26014 4846 26066
rect 4846 26014 4898 26066
rect 4898 26014 4900 26066
rect 4844 26012 4900 26014
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 3948 25452 4004 25508
rect 3724 25394 3780 25396
rect 3724 25342 3726 25394
rect 3726 25342 3778 25394
rect 3778 25342 3780 25394
rect 3724 25340 3780 25342
rect 2604 23884 2660 23940
rect 4284 25228 4340 25284
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 4060 24108 4116 24164
rect 3948 23884 4004 23940
rect 5180 23884 5236 23940
rect 4732 23042 4788 23044
rect 4732 22990 4734 23042
rect 4734 22990 4786 23042
rect 4786 22990 4788 23042
rect 4732 22988 4788 22990
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 5068 22540 5124 22596
rect 4620 22482 4676 22484
rect 4620 22430 4622 22482
rect 4622 22430 4674 22482
rect 4674 22430 4676 22482
rect 4620 22428 4676 22430
rect 1820 22370 1876 22372
rect 1820 22318 1822 22370
rect 1822 22318 1874 22370
rect 1874 22318 1876 22370
rect 1820 22316 1876 22318
rect 4396 21474 4452 21476
rect 4396 21422 4398 21474
rect 4398 21422 4450 21474
rect 4450 21422 4452 21474
rect 4396 21420 4452 21422
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 4172 19458 4228 19460
rect 4172 19406 4174 19458
rect 4174 19406 4226 19458
rect 4226 19406 4228 19458
rect 4172 19404 4228 19406
rect 2604 18284 2660 18340
rect 5068 20802 5124 20804
rect 5068 20750 5070 20802
rect 5070 20750 5122 20802
rect 5122 20750 5124 20802
rect 5068 20748 5124 20750
rect 6076 28476 6132 28532
rect 5628 25282 5684 25284
rect 5628 25230 5630 25282
rect 5630 25230 5682 25282
rect 5682 25230 5684 25282
rect 5628 25228 5684 25230
rect 5628 24162 5684 24164
rect 5628 24110 5630 24162
rect 5630 24110 5682 24162
rect 5682 24110 5684 24162
rect 5628 24108 5684 24110
rect 6748 35196 6804 35252
rect 6748 34188 6804 34244
rect 7196 35644 7252 35700
rect 7084 35308 7140 35364
rect 6972 34354 7028 34356
rect 6972 34302 6974 34354
rect 6974 34302 7026 34354
rect 7026 34302 7028 34354
rect 6972 34300 7028 34302
rect 6860 33852 6916 33908
rect 6972 33346 7028 33348
rect 6972 33294 6974 33346
rect 6974 33294 7026 33346
rect 7026 33294 7028 33346
rect 6972 33292 7028 33294
rect 6748 32450 6804 32452
rect 6748 32398 6750 32450
rect 6750 32398 6802 32450
rect 6802 32398 6804 32450
rect 6748 32396 6804 32398
rect 6300 28642 6356 28644
rect 6300 28590 6302 28642
rect 6302 28590 6354 28642
rect 6354 28590 6356 28642
rect 6300 28588 6356 28590
rect 6188 27916 6244 27972
rect 6636 28530 6692 28532
rect 6636 28478 6638 28530
rect 6638 28478 6690 28530
rect 6690 28478 6692 28530
rect 6636 28476 6692 28478
rect 6636 27916 6692 27972
rect 6524 26908 6580 26964
rect 7196 35196 7252 35252
rect 7420 34860 7476 34916
rect 7196 34076 7252 34132
rect 7308 34188 7364 34244
rect 7756 34130 7812 34132
rect 7756 34078 7758 34130
rect 7758 34078 7810 34130
rect 7810 34078 7812 34130
rect 7756 34076 7812 34078
rect 7420 33964 7476 34020
rect 7420 33068 7476 33124
rect 7308 32620 7364 32676
rect 7084 32450 7140 32452
rect 7084 32398 7086 32450
rect 7086 32398 7138 32450
rect 7138 32398 7140 32450
rect 7084 32396 7140 32398
rect 7756 32620 7812 32676
rect 7308 31778 7364 31780
rect 7308 31726 7310 31778
rect 7310 31726 7362 31778
rect 7362 31726 7364 31778
rect 7308 31724 7364 31726
rect 7756 31164 7812 31220
rect 7308 30156 7364 30212
rect 6972 27804 7028 27860
rect 6972 26908 7028 26964
rect 7084 28588 7140 28644
rect 5964 23938 6020 23940
rect 5964 23886 5966 23938
rect 5966 23886 6018 23938
rect 6018 23886 6020 23938
rect 5964 23884 6020 23886
rect 6188 23938 6244 23940
rect 6188 23886 6190 23938
rect 6190 23886 6242 23938
rect 6242 23886 6244 23938
rect 6188 23884 6244 23886
rect 5852 23324 5908 23380
rect 5404 23154 5460 23156
rect 5404 23102 5406 23154
rect 5406 23102 5458 23154
rect 5458 23102 5460 23154
rect 5404 23100 5460 23102
rect 5292 22988 5348 23044
rect 6300 23154 6356 23156
rect 6300 23102 6302 23154
rect 6302 23102 6354 23154
rect 6354 23102 6356 23154
rect 6300 23100 6356 23102
rect 5628 22428 5684 22484
rect 5852 22540 5908 22596
rect 6748 23548 6804 23604
rect 7308 28588 7364 28644
rect 7308 23548 7364 23604
rect 6748 23378 6804 23380
rect 6748 23326 6750 23378
rect 6750 23326 6802 23378
rect 6802 23326 6804 23378
rect 6748 23324 6804 23326
rect 6860 23100 6916 23156
rect 5852 21420 5908 21476
rect 5964 20802 6020 20804
rect 5964 20750 5966 20802
rect 5966 20750 6018 20802
rect 6018 20750 6020 20802
rect 5964 20748 6020 20750
rect 4956 19404 5012 19460
rect 5068 18508 5124 18564
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 6300 22146 6356 22148
rect 6300 22094 6302 22146
rect 6302 22094 6354 22146
rect 6354 22094 6356 22146
rect 6300 22092 6356 22094
rect 7308 22092 7364 22148
rect 7420 21084 7476 21140
rect 5516 18338 5572 18340
rect 5516 18286 5518 18338
rect 5518 18286 5570 18338
rect 5570 18286 5572 18338
rect 5516 18284 5572 18286
rect 6300 20188 6356 20244
rect 5852 18508 5908 18564
rect 5516 17052 5572 17108
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 7084 15932 7140 15988
rect 6860 15314 6916 15316
rect 6860 15262 6862 15314
rect 6862 15262 6914 15314
rect 6914 15262 6916 15314
rect 6860 15260 6916 15262
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 4732 13746 4788 13748
rect 4732 13694 4734 13746
rect 4734 13694 4786 13746
rect 4786 13694 4788 13746
rect 4732 13692 4788 13694
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 6972 12348 7028 12404
rect 4844 12012 4900 12068
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4732 9938 4788 9940
rect 4732 9886 4734 9938
rect 4734 9886 4786 9938
rect 4786 9886 4788 9938
rect 4732 9884 4788 9886
rect 4284 9212 4340 9268
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 3836 1874 3892 1876
rect 3836 1822 3838 1874
rect 3838 1822 3890 1874
rect 3890 1822 3892 1874
rect 3836 1820 3892 1822
rect 4476 2378 4532 2380
rect 4476 2326 4478 2378
rect 4478 2326 4530 2378
rect 4530 2326 4532 2378
rect 4476 2324 4532 2326
rect 4580 2378 4636 2380
rect 4580 2326 4582 2378
rect 4582 2326 4634 2378
rect 4634 2326 4636 2378
rect 4580 2324 4636 2326
rect 4684 2378 4740 2380
rect 4684 2326 4686 2378
rect 4686 2326 4738 2378
rect 4738 2326 4740 2378
rect 4684 2324 4740 2326
rect 5740 11676 5796 11732
rect 7420 20802 7476 20804
rect 7420 20750 7422 20802
rect 7422 20750 7474 20802
rect 7474 20750 7476 20802
rect 7420 20748 7476 20750
rect 7532 16716 7588 16772
rect 7532 15260 7588 15316
rect 7644 13692 7700 13748
rect 5516 9884 5572 9940
rect 5068 9714 5124 9716
rect 5068 9662 5070 9714
rect 5070 9662 5122 9714
rect 5122 9662 5124 9714
rect 5068 9660 5124 9662
rect 7644 12066 7700 12068
rect 7644 12014 7646 12066
rect 7646 12014 7698 12066
rect 7698 12014 7700 12066
rect 7644 12012 7700 12014
rect 7532 11676 7588 11732
rect 7196 10556 7252 10612
rect 7084 9660 7140 9716
rect 6636 7362 6692 7364
rect 6636 7310 6638 7362
rect 6638 7310 6690 7362
rect 6690 7310 6692 7362
rect 6636 7308 6692 7310
rect 5964 7196 6020 7252
rect 7420 7196 7476 7252
rect 7308 6524 7364 6580
rect 9660 69132 9716 69188
rect 9548 68514 9604 68516
rect 9548 68462 9550 68514
rect 9550 68462 9602 68514
rect 9602 68462 9604 68514
rect 9548 68460 9604 68462
rect 8988 68348 9044 68404
rect 10332 70082 10388 70084
rect 10332 70030 10334 70082
rect 10334 70030 10386 70082
rect 10386 70030 10388 70082
rect 10332 70028 10388 70030
rect 10108 68514 10164 68516
rect 10108 68462 10110 68514
rect 10110 68462 10162 68514
rect 10162 68462 10164 68514
rect 10108 68460 10164 68462
rect 9100 68236 9156 68292
rect 8764 66444 8820 66500
rect 8764 66220 8820 66276
rect 8652 59948 8708 60004
rect 9324 68236 9380 68292
rect 9884 68236 9940 68292
rect 9996 66444 10052 66500
rect 9324 66274 9380 66276
rect 9324 66222 9326 66274
rect 9326 66222 9378 66274
rect 9378 66222 9380 66274
rect 9324 66220 9380 66222
rect 10220 66274 10276 66276
rect 10220 66222 10222 66274
rect 10222 66222 10274 66274
rect 10274 66222 10276 66274
rect 10220 66220 10276 66222
rect 9660 66050 9716 66052
rect 9660 65998 9662 66050
rect 9662 65998 9714 66050
rect 9714 65998 9716 66050
rect 9660 65996 9716 65998
rect 11452 74620 11508 74676
rect 11004 72268 11060 72324
rect 11116 71762 11172 71764
rect 11116 71710 11118 71762
rect 11118 71710 11170 71762
rect 11170 71710 11172 71762
rect 11116 71708 11172 71710
rect 10556 68684 10612 68740
rect 10668 69692 10724 69748
rect 10556 68236 10612 68292
rect 10556 67452 10612 67508
rect 10668 66332 10724 66388
rect 10892 68460 10948 68516
rect 11228 69970 11284 69972
rect 11228 69918 11230 69970
rect 11230 69918 11282 69970
rect 11282 69918 11284 69970
rect 11228 69916 11284 69918
rect 13804 77362 13860 77364
rect 13804 77310 13806 77362
rect 13806 77310 13858 77362
rect 13858 77310 13860 77362
rect 13804 77308 13860 77310
rect 13692 77138 13748 77140
rect 13692 77086 13694 77138
rect 13694 77086 13746 77138
rect 13746 77086 13748 77138
rect 13692 77084 13748 77086
rect 13916 75516 13972 75572
rect 13692 74786 13748 74788
rect 13692 74734 13694 74786
rect 13694 74734 13746 74786
rect 13746 74734 13748 74786
rect 13692 74732 13748 74734
rect 14140 77868 14196 77924
rect 15820 78594 15876 78596
rect 15820 78542 15822 78594
rect 15822 78542 15874 78594
rect 15874 78542 15876 78594
rect 15820 78540 15876 78542
rect 15820 78092 15876 78148
rect 15260 77868 15316 77924
rect 14812 77084 14868 77140
rect 15148 77138 15204 77140
rect 15148 77086 15150 77138
rect 15150 77086 15202 77138
rect 15202 77086 15204 77138
rect 15148 77084 15204 77086
rect 15036 75964 15092 76020
rect 14476 75628 14532 75684
rect 15484 76972 15540 77028
rect 19516 89570 19572 89572
rect 19516 89518 19518 89570
rect 19518 89518 19570 89570
rect 19570 89518 19572 89570
rect 19516 89516 19572 89518
rect 19836 89402 19892 89404
rect 19836 89350 19838 89402
rect 19838 89350 19890 89402
rect 19890 89350 19892 89402
rect 19836 89348 19892 89350
rect 19940 89402 19996 89404
rect 19940 89350 19942 89402
rect 19942 89350 19994 89402
rect 19994 89350 19996 89402
rect 19940 89348 19996 89350
rect 20044 89402 20100 89404
rect 20044 89350 20046 89402
rect 20046 89350 20098 89402
rect 20098 89350 20100 89402
rect 20044 89348 20100 89350
rect 19628 89068 19684 89124
rect 18284 88898 18340 88900
rect 18284 88846 18286 88898
rect 18286 88846 18338 88898
rect 18338 88846 18340 88898
rect 18284 88844 18340 88846
rect 19516 88844 19572 88900
rect 19180 88732 19236 88788
rect 19068 88620 19124 88676
rect 16940 88338 16996 88340
rect 16940 88286 16942 88338
rect 16942 88286 16994 88338
rect 16994 88286 16996 88338
rect 16940 88284 16996 88286
rect 17500 87666 17556 87668
rect 17500 87614 17502 87666
rect 17502 87614 17554 87666
rect 17554 87614 17556 87666
rect 17500 87612 17556 87614
rect 18732 87612 18788 87668
rect 17836 87442 17892 87444
rect 17836 87390 17838 87442
rect 17838 87390 17890 87442
rect 17890 87390 17892 87442
rect 17836 87388 17892 87390
rect 20636 88396 20692 88452
rect 19740 88002 19796 88004
rect 19740 87950 19742 88002
rect 19742 87950 19794 88002
rect 19794 87950 19796 88002
rect 19740 87948 19796 87950
rect 20188 87948 20244 88004
rect 19836 87834 19892 87836
rect 19836 87782 19838 87834
rect 19838 87782 19890 87834
rect 19890 87782 19892 87834
rect 19836 87780 19892 87782
rect 19940 87834 19996 87836
rect 19940 87782 19942 87834
rect 19942 87782 19994 87834
rect 19994 87782 19996 87834
rect 19940 87780 19996 87782
rect 20044 87834 20100 87836
rect 20044 87782 20046 87834
rect 20046 87782 20098 87834
rect 20098 87782 20100 87834
rect 20044 87780 20100 87782
rect 20076 87666 20132 87668
rect 20076 87614 20078 87666
rect 20078 87614 20130 87666
rect 20130 87614 20132 87666
rect 20076 87612 20132 87614
rect 16940 86658 16996 86660
rect 16940 86606 16942 86658
rect 16942 86606 16994 86658
rect 16994 86606 16996 86658
rect 16940 86604 16996 86606
rect 19628 87442 19684 87444
rect 19628 87390 19630 87442
rect 19630 87390 19682 87442
rect 19682 87390 19684 87442
rect 19628 87388 19684 87390
rect 19836 86266 19892 86268
rect 19836 86214 19838 86266
rect 19838 86214 19890 86266
rect 19890 86214 19892 86266
rect 19836 86212 19892 86214
rect 19940 86266 19996 86268
rect 19940 86214 19942 86266
rect 19942 86214 19994 86266
rect 19994 86214 19996 86266
rect 19940 86212 19996 86214
rect 20044 86266 20100 86268
rect 20044 86214 20046 86266
rect 20046 86214 20098 86266
rect 20098 86214 20100 86266
rect 20044 86212 20100 86214
rect 17612 84530 17668 84532
rect 17612 84478 17614 84530
rect 17614 84478 17666 84530
rect 17666 84478 17668 84530
rect 17612 84476 17668 84478
rect 16156 84028 16212 84084
rect 17724 83692 17780 83748
rect 17836 83356 17892 83412
rect 16604 83298 16660 83300
rect 16604 83246 16606 83298
rect 16606 83246 16658 83298
rect 16658 83246 16660 83298
rect 16604 83244 16660 83246
rect 17164 83298 17220 83300
rect 17164 83246 17166 83298
rect 17166 83246 17218 83298
rect 17218 83246 17220 83298
rect 17164 83244 17220 83246
rect 16156 83020 16212 83076
rect 16940 82460 16996 82516
rect 16380 82236 16436 82292
rect 16380 81058 16436 81060
rect 16380 81006 16382 81058
rect 16382 81006 16434 81058
rect 16434 81006 16436 81058
rect 16380 81004 16436 81006
rect 16268 79772 16324 79828
rect 16492 81228 16548 81284
rect 17052 81004 17108 81060
rect 17388 81004 17444 81060
rect 17388 80610 17444 80612
rect 17388 80558 17390 80610
rect 17390 80558 17442 80610
rect 17442 80558 17444 80610
rect 17388 80556 17444 80558
rect 17052 80498 17108 80500
rect 17052 80446 17054 80498
rect 17054 80446 17106 80498
rect 17106 80446 17108 80498
rect 17052 80444 17108 80446
rect 17836 80332 17892 80388
rect 16044 76972 16100 77028
rect 16828 79490 16884 79492
rect 16828 79438 16830 79490
rect 16830 79438 16882 79490
rect 16882 79438 16884 79490
rect 16828 79436 16884 79438
rect 18844 85148 18900 85204
rect 18732 84866 18788 84868
rect 18732 84814 18734 84866
rect 18734 84814 18786 84866
rect 18786 84814 18788 84866
rect 18732 84812 18788 84814
rect 18844 84530 18900 84532
rect 18844 84478 18846 84530
rect 18846 84478 18898 84530
rect 18898 84478 18900 84530
rect 18844 84476 18900 84478
rect 19180 85090 19236 85092
rect 19180 85038 19182 85090
rect 19182 85038 19234 85090
rect 19234 85038 19236 85090
rect 19180 85036 19236 85038
rect 18844 84252 18900 84308
rect 18060 83356 18116 83412
rect 18508 83522 18564 83524
rect 18508 83470 18510 83522
rect 18510 83470 18562 83522
rect 18562 83470 18564 83522
rect 18508 83468 18564 83470
rect 18284 83298 18340 83300
rect 18284 83246 18286 83298
rect 18286 83246 18338 83298
rect 18338 83246 18340 83298
rect 18284 83244 18340 83246
rect 18172 82460 18228 82516
rect 19180 83692 19236 83748
rect 19292 83634 19348 83636
rect 19292 83582 19294 83634
rect 19294 83582 19346 83634
rect 19346 83582 19348 83634
rect 19292 83580 19348 83582
rect 19292 83356 19348 83412
rect 18396 82460 18452 82516
rect 18508 81228 18564 81284
rect 18620 81004 18676 81060
rect 18060 79772 18116 79828
rect 17500 78876 17556 78932
rect 18060 79436 18116 79492
rect 16716 78316 16772 78372
rect 17612 78146 17668 78148
rect 17612 78094 17614 78146
rect 17614 78094 17666 78146
rect 17666 78094 17668 78146
rect 17612 78092 17668 78094
rect 16268 77868 16324 77924
rect 16716 77980 16772 78036
rect 15932 76690 15988 76692
rect 15932 76638 15934 76690
rect 15934 76638 15986 76690
rect 15986 76638 15988 76690
rect 15932 76636 15988 76638
rect 15932 75682 15988 75684
rect 15932 75630 15934 75682
rect 15934 75630 15986 75682
rect 15986 75630 15988 75682
rect 15932 75628 15988 75630
rect 16604 76690 16660 76692
rect 16604 76638 16606 76690
rect 16606 76638 16658 76690
rect 16658 76638 16660 76690
rect 16604 76636 16660 76638
rect 17388 78034 17444 78036
rect 17388 77982 17390 78034
rect 17390 77982 17442 78034
rect 17442 77982 17444 78034
rect 17388 77980 17444 77982
rect 16828 77922 16884 77924
rect 16828 77870 16830 77922
rect 16830 77870 16882 77922
rect 16882 77870 16884 77922
rect 16828 77868 16884 77870
rect 16828 77138 16884 77140
rect 16828 77086 16830 77138
rect 16830 77086 16882 77138
rect 16882 77086 16884 77138
rect 16828 77084 16884 77086
rect 17948 77084 18004 77140
rect 17724 76972 17780 77028
rect 15036 75458 15092 75460
rect 15036 75406 15038 75458
rect 15038 75406 15090 75458
rect 15090 75406 15092 75458
rect 15036 75404 15092 75406
rect 15036 73948 15092 74004
rect 11564 72322 11620 72324
rect 11564 72270 11566 72322
rect 11566 72270 11618 72322
rect 11618 72270 11620 72322
rect 11564 72268 11620 72270
rect 12684 71372 12740 71428
rect 11900 70812 11956 70868
rect 13468 71372 13524 71428
rect 15260 74732 15316 74788
rect 13916 72156 13972 72212
rect 14476 71762 14532 71764
rect 14476 71710 14478 71762
rect 14478 71710 14530 71762
rect 14530 71710 14532 71762
rect 14476 71708 14532 71710
rect 15036 71708 15092 71764
rect 12908 70588 12964 70644
rect 11900 69468 11956 69524
rect 14028 70588 14084 70644
rect 14588 70252 14644 70308
rect 13692 69916 13748 69972
rect 13468 68348 13524 68404
rect 11676 67452 11732 67508
rect 11116 66274 11172 66276
rect 11116 66222 11118 66274
rect 11118 66222 11170 66274
rect 11170 66222 11172 66274
rect 11116 66220 11172 66222
rect 10556 66050 10612 66052
rect 10556 65998 10558 66050
rect 10558 65998 10610 66050
rect 10610 65998 10612 66050
rect 10556 65996 10612 65998
rect 8876 63644 8932 63700
rect 8988 63138 9044 63140
rect 8988 63086 8990 63138
rect 8990 63086 9042 63138
rect 9042 63086 9044 63138
rect 8988 63084 9044 63086
rect 9212 63308 9268 63364
rect 8988 61628 9044 61684
rect 8316 59052 8372 59108
rect 9100 61346 9156 61348
rect 9100 61294 9102 61346
rect 9102 61294 9154 61346
rect 9154 61294 9156 61346
rect 9100 61292 9156 61294
rect 9660 63084 9716 63140
rect 9660 62578 9716 62580
rect 9660 62526 9662 62578
rect 9662 62526 9714 62578
rect 9714 62526 9716 62578
rect 9660 62524 9716 62526
rect 9996 61682 10052 61684
rect 9996 61630 9998 61682
rect 9998 61630 10050 61682
rect 10050 61630 10052 61682
rect 9996 61628 10052 61630
rect 8428 58156 8484 58212
rect 8204 57596 8260 57652
rect 8204 56476 8260 56532
rect 9548 59948 9604 60004
rect 9772 58156 9828 58212
rect 8540 55356 8596 55412
rect 8204 53676 8260 53732
rect 8428 54460 8484 54516
rect 9324 55074 9380 55076
rect 9324 55022 9326 55074
rect 9326 55022 9378 55074
rect 9378 55022 9380 55074
rect 9324 55020 9380 55022
rect 9548 54626 9604 54628
rect 9548 54574 9550 54626
rect 9550 54574 9602 54626
rect 9602 54574 9604 54626
rect 9548 54572 9604 54574
rect 8988 54460 9044 54516
rect 8428 53564 8484 53620
rect 8652 53676 8708 53732
rect 8988 53730 9044 53732
rect 8988 53678 8990 53730
rect 8990 53678 9042 53730
rect 9042 53678 9044 53730
rect 8988 53676 9044 53678
rect 9660 53564 9716 53620
rect 8204 52556 8260 52612
rect 8316 52444 8372 52500
rect 8316 48636 8372 48692
rect 9324 51212 9380 51268
rect 9436 50706 9492 50708
rect 9436 50654 9438 50706
rect 9438 50654 9490 50706
rect 9490 50654 9492 50706
rect 9436 50652 9492 50654
rect 10108 53452 10164 53508
rect 10220 51996 10276 52052
rect 8876 49196 8932 49252
rect 8876 48130 8932 48132
rect 8876 48078 8878 48130
rect 8878 48078 8930 48130
rect 8930 48078 8932 48130
rect 8876 48076 8932 48078
rect 8764 47964 8820 48020
rect 10108 49980 10164 50036
rect 11228 63756 11284 63812
rect 10668 61628 10724 61684
rect 10892 59218 10948 59220
rect 10892 59166 10894 59218
rect 10894 59166 10946 59218
rect 10946 59166 10948 59218
rect 10892 59164 10948 59166
rect 11452 65660 11508 65716
rect 11452 64204 11508 64260
rect 11900 66220 11956 66276
rect 12460 65378 12516 65380
rect 12460 65326 12462 65378
rect 12462 65326 12514 65378
rect 12514 65326 12516 65378
rect 12460 65324 12516 65326
rect 12460 64876 12516 64932
rect 13468 64930 13524 64932
rect 13468 64878 13470 64930
rect 13470 64878 13522 64930
rect 13522 64878 13524 64930
rect 13468 64876 13524 64878
rect 13580 65324 13636 65380
rect 13020 64818 13076 64820
rect 13020 64766 13022 64818
rect 13022 64766 13074 64818
rect 13074 64766 13076 64818
rect 13020 64764 13076 64766
rect 13692 64764 13748 64820
rect 13804 64706 13860 64708
rect 13804 64654 13806 64706
rect 13806 64654 13858 64706
rect 13858 64654 13860 64706
rect 13804 64652 13860 64654
rect 11900 64316 11956 64372
rect 12124 64428 12180 64484
rect 11788 64204 11844 64260
rect 11900 63756 11956 63812
rect 11900 63250 11956 63252
rect 11900 63198 11902 63250
rect 11902 63198 11954 63250
rect 11954 63198 11956 63250
rect 11900 63196 11956 63198
rect 13468 63308 13524 63364
rect 12012 62524 12068 62580
rect 10892 55356 10948 55412
rect 11228 54514 11284 54516
rect 11228 54462 11230 54514
rect 11230 54462 11282 54514
rect 11282 54462 11284 54514
rect 11228 54460 11284 54462
rect 10892 53900 10948 53956
rect 10780 53842 10836 53844
rect 10780 53790 10782 53842
rect 10782 53790 10834 53842
rect 10834 53790 10836 53842
rect 10780 53788 10836 53790
rect 10780 51266 10836 51268
rect 10780 51214 10782 51266
rect 10782 51214 10834 51266
rect 10834 51214 10836 51266
rect 10780 51212 10836 51214
rect 13692 64316 13748 64372
rect 14028 69522 14084 69524
rect 14028 69470 14030 69522
rect 14030 69470 14082 69522
rect 14082 69470 14084 69522
rect 14028 69468 14084 69470
rect 14476 69522 14532 69524
rect 14476 69470 14478 69522
rect 14478 69470 14530 69522
rect 14530 69470 14532 69522
rect 14476 69468 14532 69470
rect 14364 68684 14420 68740
rect 14028 65436 14084 65492
rect 14028 64652 14084 64708
rect 14364 64764 14420 64820
rect 14028 64482 14084 64484
rect 14028 64430 14030 64482
rect 14030 64430 14082 64482
rect 14082 64430 14084 64482
rect 14028 64428 14084 64430
rect 14028 63980 14084 64036
rect 14364 63868 14420 63924
rect 14812 69468 14868 69524
rect 15260 70140 15316 70196
rect 14924 68796 14980 68852
rect 15148 68796 15204 68852
rect 15260 68684 15316 68740
rect 15372 73948 15428 74004
rect 15932 73948 15988 74004
rect 16044 75068 16100 75124
rect 17500 75068 17556 75124
rect 17724 75122 17780 75124
rect 17724 75070 17726 75122
rect 17726 75070 17778 75122
rect 17778 75070 17780 75122
rect 17724 75068 17780 75070
rect 17500 73836 17556 73892
rect 18060 75516 18116 75572
rect 18284 79602 18340 79604
rect 18284 79550 18286 79602
rect 18286 79550 18338 79602
rect 18338 79550 18340 79602
rect 18284 79548 18340 79550
rect 18620 79602 18676 79604
rect 18620 79550 18622 79602
rect 18622 79550 18674 79602
rect 18674 79550 18676 79602
rect 18620 79548 18676 79550
rect 18844 80668 18900 80724
rect 20412 87724 20468 87780
rect 20188 85036 20244 85092
rect 20748 86828 20804 86884
rect 20636 86716 20692 86772
rect 20748 86658 20804 86660
rect 20748 86606 20750 86658
rect 20750 86606 20802 86658
rect 20802 86606 20804 86658
rect 20748 86604 20804 86606
rect 21420 95788 21476 95844
rect 22092 95788 22148 95844
rect 21196 95282 21252 95284
rect 21196 95230 21198 95282
rect 21198 95230 21250 95282
rect 21250 95230 21252 95282
rect 21196 95228 21252 95230
rect 22316 95228 22372 95284
rect 25340 96124 25396 96180
rect 24220 95954 24276 95956
rect 24220 95902 24222 95954
rect 24222 95902 24274 95954
rect 24274 95902 24276 95954
rect 24220 95900 24276 95902
rect 23548 95452 23604 95508
rect 23324 95228 23380 95284
rect 21980 94386 22036 94388
rect 21980 94334 21982 94386
rect 21982 94334 22034 94386
rect 22034 94334 22036 94386
rect 21980 94332 22036 94334
rect 21532 93884 21588 93940
rect 20972 92988 21028 93044
rect 23212 93324 23268 93380
rect 22204 92652 22260 92708
rect 21644 91980 21700 92036
rect 20972 91868 21028 91924
rect 23324 92034 23380 92036
rect 23324 91982 23326 92034
rect 23326 91982 23378 92034
rect 23378 91982 23380 92034
rect 23324 91980 23380 91982
rect 22428 91868 22484 91924
rect 21868 90412 21924 90468
rect 21644 89906 21700 89908
rect 21644 89854 21646 89906
rect 21646 89854 21698 89906
rect 21698 89854 21700 89906
rect 21644 89852 21700 89854
rect 21756 89516 21812 89572
rect 21196 88956 21252 89012
rect 21868 89404 21924 89460
rect 21980 89852 22036 89908
rect 22092 89682 22148 89684
rect 22092 89630 22094 89682
rect 22094 89630 22146 89682
rect 22146 89630 22148 89682
rect 22092 89628 22148 89630
rect 22092 89068 22148 89124
rect 22204 88956 22260 89012
rect 22988 90578 23044 90580
rect 22988 90526 22990 90578
rect 22990 90526 23042 90578
rect 23042 90526 23044 90578
rect 22988 90524 23044 90526
rect 21532 88226 21588 88228
rect 21532 88174 21534 88226
rect 21534 88174 21586 88226
rect 21586 88174 21588 88226
rect 21532 88172 21588 88174
rect 22204 88172 22260 88228
rect 21196 87948 21252 88004
rect 21196 87612 21252 87668
rect 21084 87554 21140 87556
rect 21084 87502 21086 87554
rect 21086 87502 21138 87554
rect 21138 87502 21140 87554
rect 21084 87500 21140 87502
rect 20972 87442 21028 87444
rect 20972 87390 20974 87442
rect 20974 87390 21026 87442
rect 21026 87390 21028 87442
rect 20972 87388 21028 87390
rect 21980 86716 22036 86772
rect 21084 86380 21140 86436
rect 20076 84866 20132 84868
rect 20076 84814 20078 84866
rect 20078 84814 20130 84866
rect 20130 84814 20132 84866
rect 20076 84812 20132 84814
rect 19836 84698 19892 84700
rect 19836 84646 19838 84698
rect 19838 84646 19890 84698
rect 19890 84646 19892 84698
rect 19836 84644 19892 84646
rect 19940 84698 19996 84700
rect 19940 84646 19942 84698
rect 19942 84646 19994 84698
rect 19994 84646 19996 84698
rect 19940 84644 19996 84646
rect 20044 84698 20100 84700
rect 20044 84646 20046 84698
rect 20046 84646 20098 84698
rect 20098 84646 20100 84698
rect 20044 84644 20100 84646
rect 20412 84588 20468 84644
rect 19964 84418 20020 84420
rect 19964 84366 19966 84418
rect 19966 84366 20018 84418
rect 20018 84366 20020 84418
rect 19964 84364 20020 84366
rect 19740 84028 19796 84084
rect 19516 83468 19572 83524
rect 20748 85820 20804 85876
rect 21756 86156 21812 86212
rect 21980 85708 22036 85764
rect 20076 83692 20132 83748
rect 19964 83580 20020 83636
rect 19836 83130 19892 83132
rect 19836 83078 19838 83130
rect 19838 83078 19890 83130
rect 19890 83078 19892 83130
rect 19836 83076 19892 83078
rect 19940 83130 19996 83132
rect 19940 83078 19942 83130
rect 19942 83078 19994 83130
rect 19994 83078 19996 83130
rect 19940 83076 19996 83078
rect 20044 83130 20100 83132
rect 20044 83078 20046 83130
rect 20046 83078 20098 83130
rect 20098 83078 20100 83130
rect 20044 83076 20100 83078
rect 19404 82572 19460 82628
rect 20300 83356 20356 83412
rect 20412 83692 20468 83748
rect 20412 83244 20468 83300
rect 21420 85090 21476 85092
rect 21420 85038 21422 85090
rect 21422 85038 21474 85090
rect 21474 85038 21476 85090
rect 21420 85036 21476 85038
rect 20636 84306 20692 84308
rect 20636 84254 20638 84306
rect 20638 84254 20690 84306
rect 20690 84254 20692 84306
rect 20636 84252 20692 84254
rect 20524 82796 20580 82852
rect 20412 82460 20468 82516
rect 20972 82572 21028 82628
rect 19836 81562 19892 81564
rect 19836 81510 19838 81562
rect 19838 81510 19890 81562
rect 19890 81510 19892 81562
rect 19836 81508 19892 81510
rect 19940 81562 19996 81564
rect 19940 81510 19942 81562
rect 19942 81510 19994 81562
rect 19994 81510 19996 81562
rect 19940 81508 19996 81510
rect 20044 81562 20100 81564
rect 20044 81510 20046 81562
rect 20046 81510 20098 81562
rect 20098 81510 20100 81562
rect 20044 81508 20100 81510
rect 20188 81228 20244 81284
rect 21084 82460 21140 82516
rect 20300 81058 20356 81060
rect 20300 81006 20302 81058
rect 20302 81006 20354 81058
rect 20354 81006 20356 81058
rect 20300 81004 20356 81006
rect 20076 80668 20132 80724
rect 19404 80108 19460 80164
rect 20076 80108 20132 80164
rect 19836 79994 19892 79996
rect 19836 79942 19838 79994
rect 19838 79942 19890 79994
rect 19890 79942 19892 79994
rect 19836 79940 19892 79942
rect 19940 79994 19996 79996
rect 19940 79942 19942 79994
rect 19942 79942 19994 79994
rect 19994 79942 19996 79994
rect 19940 79940 19996 79942
rect 20044 79994 20100 79996
rect 20044 79942 20046 79994
rect 20046 79942 20098 79994
rect 20098 79942 20100 79994
rect 20044 79940 20100 79942
rect 18396 78764 18452 78820
rect 20076 78540 20132 78596
rect 18620 78258 18676 78260
rect 18620 78206 18622 78258
rect 18622 78206 18674 78258
rect 18674 78206 18676 78258
rect 18620 78204 18676 78206
rect 18732 78316 18788 78372
rect 19836 78426 19892 78428
rect 19836 78374 19838 78426
rect 19838 78374 19890 78426
rect 19890 78374 19892 78426
rect 19836 78372 19892 78374
rect 19940 78426 19996 78428
rect 19940 78374 19942 78426
rect 19942 78374 19994 78426
rect 19994 78374 19996 78426
rect 19940 78372 19996 78374
rect 20044 78426 20100 78428
rect 20044 78374 20046 78426
rect 20046 78374 20098 78426
rect 20098 78374 20100 78426
rect 20044 78372 20100 78374
rect 19628 78204 19684 78260
rect 21868 83522 21924 83524
rect 21868 83470 21870 83522
rect 21870 83470 21922 83522
rect 21922 83470 21924 83522
rect 21868 83468 21924 83470
rect 22204 86716 22260 86772
rect 22876 89628 22932 89684
rect 22540 89404 22596 89460
rect 22428 88226 22484 88228
rect 22428 88174 22430 88226
rect 22430 88174 22482 88226
rect 22482 88174 22484 88226
rect 22428 88172 22484 88174
rect 22876 89180 22932 89236
rect 22764 88396 22820 88452
rect 22988 88844 23044 88900
rect 22764 87724 22820 87780
rect 23548 90466 23604 90468
rect 23548 90414 23550 90466
rect 23550 90414 23602 90466
rect 23602 90414 23604 90466
rect 23548 90412 23604 90414
rect 23436 89852 23492 89908
rect 23884 92428 23940 92484
rect 26012 95676 26068 95732
rect 24668 95282 24724 95284
rect 24668 95230 24670 95282
rect 24670 95230 24722 95282
rect 24722 95230 24724 95282
rect 24668 95228 24724 95230
rect 24444 93436 24500 93492
rect 26012 95282 26068 95284
rect 26012 95230 26014 95282
rect 26014 95230 26066 95282
rect 26066 95230 26068 95282
rect 26012 95228 26068 95230
rect 26236 94610 26292 94612
rect 26236 94558 26238 94610
rect 26238 94558 26290 94610
rect 26290 94558 26292 94610
rect 26236 94556 26292 94558
rect 24668 93324 24724 93380
rect 25228 92652 25284 92708
rect 23996 91868 24052 91924
rect 23324 89570 23380 89572
rect 23324 89518 23326 89570
rect 23326 89518 23378 89570
rect 23378 89518 23380 89570
rect 23324 89516 23380 89518
rect 23212 89404 23268 89460
rect 23548 89292 23604 89348
rect 23660 89180 23716 89236
rect 23436 88956 23492 89012
rect 24108 90690 24164 90692
rect 24108 90638 24110 90690
rect 24110 90638 24162 90690
rect 24162 90638 24164 90690
rect 24108 90636 24164 90638
rect 24668 91868 24724 91924
rect 25340 92146 25396 92148
rect 25340 92094 25342 92146
rect 25342 92094 25394 92146
rect 25394 92094 25396 92146
rect 25340 92092 25396 92094
rect 26124 92706 26180 92708
rect 26124 92654 26126 92706
rect 26126 92654 26178 92706
rect 26178 92654 26180 92706
rect 26124 92652 26180 92654
rect 26236 92764 26292 92820
rect 25564 92428 25620 92484
rect 26124 92258 26180 92260
rect 26124 92206 26126 92258
rect 26126 92206 26178 92258
rect 26178 92206 26180 92258
rect 26124 92204 26180 92206
rect 25116 90524 25172 90580
rect 25676 92092 25732 92148
rect 24108 89292 24164 89348
rect 23996 88844 24052 88900
rect 23884 88508 23940 88564
rect 24444 89404 24500 89460
rect 24220 89068 24276 89124
rect 24780 89068 24836 89124
rect 24892 89180 24948 89236
rect 24444 89010 24500 89012
rect 24444 88958 24446 89010
rect 24446 88958 24498 89010
rect 24498 88958 24500 89010
rect 24444 88956 24500 88958
rect 23884 88284 23940 88340
rect 22092 83244 22148 83300
rect 21196 81900 21252 81956
rect 21420 83020 21476 83076
rect 22652 86828 22708 86884
rect 21980 81282 22036 81284
rect 21980 81230 21982 81282
rect 21982 81230 22034 81282
rect 22034 81230 22036 81282
rect 21980 81228 22036 81230
rect 21868 81116 21924 81172
rect 22092 81004 22148 81060
rect 21980 80946 22036 80948
rect 21980 80894 21982 80946
rect 21982 80894 22034 80946
rect 22034 80894 22036 80946
rect 21980 80892 22036 80894
rect 20524 80386 20580 80388
rect 20524 80334 20526 80386
rect 20526 80334 20578 80386
rect 20578 80334 20580 80386
rect 20524 80332 20580 80334
rect 19516 77196 19572 77252
rect 19292 75964 19348 76020
rect 19836 76858 19892 76860
rect 19836 76806 19838 76858
rect 19838 76806 19890 76858
rect 19890 76806 19892 76858
rect 19836 76804 19892 76806
rect 19940 76858 19996 76860
rect 19940 76806 19942 76858
rect 19942 76806 19994 76858
rect 19994 76806 19996 76858
rect 19940 76804 19996 76806
rect 20044 76858 20100 76860
rect 20044 76806 20046 76858
rect 20046 76806 20098 76858
rect 20098 76806 20100 76858
rect 20044 76804 20100 76806
rect 18172 75068 18228 75124
rect 19068 75516 19124 75572
rect 18060 74786 18116 74788
rect 18060 74734 18062 74786
rect 18062 74734 18114 74786
rect 18114 74734 18116 74786
rect 18060 74732 18116 74734
rect 19068 74226 19124 74228
rect 19068 74174 19070 74226
rect 19070 74174 19122 74226
rect 19122 74174 19124 74226
rect 19068 74172 19124 74174
rect 17948 74060 18004 74116
rect 18844 73836 18900 73892
rect 17724 73164 17780 73220
rect 18396 73218 18452 73220
rect 18396 73166 18398 73218
rect 18398 73166 18450 73218
rect 18450 73166 18452 73218
rect 18396 73164 18452 73166
rect 18844 72156 18900 72212
rect 16828 71708 16884 71764
rect 17500 71762 17556 71764
rect 17500 71710 17502 71762
rect 17502 71710 17554 71762
rect 17554 71710 17556 71762
rect 17500 71708 17556 71710
rect 19180 71708 19236 71764
rect 15484 70588 15540 70644
rect 15708 70306 15764 70308
rect 15708 70254 15710 70306
rect 15710 70254 15762 70306
rect 15762 70254 15764 70306
rect 15708 70252 15764 70254
rect 16604 70252 16660 70308
rect 15596 70194 15652 70196
rect 15596 70142 15598 70194
rect 15598 70142 15650 70194
rect 15650 70142 15652 70194
rect 15596 70140 15652 70142
rect 16268 69468 16324 69524
rect 15372 68348 15428 68404
rect 15036 67058 15092 67060
rect 15036 67006 15038 67058
rect 15038 67006 15090 67058
rect 15090 67006 15092 67058
rect 15036 67004 15092 67006
rect 15484 67004 15540 67060
rect 15484 66556 15540 66612
rect 14924 64204 14980 64260
rect 13916 62748 13972 62804
rect 14476 63026 14532 63028
rect 14476 62974 14478 63026
rect 14478 62974 14530 63026
rect 14530 62974 14532 63026
rect 14476 62972 14532 62974
rect 14476 62636 14532 62692
rect 13580 61404 13636 61460
rect 13468 59164 13524 59220
rect 13468 58492 13524 58548
rect 11676 58210 11732 58212
rect 11676 58158 11678 58210
rect 11678 58158 11730 58210
rect 11730 58158 11732 58210
rect 11676 58156 11732 58158
rect 12460 57650 12516 57652
rect 12460 57598 12462 57650
rect 12462 57598 12514 57650
rect 12514 57598 12516 57650
rect 12460 57596 12516 57598
rect 13020 56588 13076 56644
rect 11564 56082 11620 56084
rect 11564 56030 11566 56082
rect 11566 56030 11618 56082
rect 11618 56030 11620 56082
rect 11564 56028 11620 56030
rect 12236 56082 12292 56084
rect 12236 56030 12238 56082
rect 12238 56030 12290 56082
rect 12290 56030 12292 56082
rect 12236 56028 12292 56030
rect 11452 54796 11508 54852
rect 11676 54738 11732 54740
rect 11676 54686 11678 54738
rect 11678 54686 11730 54738
rect 11730 54686 11732 54738
rect 11676 54684 11732 54686
rect 11564 53452 11620 53508
rect 11452 53170 11508 53172
rect 11452 53118 11454 53170
rect 11454 53118 11506 53170
rect 11506 53118 11508 53170
rect 11452 53116 11508 53118
rect 10444 49810 10500 49812
rect 10444 49758 10446 49810
rect 10446 49758 10498 49810
rect 10498 49758 10500 49810
rect 10444 49756 10500 49758
rect 10332 49308 10388 49364
rect 9660 48524 9716 48580
rect 10108 48972 10164 49028
rect 9996 48076 10052 48132
rect 9436 47458 9492 47460
rect 9436 47406 9438 47458
rect 9438 47406 9490 47458
rect 9490 47406 9492 47458
rect 9436 47404 9492 47406
rect 8316 47180 8372 47236
rect 10108 47458 10164 47460
rect 10108 47406 10110 47458
rect 10110 47406 10162 47458
rect 10162 47406 10164 47458
rect 10108 47404 10164 47406
rect 10220 48524 10276 48580
rect 8316 44882 8372 44884
rect 8316 44830 8318 44882
rect 8318 44830 8370 44882
rect 8370 44830 8372 44882
rect 8316 44828 8372 44830
rect 8092 41970 8148 41972
rect 8092 41918 8094 41970
rect 8094 41918 8146 41970
rect 8146 41918 8148 41970
rect 8092 41916 8148 41918
rect 7980 39340 8036 39396
rect 8092 32674 8148 32676
rect 8092 32622 8094 32674
rect 8094 32622 8146 32674
rect 8146 32622 8148 32674
rect 8092 32620 8148 32622
rect 8092 30156 8148 30212
rect 7980 28700 8036 28756
rect 8204 28700 8260 28756
rect 8988 43426 9044 43428
rect 8988 43374 8990 43426
rect 8990 43374 9042 43426
rect 9042 43374 9044 43426
rect 8988 43372 9044 43374
rect 10444 48636 10500 48692
rect 10220 43372 10276 43428
rect 9324 42476 9380 42532
rect 9884 42700 9940 42756
rect 9772 41858 9828 41860
rect 9772 41806 9774 41858
rect 9774 41806 9826 41858
rect 9826 41806 9828 41858
rect 9772 41804 9828 41806
rect 10668 48076 10724 48132
rect 10556 44268 10612 44324
rect 10332 42754 10388 42756
rect 10332 42702 10334 42754
rect 10334 42702 10386 42754
rect 10386 42702 10388 42754
rect 10332 42700 10388 42702
rect 9996 42642 10052 42644
rect 9996 42590 9998 42642
rect 9998 42590 10050 42642
rect 10050 42590 10052 42642
rect 9996 42588 10052 42590
rect 10108 42530 10164 42532
rect 10108 42478 10110 42530
rect 10110 42478 10162 42530
rect 10162 42478 10164 42530
rect 10108 42476 10164 42478
rect 9996 42028 10052 42084
rect 10332 42028 10388 42084
rect 11116 50034 11172 50036
rect 11116 49982 11118 50034
rect 11118 49982 11170 50034
rect 11170 49982 11172 50034
rect 11116 49980 11172 49982
rect 11004 49756 11060 49812
rect 11788 53676 11844 53732
rect 11900 55356 11956 55412
rect 11900 54348 11956 54404
rect 11788 52220 11844 52276
rect 12684 54684 12740 54740
rect 12348 54012 12404 54068
rect 14812 62860 14868 62916
rect 15036 62860 15092 62916
rect 14588 62300 14644 62356
rect 14700 61458 14756 61460
rect 14700 61406 14702 61458
rect 14702 61406 14754 61458
rect 14754 61406 14756 61458
rect 14700 61404 14756 61406
rect 14252 59052 14308 59108
rect 14476 59276 14532 59332
rect 13804 58604 13860 58660
rect 14028 58434 14084 58436
rect 14028 58382 14030 58434
rect 14030 58382 14082 58434
rect 14082 58382 14084 58434
rect 14028 58380 14084 58382
rect 13692 57596 13748 57652
rect 12236 53900 12292 53956
rect 12908 53676 12964 53732
rect 12012 53116 12068 53172
rect 12348 53564 12404 53620
rect 13468 53788 13524 53844
rect 13020 52834 13076 52836
rect 13020 52782 13022 52834
rect 13022 52782 13074 52834
rect 13074 52782 13076 52834
rect 13020 52780 13076 52782
rect 12908 52274 12964 52276
rect 12908 52222 12910 52274
rect 12910 52222 12962 52274
rect 12962 52222 12964 52274
rect 12908 52220 12964 52222
rect 13020 52108 13076 52164
rect 12012 51212 12068 51268
rect 11676 49980 11732 50036
rect 11676 49810 11732 49812
rect 11676 49758 11678 49810
rect 11678 49758 11730 49810
rect 11730 49758 11732 49810
rect 11676 49756 11732 49758
rect 11228 49026 11284 49028
rect 11228 48974 11230 49026
rect 11230 48974 11282 49026
rect 11282 48974 11284 49026
rect 11228 48972 11284 48974
rect 11452 48636 11508 48692
rect 11676 48018 11732 48020
rect 11676 47966 11678 48018
rect 11678 47966 11730 48018
rect 11730 47966 11732 48018
rect 11676 47964 11732 47966
rect 11564 46844 11620 46900
rect 11004 42530 11060 42532
rect 11004 42478 11006 42530
rect 11006 42478 11058 42530
rect 11058 42478 11060 42530
rect 11004 42476 11060 42478
rect 9996 40572 10052 40628
rect 8540 36594 8596 36596
rect 8540 36542 8542 36594
rect 8542 36542 8594 36594
rect 8594 36542 8596 36594
rect 8540 36540 8596 36542
rect 9100 36540 9156 36596
rect 9548 37938 9604 37940
rect 9548 37886 9550 37938
rect 9550 37886 9602 37938
rect 9602 37886 9604 37938
rect 9548 37884 9604 37886
rect 9772 37772 9828 37828
rect 10220 38050 10276 38052
rect 10220 37998 10222 38050
rect 10222 37998 10274 38050
rect 10274 37998 10276 38050
rect 10220 37996 10276 37998
rect 9100 35868 9156 35924
rect 10220 37100 10276 37156
rect 9772 36428 9828 36484
rect 9884 36258 9940 36260
rect 9884 36206 9886 36258
rect 9886 36206 9938 36258
rect 9938 36206 9940 36258
rect 9884 36204 9940 36206
rect 9884 35922 9940 35924
rect 9884 35870 9886 35922
rect 9886 35870 9938 35922
rect 9938 35870 9940 35922
rect 9884 35868 9940 35870
rect 10108 35698 10164 35700
rect 10108 35646 10110 35698
rect 10110 35646 10162 35698
rect 10162 35646 10164 35698
rect 10108 35644 10164 35646
rect 9884 34018 9940 34020
rect 9884 33966 9886 34018
rect 9886 33966 9938 34018
rect 9938 33966 9940 34018
rect 9884 33964 9940 33966
rect 10108 33964 10164 34020
rect 9324 31836 9380 31892
rect 7980 28252 8036 28308
rect 8092 27580 8148 27636
rect 8428 23548 8484 23604
rect 8988 31218 9044 31220
rect 8988 31166 8990 31218
rect 8990 31166 9042 31218
rect 9042 31166 9044 31218
rect 8988 31164 9044 31166
rect 10108 31164 10164 31220
rect 10108 30716 10164 30772
rect 9884 29650 9940 29652
rect 9884 29598 9886 29650
rect 9886 29598 9938 29650
rect 9938 29598 9940 29650
rect 9884 29596 9940 29598
rect 10108 28642 10164 28644
rect 10108 28590 10110 28642
rect 10110 28590 10162 28642
rect 10162 28590 10164 28642
rect 10108 28588 10164 28590
rect 9884 27858 9940 27860
rect 9884 27806 9886 27858
rect 9886 27806 9938 27858
rect 9938 27806 9940 27858
rect 9884 27804 9940 27806
rect 10108 27746 10164 27748
rect 10108 27694 10110 27746
rect 10110 27694 10162 27746
rect 10162 27694 10164 27746
rect 10108 27692 10164 27694
rect 9548 27634 9604 27636
rect 9548 27582 9550 27634
rect 9550 27582 9602 27634
rect 9602 27582 9604 27634
rect 9548 27580 9604 27582
rect 9996 24556 10052 24612
rect 9212 23548 9268 23604
rect 9772 23324 9828 23380
rect 8764 23154 8820 23156
rect 8764 23102 8766 23154
rect 8766 23102 8818 23154
rect 8818 23102 8820 23154
rect 8764 23100 8820 23102
rect 8204 21084 8260 21140
rect 8652 22540 8708 22596
rect 10668 37938 10724 37940
rect 10668 37886 10670 37938
rect 10670 37886 10722 37938
rect 10722 37886 10724 37938
rect 10668 37884 10724 37886
rect 10556 37772 10612 37828
rect 10668 36428 10724 36484
rect 10556 33964 10612 34020
rect 10556 31890 10612 31892
rect 10556 31838 10558 31890
rect 10558 31838 10610 31890
rect 10610 31838 10612 31890
rect 10556 31836 10612 31838
rect 10556 30156 10612 30212
rect 11004 37938 11060 37940
rect 11004 37886 11006 37938
rect 11006 37886 11058 37938
rect 11058 37886 11060 37938
rect 11004 37884 11060 37886
rect 11228 42700 11284 42756
rect 11452 42476 11508 42532
rect 11340 41858 11396 41860
rect 11340 41806 11342 41858
rect 11342 41806 11394 41858
rect 11394 41806 11396 41858
rect 11340 41804 11396 41806
rect 11676 41916 11732 41972
rect 11452 39564 11508 39620
rect 12348 49698 12404 49700
rect 12348 49646 12350 49698
rect 12350 49646 12402 49698
rect 12402 49646 12404 49698
rect 12348 49644 12404 49646
rect 12460 49196 12516 49252
rect 13468 49250 13524 49252
rect 13468 49198 13470 49250
rect 13470 49198 13522 49250
rect 13522 49198 13524 49250
rect 13468 49196 13524 49198
rect 13580 49644 13636 49700
rect 15596 65490 15652 65492
rect 15596 65438 15598 65490
rect 15598 65438 15650 65490
rect 15650 65438 15652 65490
rect 15596 65436 15652 65438
rect 15820 68850 15876 68852
rect 15820 68798 15822 68850
rect 15822 68798 15874 68850
rect 15874 68798 15876 68850
rect 15820 68796 15876 68798
rect 16156 68402 16212 68404
rect 16156 68350 16158 68402
rect 16158 68350 16210 68402
rect 16210 68350 16212 68402
rect 16156 68348 16212 68350
rect 16156 67676 16212 67732
rect 16940 68796 16996 68852
rect 16828 67730 16884 67732
rect 16828 67678 16830 67730
rect 16830 67678 16882 67730
rect 16882 67678 16884 67730
rect 16828 67676 16884 67678
rect 17500 68796 17556 68852
rect 18508 70082 18564 70084
rect 18508 70030 18510 70082
rect 18510 70030 18562 70082
rect 18562 70030 18564 70082
rect 18508 70028 18564 70030
rect 17612 67730 17668 67732
rect 17612 67678 17614 67730
rect 17614 67678 17666 67730
rect 17666 67678 17668 67730
rect 17612 67676 17668 67678
rect 16492 66274 16548 66276
rect 16492 66222 16494 66274
rect 16494 66222 16546 66274
rect 16546 66222 16548 66274
rect 16492 66220 16548 66222
rect 16380 66108 16436 66164
rect 16268 65602 16324 65604
rect 16268 65550 16270 65602
rect 16270 65550 16322 65602
rect 16322 65550 16324 65602
rect 16268 65548 16324 65550
rect 18620 67954 18676 67956
rect 18620 67902 18622 67954
rect 18622 67902 18674 67954
rect 18674 67902 18676 67954
rect 18620 67900 18676 67902
rect 17948 67058 18004 67060
rect 17948 67006 17950 67058
rect 17950 67006 18002 67058
rect 18002 67006 18004 67058
rect 17948 67004 18004 67006
rect 16828 64204 16884 64260
rect 15708 63922 15764 63924
rect 15708 63870 15710 63922
rect 15710 63870 15762 63922
rect 15762 63870 15764 63922
rect 15708 63868 15764 63870
rect 15708 63084 15764 63140
rect 15484 62748 15540 62804
rect 15260 62636 15316 62692
rect 15372 62354 15428 62356
rect 15372 62302 15374 62354
rect 15374 62302 15426 62354
rect 15426 62302 15428 62354
rect 15372 62300 15428 62302
rect 16380 63868 16436 63924
rect 16044 63138 16100 63140
rect 16044 63086 16046 63138
rect 16046 63086 16098 63138
rect 16098 63086 16100 63138
rect 16044 63084 16100 63086
rect 16156 63026 16212 63028
rect 16156 62974 16158 63026
rect 16158 62974 16210 63026
rect 16210 62974 16212 63026
rect 16156 62972 16212 62974
rect 15148 61570 15204 61572
rect 15148 61518 15150 61570
rect 15150 61518 15202 61570
rect 15202 61518 15204 61570
rect 15148 61516 15204 61518
rect 17388 66892 17444 66948
rect 18620 67004 18676 67060
rect 18956 70194 19012 70196
rect 18956 70142 18958 70194
rect 18958 70142 19010 70194
rect 19010 70142 19012 70194
rect 18956 70140 19012 70142
rect 18844 68796 18900 68852
rect 19628 76524 19684 76580
rect 20860 80220 20916 80276
rect 20636 80162 20692 80164
rect 20636 80110 20638 80162
rect 20638 80110 20690 80162
rect 20690 80110 20692 80162
rect 20636 80108 20692 80110
rect 20972 79996 21028 80052
rect 22092 80108 22148 80164
rect 21532 79996 21588 80052
rect 22876 86716 22932 86772
rect 22316 84476 22372 84532
rect 22316 84028 22372 84084
rect 22316 82684 22372 82740
rect 23772 87666 23828 87668
rect 23772 87614 23774 87666
rect 23774 87614 23826 87666
rect 23826 87614 23828 87666
rect 23772 87612 23828 87614
rect 23660 86604 23716 86660
rect 23660 86434 23716 86436
rect 23660 86382 23662 86434
rect 23662 86382 23714 86434
rect 23714 86382 23716 86434
rect 23660 86380 23716 86382
rect 23548 86044 23604 86100
rect 23324 84418 23380 84420
rect 23324 84366 23326 84418
rect 23326 84366 23378 84418
rect 23378 84366 23380 84418
rect 23324 84364 23380 84366
rect 22876 83020 22932 83076
rect 22988 82684 23044 82740
rect 23100 81676 23156 81732
rect 22428 80220 22484 80276
rect 22204 79772 22260 79828
rect 22316 79996 22372 80052
rect 22652 81228 22708 81284
rect 23100 81170 23156 81172
rect 23100 81118 23102 81170
rect 23102 81118 23154 81170
rect 23154 81118 23156 81170
rect 23100 81116 23156 81118
rect 23324 81004 23380 81060
rect 22764 80780 22820 80836
rect 20524 78818 20580 78820
rect 20524 78766 20526 78818
rect 20526 78766 20578 78818
rect 20578 78766 20580 78818
rect 20524 78764 20580 78766
rect 20636 78706 20692 78708
rect 20636 78654 20638 78706
rect 20638 78654 20690 78706
rect 20690 78654 20692 78706
rect 20636 78652 20692 78654
rect 21644 78594 21700 78596
rect 21644 78542 21646 78594
rect 21646 78542 21698 78594
rect 21698 78542 21700 78594
rect 21644 78540 21700 78542
rect 23436 79602 23492 79604
rect 23436 79550 23438 79602
rect 23438 79550 23490 79602
rect 23490 79550 23492 79602
rect 23436 79548 23492 79550
rect 21868 77644 21924 77700
rect 20636 76578 20692 76580
rect 20636 76526 20638 76578
rect 20638 76526 20690 76578
rect 20690 76526 20692 76578
rect 20636 76524 20692 76526
rect 21644 76636 21700 76692
rect 20412 75516 20468 75572
rect 22540 78594 22596 78596
rect 22540 78542 22542 78594
rect 22542 78542 22594 78594
rect 22594 78542 22596 78594
rect 22540 78540 22596 78542
rect 22092 77756 22148 77812
rect 22540 77980 22596 78036
rect 21980 75852 22036 75908
rect 19836 75290 19892 75292
rect 19836 75238 19838 75290
rect 19838 75238 19890 75290
rect 19890 75238 19892 75290
rect 19836 75236 19892 75238
rect 19940 75290 19996 75292
rect 19940 75238 19942 75290
rect 19942 75238 19994 75290
rect 19994 75238 19996 75290
rect 19940 75236 19996 75238
rect 20044 75290 20100 75292
rect 20044 75238 20046 75290
rect 20046 75238 20098 75290
rect 20098 75238 20100 75290
rect 20044 75236 20100 75238
rect 19740 74786 19796 74788
rect 19740 74734 19742 74786
rect 19742 74734 19794 74786
rect 19794 74734 19796 74786
rect 19740 74732 19796 74734
rect 20076 74284 20132 74340
rect 19852 74114 19908 74116
rect 19852 74062 19854 74114
rect 19854 74062 19906 74114
rect 19906 74062 19908 74114
rect 19852 74060 19908 74062
rect 21420 74284 21476 74340
rect 21644 74172 21700 74228
rect 19740 73948 19796 74004
rect 20524 73948 20580 74004
rect 19516 73890 19572 73892
rect 19516 73838 19518 73890
rect 19518 73838 19570 73890
rect 19570 73838 19572 73890
rect 19516 73836 19572 73838
rect 19836 73722 19892 73724
rect 19836 73670 19838 73722
rect 19838 73670 19890 73722
rect 19890 73670 19892 73722
rect 19836 73668 19892 73670
rect 19940 73722 19996 73724
rect 19940 73670 19942 73722
rect 19942 73670 19994 73722
rect 19994 73670 19996 73722
rect 19940 73668 19996 73670
rect 20044 73722 20100 73724
rect 20044 73670 20046 73722
rect 20046 73670 20098 73722
rect 20098 73670 20100 73722
rect 20044 73668 20100 73670
rect 21084 73164 21140 73220
rect 19964 72546 20020 72548
rect 19964 72494 19966 72546
rect 19966 72494 20018 72546
rect 20018 72494 20020 72546
rect 19964 72492 20020 72494
rect 20412 72546 20468 72548
rect 20412 72494 20414 72546
rect 20414 72494 20466 72546
rect 20466 72494 20468 72546
rect 20412 72492 20468 72494
rect 19836 72154 19892 72156
rect 19836 72102 19838 72154
rect 19838 72102 19890 72154
rect 19890 72102 19892 72154
rect 19836 72100 19892 72102
rect 19940 72154 19996 72156
rect 19940 72102 19942 72154
rect 19942 72102 19994 72154
rect 19994 72102 19996 72154
rect 19940 72100 19996 72102
rect 20044 72154 20100 72156
rect 20044 72102 20046 72154
rect 20046 72102 20098 72154
rect 20098 72102 20100 72154
rect 20044 72100 20100 72102
rect 19836 70586 19892 70588
rect 19836 70534 19838 70586
rect 19838 70534 19890 70586
rect 19890 70534 19892 70586
rect 19836 70532 19892 70534
rect 19940 70586 19996 70588
rect 19940 70534 19942 70586
rect 19942 70534 19994 70586
rect 19994 70534 19996 70586
rect 19940 70532 19996 70534
rect 20044 70586 20100 70588
rect 20044 70534 20046 70586
rect 20046 70534 20098 70586
rect 20098 70534 20100 70586
rect 20044 70532 20100 70534
rect 19628 70082 19684 70084
rect 19628 70030 19630 70082
rect 19630 70030 19682 70082
rect 19682 70030 19684 70082
rect 19628 70028 19684 70030
rect 19836 69018 19892 69020
rect 19836 68966 19838 69018
rect 19838 68966 19890 69018
rect 19890 68966 19892 69018
rect 19836 68964 19892 68966
rect 19940 69018 19996 69020
rect 19940 68966 19942 69018
rect 19942 68966 19994 69018
rect 19994 68966 19996 69018
rect 19940 68964 19996 68966
rect 20044 69018 20100 69020
rect 20044 68966 20046 69018
rect 20046 68966 20098 69018
rect 20098 68966 20100 69018
rect 20044 68964 20100 68966
rect 20748 68738 20804 68740
rect 20748 68686 20750 68738
rect 20750 68686 20802 68738
rect 20802 68686 20804 68738
rect 20748 68684 20804 68686
rect 20188 67954 20244 67956
rect 20188 67902 20190 67954
rect 20190 67902 20242 67954
rect 20242 67902 20244 67954
rect 20188 67900 20244 67902
rect 21868 71762 21924 71764
rect 21868 71710 21870 71762
rect 21870 71710 21922 71762
rect 21922 71710 21924 71762
rect 21868 71708 21924 71710
rect 21084 68684 21140 68740
rect 19404 67618 19460 67620
rect 19404 67566 19406 67618
rect 19406 67566 19458 67618
rect 19458 67566 19460 67618
rect 19404 67564 19460 67566
rect 18172 66946 18228 66948
rect 18172 66894 18174 66946
rect 18174 66894 18226 66946
rect 18226 66894 18228 66946
rect 18172 66892 18228 66894
rect 18172 66332 18228 66388
rect 18620 66444 18676 66500
rect 17948 66108 18004 66164
rect 17500 65602 17556 65604
rect 17500 65550 17502 65602
rect 17502 65550 17554 65602
rect 17554 65550 17556 65602
rect 17500 65548 17556 65550
rect 18732 66386 18788 66388
rect 18732 66334 18734 66386
rect 18734 66334 18786 66386
rect 18786 66334 18788 66386
rect 18732 66332 18788 66334
rect 17948 64204 18004 64260
rect 17500 63868 17556 63924
rect 16604 63084 16660 63140
rect 17052 62914 17108 62916
rect 17052 62862 17054 62914
rect 17054 62862 17106 62914
rect 17106 62862 17108 62914
rect 17052 62860 17108 62862
rect 17276 62860 17332 62916
rect 16716 62748 16772 62804
rect 16604 62188 16660 62244
rect 16828 62636 16884 62692
rect 18172 62748 18228 62804
rect 18172 62300 18228 62356
rect 17724 62242 17780 62244
rect 17724 62190 17726 62242
rect 17726 62190 17778 62242
rect 17778 62190 17780 62242
rect 17724 62188 17780 62190
rect 15484 59330 15540 59332
rect 15484 59278 15486 59330
rect 15486 59278 15538 59330
rect 15538 59278 15540 59330
rect 15484 59276 15540 59278
rect 14588 58940 14644 58996
rect 14588 57820 14644 57876
rect 14364 56642 14420 56644
rect 14364 56590 14366 56642
rect 14366 56590 14418 56642
rect 14418 56590 14420 56642
rect 14364 56588 14420 56590
rect 15036 58940 15092 58996
rect 16044 58716 16100 58772
rect 15036 58380 15092 58436
rect 15596 58604 15652 58660
rect 14812 55356 14868 55412
rect 16044 57874 16100 57876
rect 16044 57822 16046 57874
rect 16046 57822 16098 57874
rect 16098 57822 16100 57874
rect 16044 57820 16100 57822
rect 16268 59164 16324 59220
rect 16380 59106 16436 59108
rect 16380 59054 16382 59106
rect 16382 59054 16434 59106
rect 16434 59054 16436 59106
rect 16380 59052 16436 59054
rect 17164 61292 17220 61348
rect 16716 58604 16772 58660
rect 16828 58156 16884 58212
rect 17948 61292 18004 61348
rect 17836 60284 17892 60340
rect 17500 59330 17556 59332
rect 17500 59278 17502 59330
rect 17502 59278 17554 59330
rect 17554 59278 17556 59330
rect 17500 59276 17556 59278
rect 17388 59218 17444 59220
rect 17388 59166 17390 59218
rect 17390 59166 17442 59218
rect 17442 59166 17444 59218
rect 17388 59164 17444 59166
rect 17612 58716 17668 58772
rect 17276 58044 17332 58100
rect 17612 58156 17668 58212
rect 16940 57932 16996 57988
rect 16828 57708 16884 57764
rect 14028 55244 14084 55300
rect 13804 53618 13860 53620
rect 13804 53566 13806 53618
rect 13806 53566 13858 53618
rect 13858 53566 13860 53618
rect 13804 53564 13860 53566
rect 13804 49026 13860 49028
rect 13804 48974 13806 49026
rect 13806 48974 13858 49026
rect 13858 48974 13860 49026
rect 13804 48972 13860 48974
rect 13020 48860 13076 48916
rect 11900 48748 11956 48804
rect 12908 48748 12964 48804
rect 12348 48130 12404 48132
rect 12348 48078 12350 48130
rect 12350 48078 12402 48130
rect 12402 48078 12404 48130
rect 12348 48076 12404 48078
rect 12796 47964 12852 48020
rect 13020 48076 13076 48132
rect 13132 47292 13188 47348
rect 12908 45890 12964 45892
rect 12908 45838 12910 45890
rect 12910 45838 12962 45890
rect 12962 45838 12964 45890
rect 12908 45836 12964 45838
rect 12236 45612 12292 45668
rect 11900 44994 11956 44996
rect 11900 44942 11902 44994
rect 11902 44942 11954 44994
rect 11954 44942 11956 44994
rect 11900 44940 11956 44942
rect 12460 44994 12516 44996
rect 12460 44942 12462 44994
rect 12462 44942 12514 44994
rect 12514 44942 12516 44994
rect 12460 44940 12516 44942
rect 13916 48466 13972 48468
rect 13916 48414 13918 48466
rect 13918 48414 13970 48466
rect 13970 48414 13972 48466
rect 13916 48412 13972 48414
rect 13692 47516 13748 47572
rect 13580 47234 13636 47236
rect 13580 47182 13582 47234
rect 13582 47182 13634 47234
rect 13634 47182 13636 47234
rect 13580 47180 13636 47182
rect 14252 53506 14308 53508
rect 14252 53454 14254 53506
rect 14254 53454 14306 53506
rect 14306 53454 14308 53506
rect 14252 53452 14308 53454
rect 14812 54012 14868 54068
rect 14364 49756 14420 49812
rect 15596 54012 15652 54068
rect 15820 53730 15876 53732
rect 15820 53678 15822 53730
rect 15822 53678 15874 53730
rect 15874 53678 15876 53730
rect 15820 53676 15876 53678
rect 15260 53116 15316 53172
rect 16044 52892 16100 52948
rect 15596 52162 15652 52164
rect 15596 52110 15598 52162
rect 15598 52110 15650 52162
rect 15650 52110 15652 52162
rect 15596 52108 15652 52110
rect 15820 51660 15876 51716
rect 14140 48914 14196 48916
rect 14140 48862 14142 48914
rect 14142 48862 14194 48914
rect 14194 48862 14196 48914
rect 14140 48860 14196 48862
rect 14252 48802 14308 48804
rect 14252 48750 14254 48802
rect 14254 48750 14306 48802
rect 14306 48750 14308 48802
rect 14252 48748 14308 48750
rect 14476 49196 14532 49252
rect 14364 47180 14420 47236
rect 13804 45890 13860 45892
rect 13804 45838 13806 45890
rect 13806 45838 13858 45890
rect 13858 45838 13860 45890
rect 13804 45836 13860 45838
rect 12460 39394 12516 39396
rect 12460 39342 12462 39394
rect 12462 39342 12514 39394
rect 12514 39342 12516 39394
rect 12460 39340 12516 39342
rect 11452 38050 11508 38052
rect 11452 37998 11454 38050
rect 11454 37998 11506 38050
rect 11506 37998 11508 38050
rect 11452 37996 11508 37998
rect 11676 37154 11732 37156
rect 11676 37102 11678 37154
rect 11678 37102 11730 37154
rect 11730 37102 11732 37154
rect 11676 37100 11732 37102
rect 12012 36540 12068 36596
rect 11116 35698 11172 35700
rect 11116 35646 11118 35698
rect 11118 35646 11170 35698
rect 11170 35646 11172 35698
rect 11116 35644 11172 35646
rect 11564 33964 11620 34020
rect 11676 33516 11732 33572
rect 11004 30156 11060 30212
rect 10556 29596 10612 29652
rect 10556 27858 10612 27860
rect 10556 27806 10558 27858
rect 10558 27806 10610 27858
rect 10610 27806 10612 27858
rect 10556 27804 10612 27806
rect 10332 24610 10388 24612
rect 10332 24558 10334 24610
rect 10334 24558 10386 24610
rect 10386 24558 10388 24610
rect 10332 24556 10388 24558
rect 9772 22540 9828 22596
rect 8092 20188 8148 20244
rect 8652 20188 8708 20244
rect 9324 18396 9380 18452
rect 7980 15932 8036 15988
rect 8652 17106 8708 17108
rect 8652 17054 8654 17106
rect 8654 17054 8706 17106
rect 8706 17054 8708 17106
rect 8652 17052 8708 17054
rect 10220 18396 10276 18452
rect 10556 23378 10612 23380
rect 10556 23326 10558 23378
rect 10558 23326 10610 23378
rect 10610 23326 10612 23378
rect 10556 23324 10612 23326
rect 10780 29538 10836 29540
rect 10780 29486 10782 29538
rect 10782 29486 10834 29538
rect 10834 29486 10836 29538
rect 10780 29484 10836 29486
rect 11340 29484 11396 29540
rect 12236 37100 12292 37156
rect 12236 33852 12292 33908
rect 12236 31612 12292 31668
rect 11004 23100 11060 23156
rect 11452 22482 11508 22484
rect 11452 22430 11454 22482
rect 11454 22430 11506 22482
rect 11506 22430 11508 22482
rect 11452 22428 11508 22430
rect 11004 22092 11060 22148
rect 10892 21586 10948 21588
rect 10892 21534 10894 21586
rect 10894 21534 10946 21586
rect 10946 21534 10948 21586
rect 10892 21532 10948 21534
rect 10220 16156 10276 16212
rect 8092 15484 8148 15540
rect 8988 15538 9044 15540
rect 8988 15486 8990 15538
rect 8990 15486 9042 15538
rect 9042 15486 9044 15538
rect 8988 15484 9044 15486
rect 10220 15484 10276 15540
rect 8316 13804 8372 13860
rect 7980 13746 8036 13748
rect 7980 13694 7982 13746
rect 7982 13694 8034 13746
rect 8034 13694 8036 13746
rect 7980 13692 8036 13694
rect 9548 13858 9604 13860
rect 9548 13806 9550 13858
rect 9550 13806 9602 13858
rect 9602 13806 9604 13858
rect 9548 13804 9604 13806
rect 8092 12402 8148 12404
rect 8092 12350 8094 12402
rect 8094 12350 8146 12402
rect 8146 12350 8148 12402
rect 8092 12348 8148 12350
rect 9884 12348 9940 12404
rect 8428 12012 8484 12068
rect 8988 12066 9044 12068
rect 8988 12014 8990 12066
rect 8990 12014 9042 12066
rect 9042 12014 9044 12066
rect 8988 12012 9044 12014
rect 8988 11676 9044 11732
rect 8540 10332 8596 10388
rect 9996 10332 10052 10388
rect 10108 10668 10164 10724
rect 8988 9266 9044 9268
rect 8988 9214 8990 9266
rect 8990 9214 9042 9266
rect 9042 9214 9044 9266
rect 8988 9212 9044 9214
rect 9884 9212 9940 9268
rect 10220 10610 10276 10612
rect 10220 10558 10222 10610
rect 10222 10558 10274 10610
rect 10274 10558 10276 10610
rect 10220 10556 10276 10558
rect 8652 7196 8708 7252
rect 5292 5180 5348 5236
rect 6412 5180 6468 5236
rect 5628 4844 5684 4900
rect 5852 1874 5908 1876
rect 5852 1822 5854 1874
rect 5854 1822 5906 1874
rect 5906 1822 5908 1874
rect 5852 1820 5908 1822
rect 5068 1762 5124 1764
rect 5068 1710 5070 1762
rect 5070 1710 5122 1762
rect 5122 1710 5124 1762
rect 5068 1708 5124 1710
rect 6300 3442 6356 3444
rect 6300 3390 6302 3442
rect 6302 3390 6354 3442
rect 6354 3390 6356 3442
rect 6300 3388 6356 3390
rect 8652 5516 8708 5572
rect 8988 7084 9044 7140
rect 8092 4508 8148 4564
rect 8204 4060 8260 4116
rect 7532 3500 7588 3556
rect 7420 3442 7476 3444
rect 7420 3390 7422 3442
rect 7422 3390 7474 3442
rect 7474 3390 7476 3442
rect 7420 3388 7476 3390
rect 10108 6802 10164 6804
rect 10108 6750 10110 6802
rect 10110 6750 10162 6802
rect 10162 6750 10164 6802
rect 10108 6748 10164 6750
rect 9996 6636 10052 6692
rect 9660 6524 9716 6580
rect 10444 15314 10500 15316
rect 10444 15262 10446 15314
rect 10446 15262 10498 15314
rect 10498 15262 10500 15314
rect 10444 15260 10500 15262
rect 11116 20188 11172 20244
rect 11116 19740 11172 19796
rect 11788 19794 11844 19796
rect 11788 19742 11790 19794
rect 11790 19742 11842 19794
rect 11842 19742 11844 19794
rect 11788 19740 11844 19742
rect 11788 17500 11844 17556
rect 10780 17052 10836 17108
rect 11452 15820 11508 15876
rect 11452 15260 11508 15316
rect 12124 22988 12180 23044
rect 12012 20860 12068 20916
rect 12124 19740 12180 19796
rect 12572 37266 12628 37268
rect 12572 37214 12574 37266
rect 12574 37214 12626 37266
rect 12626 37214 12628 37266
rect 12572 37212 12628 37214
rect 13244 41916 13300 41972
rect 12908 41298 12964 41300
rect 12908 41246 12910 41298
rect 12910 41246 12962 41298
rect 12962 41246 12964 41298
rect 12908 41244 12964 41246
rect 13020 40572 13076 40628
rect 12908 39618 12964 39620
rect 12908 39566 12910 39618
rect 12910 39566 12962 39618
rect 12962 39566 12964 39618
rect 12908 39564 12964 39566
rect 13580 40514 13636 40516
rect 13580 40462 13582 40514
rect 13582 40462 13634 40514
rect 13634 40462 13636 40514
rect 13580 40460 13636 40462
rect 13692 40572 13748 40628
rect 13804 40460 13860 40516
rect 13356 38108 13412 38164
rect 12684 36988 12740 37044
rect 13020 37154 13076 37156
rect 13020 37102 13022 37154
rect 13022 37102 13074 37154
rect 13074 37102 13076 37154
rect 13020 37100 13076 37102
rect 12908 35644 12964 35700
rect 12684 33852 12740 33908
rect 13580 33516 13636 33572
rect 13580 32508 13636 32564
rect 12684 28812 12740 28868
rect 13244 29596 13300 29652
rect 12908 28140 12964 28196
rect 13468 28866 13524 28868
rect 13468 28814 13470 28866
rect 13470 28814 13522 28866
rect 13522 28814 13524 28866
rect 13468 28812 13524 28814
rect 13580 28588 13636 28644
rect 13468 27692 13524 27748
rect 12684 25394 12740 25396
rect 12684 25342 12686 25394
rect 12686 25342 12738 25394
rect 12738 25342 12740 25394
rect 12684 25340 12740 25342
rect 13244 25340 13300 25396
rect 13020 25116 13076 25172
rect 12796 24162 12852 24164
rect 12796 24110 12798 24162
rect 12798 24110 12850 24162
rect 12850 24110 12852 24162
rect 12796 24108 12852 24110
rect 12348 23548 12404 23604
rect 12684 23548 12740 23604
rect 12348 23042 12404 23044
rect 12348 22990 12350 23042
rect 12350 22990 12402 23042
rect 12402 22990 12404 23042
rect 12348 22988 12404 22990
rect 12348 22482 12404 22484
rect 12348 22430 12350 22482
rect 12350 22430 12402 22482
rect 12402 22430 12404 22482
rect 12348 22428 12404 22430
rect 12796 22540 12852 22596
rect 14028 45106 14084 45108
rect 14028 45054 14030 45106
rect 14030 45054 14082 45106
rect 14082 45054 14084 45106
rect 14028 45052 14084 45054
rect 14364 45330 14420 45332
rect 14364 45278 14366 45330
rect 14366 45278 14418 45330
rect 14418 45278 14420 45330
rect 14364 45276 14420 45278
rect 15372 50482 15428 50484
rect 15372 50430 15374 50482
rect 15374 50430 15426 50482
rect 15426 50430 15428 50482
rect 15372 50428 15428 50430
rect 14924 49756 14980 49812
rect 14812 49196 14868 49252
rect 15260 49532 15316 49588
rect 14700 48972 14756 49028
rect 14924 48802 14980 48804
rect 14924 48750 14926 48802
rect 14926 48750 14978 48802
rect 14978 48750 14980 48802
rect 14924 48748 14980 48750
rect 14700 48188 14756 48244
rect 14812 47740 14868 47796
rect 15372 48242 15428 48244
rect 15372 48190 15374 48242
rect 15374 48190 15426 48242
rect 15426 48190 15428 48242
rect 15372 48188 15428 48190
rect 17388 57762 17444 57764
rect 17388 57710 17390 57762
rect 17390 57710 17442 57762
rect 17442 57710 17444 57762
rect 17388 57708 17444 57710
rect 16604 56476 16660 56532
rect 17164 56476 17220 56532
rect 16716 55020 16772 55076
rect 16268 53170 16324 53172
rect 16268 53118 16270 53170
rect 16270 53118 16322 53170
rect 16322 53118 16324 53170
rect 16268 53116 16324 53118
rect 16268 52668 16324 52724
rect 16604 53058 16660 53060
rect 16604 53006 16606 53058
rect 16606 53006 16658 53058
rect 16658 53006 16660 53058
rect 16604 53004 16660 53006
rect 16380 52556 16436 52612
rect 16604 51548 16660 51604
rect 16380 51378 16436 51380
rect 16380 51326 16382 51378
rect 16382 51326 16434 51378
rect 16434 51326 16436 51378
rect 16380 51324 16436 51326
rect 16268 50876 16324 50932
rect 15932 50370 15988 50372
rect 15932 50318 15934 50370
rect 15934 50318 15986 50370
rect 15986 50318 15988 50370
rect 15932 50316 15988 50318
rect 15596 49308 15652 49364
rect 17836 58604 17892 58660
rect 17836 58044 17892 58100
rect 18172 59164 18228 59220
rect 17948 56978 18004 56980
rect 17948 56926 17950 56978
rect 17950 56926 18002 56978
rect 18002 56926 18004 56978
rect 17948 56924 18004 56926
rect 18620 64428 18676 64484
rect 18620 62578 18676 62580
rect 18620 62526 18622 62578
rect 18622 62526 18674 62578
rect 18674 62526 18676 62578
rect 18620 62524 18676 62526
rect 18956 67004 19012 67060
rect 18732 62076 18788 62132
rect 18732 60620 18788 60676
rect 18844 65772 18900 65828
rect 19180 66498 19236 66500
rect 19180 66446 19182 66498
rect 19182 66446 19234 66498
rect 19234 66446 19236 66498
rect 19180 66444 19236 66446
rect 19404 66444 19460 66500
rect 19292 66220 19348 66276
rect 19836 67450 19892 67452
rect 19836 67398 19838 67450
rect 19838 67398 19890 67450
rect 19890 67398 19892 67450
rect 19836 67396 19892 67398
rect 19940 67450 19996 67452
rect 19940 67398 19942 67450
rect 19942 67398 19994 67450
rect 19994 67398 19996 67450
rect 19940 67396 19996 67398
rect 20044 67450 20100 67452
rect 20044 67398 20046 67450
rect 20046 67398 20098 67450
rect 20098 67398 20100 67450
rect 20044 67396 20100 67398
rect 20076 67116 20132 67172
rect 20412 66274 20468 66276
rect 20412 66222 20414 66274
rect 20414 66222 20466 66274
rect 20466 66222 20468 66274
rect 20412 66220 20468 66222
rect 18956 63084 19012 63140
rect 18956 62524 19012 62580
rect 19836 65882 19892 65884
rect 19836 65830 19838 65882
rect 19838 65830 19890 65882
rect 19890 65830 19892 65882
rect 19836 65828 19892 65830
rect 19940 65882 19996 65884
rect 19940 65830 19942 65882
rect 19942 65830 19994 65882
rect 19994 65830 19996 65882
rect 19940 65828 19996 65830
rect 20044 65882 20100 65884
rect 20044 65830 20046 65882
rect 20046 65830 20098 65882
rect 20098 65830 20100 65882
rect 20044 65828 20100 65830
rect 19404 65324 19460 65380
rect 19516 65660 19572 65716
rect 19836 64314 19892 64316
rect 19836 64262 19838 64314
rect 19838 64262 19890 64314
rect 19890 64262 19892 64314
rect 19836 64260 19892 64262
rect 19940 64314 19996 64316
rect 19940 64262 19942 64314
rect 19942 64262 19994 64314
rect 19994 64262 19996 64314
rect 19940 64260 19996 64262
rect 20044 64314 20100 64316
rect 20044 64262 20046 64314
rect 20046 64262 20098 64314
rect 20098 64262 20100 64314
rect 20044 64260 20100 64262
rect 19964 64034 20020 64036
rect 19964 63982 19966 64034
rect 19966 63982 20018 64034
rect 20018 63982 20020 64034
rect 19964 63980 20020 63982
rect 19404 62524 19460 62580
rect 18956 61516 19012 61572
rect 18956 61010 19012 61012
rect 18956 60958 18958 61010
rect 18958 60958 19010 61010
rect 19010 60958 19012 61010
rect 18956 60956 19012 60958
rect 18956 60732 19012 60788
rect 18732 59442 18788 59444
rect 18732 59390 18734 59442
rect 18734 59390 18786 59442
rect 18786 59390 18788 59442
rect 18732 59388 18788 59390
rect 18620 58604 18676 58660
rect 18508 57372 18564 57428
rect 18060 56364 18116 56420
rect 18284 57148 18340 57204
rect 18396 56924 18452 56980
rect 17948 55916 18004 55972
rect 17052 53842 17108 53844
rect 17052 53790 17054 53842
rect 17054 53790 17106 53842
rect 17106 53790 17108 53842
rect 17052 53788 17108 53790
rect 16828 53676 16884 53732
rect 16828 52274 16884 52276
rect 16828 52222 16830 52274
rect 16830 52222 16882 52274
rect 16882 52222 16884 52274
rect 16828 52220 16884 52222
rect 17164 52220 17220 52276
rect 16828 51996 16884 52052
rect 16716 50988 16772 51044
rect 16492 49308 16548 49364
rect 15932 48972 15988 49028
rect 16044 49084 16100 49140
rect 15820 48802 15876 48804
rect 15820 48750 15822 48802
rect 15822 48750 15874 48802
rect 15874 48750 15876 48802
rect 15820 48748 15876 48750
rect 15596 47516 15652 47572
rect 16268 48524 16324 48580
rect 15820 48300 15876 48356
rect 15820 47740 15876 47796
rect 15036 47346 15092 47348
rect 15036 47294 15038 47346
rect 15038 47294 15090 47346
rect 15090 47294 15092 47346
rect 15036 47292 15092 47294
rect 15484 47346 15540 47348
rect 15484 47294 15486 47346
rect 15486 47294 15538 47346
rect 15538 47294 15540 47346
rect 15484 47292 15540 47294
rect 15708 47180 15764 47236
rect 16492 48300 16548 48356
rect 16268 47234 16324 47236
rect 16268 47182 16270 47234
rect 16270 47182 16322 47234
rect 16322 47182 16324 47234
rect 16268 47180 16324 47182
rect 14364 42252 14420 42308
rect 14364 40514 14420 40516
rect 14364 40462 14366 40514
rect 14366 40462 14418 40514
rect 14418 40462 14420 40514
rect 14364 40460 14420 40462
rect 14028 39394 14084 39396
rect 14028 39342 14030 39394
rect 14030 39342 14082 39394
rect 14082 39342 14084 39394
rect 14028 39340 14084 39342
rect 15596 46562 15652 46564
rect 15596 46510 15598 46562
rect 15598 46510 15650 46562
rect 15650 46510 15652 46562
rect 15596 46508 15652 46510
rect 16268 46508 16324 46564
rect 15932 46284 15988 46340
rect 15148 45276 15204 45332
rect 15372 45106 15428 45108
rect 15372 45054 15374 45106
rect 15374 45054 15426 45106
rect 15426 45054 15428 45106
rect 15372 45052 15428 45054
rect 15260 44156 15316 44212
rect 15148 43596 15204 43652
rect 15596 44098 15652 44100
rect 15596 44046 15598 44098
rect 15598 44046 15650 44098
rect 15650 44046 15652 44098
rect 15596 44044 15652 44046
rect 15372 43148 15428 43204
rect 15484 43260 15540 43316
rect 15036 42588 15092 42644
rect 14812 42140 14868 42196
rect 14588 41916 14644 41972
rect 15036 41858 15092 41860
rect 15036 41806 15038 41858
rect 15038 41806 15090 41858
rect 15090 41806 15092 41858
rect 15036 41804 15092 41806
rect 15148 41244 15204 41300
rect 14812 41186 14868 41188
rect 14812 41134 14814 41186
rect 14814 41134 14866 41186
rect 14866 41134 14868 41186
rect 14812 41132 14868 41134
rect 14924 40236 14980 40292
rect 15148 39618 15204 39620
rect 15148 39566 15150 39618
rect 15150 39566 15202 39618
rect 15202 39566 15204 39618
rect 15148 39564 15204 39566
rect 14924 39394 14980 39396
rect 14924 39342 14926 39394
rect 14926 39342 14978 39394
rect 14978 39342 14980 39394
rect 14924 39340 14980 39342
rect 15036 39228 15092 39284
rect 13916 37826 13972 37828
rect 13916 37774 13918 37826
rect 13918 37774 13970 37826
rect 13970 37774 13972 37826
rect 13916 37772 13972 37774
rect 13804 30380 13860 30436
rect 13804 29596 13860 29652
rect 14252 29820 14308 29876
rect 14140 29426 14196 29428
rect 14140 29374 14142 29426
rect 14142 29374 14194 29426
rect 14194 29374 14196 29426
rect 14140 29372 14196 29374
rect 14028 28754 14084 28756
rect 14028 28702 14030 28754
rect 14030 28702 14082 28754
rect 14082 28702 14084 28754
rect 14028 28700 14084 28702
rect 14140 28588 14196 28644
rect 13692 25116 13748 25172
rect 14812 38162 14868 38164
rect 14812 38110 14814 38162
rect 14814 38110 14866 38162
rect 14866 38110 14868 38162
rect 14812 38108 14868 38110
rect 14588 37772 14644 37828
rect 14924 35420 14980 35476
rect 16044 45500 16100 45556
rect 15932 44156 15988 44212
rect 16380 45948 16436 46004
rect 17836 53452 17892 53508
rect 17388 52722 17444 52724
rect 17388 52670 17390 52722
rect 17390 52670 17442 52722
rect 17442 52670 17444 52722
rect 17388 52668 17444 52670
rect 18172 53452 18228 53508
rect 17724 52722 17780 52724
rect 17724 52670 17726 52722
rect 17726 52670 17778 52722
rect 17778 52670 17780 52722
rect 17724 52668 17780 52670
rect 18060 52892 18116 52948
rect 17500 52556 17556 52612
rect 18060 52220 18116 52276
rect 17612 50428 17668 50484
rect 17052 49980 17108 50036
rect 16828 49532 16884 49588
rect 17052 48636 17108 48692
rect 17612 49868 17668 49924
rect 17948 51996 18004 52052
rect 17836 51660 17892 51716
rect 18508 56476 18564 56532
rect 18508 56194 18564 56196
rect 18508 56142 18510 56194
rect 18510 56142 18562 56194
rect 18562 56142 18564 56194
rect 18508 56140 18564 56142
rect 19180 58604 19236 58660
rect 18844 57036 18900 57092
rect 18844 56812 18900 56868
rect 19516 62130 19572 62132
rect 19516 62078 19518 62130
rect 19518 62078 19570 62130
rect 19570 62078 19572 62130
rect 19516 62076 19572 62078
rect 19404 61292 19460 61348
rect 19516 60956 19572 61012
rect 19516 59330 19572 59332
rect 19516 59278 19518 59330
rect 19518 59278 19570 59330
rect 19570 59278 19572 59330
rect 19516 59276 19572 59278
rect 19292 57036 19348 57092
rect 19404 59052 19460 59108
rect 19404 57148 19460 57204
rect 19180 56812 19236 56868
rect 18732 55916 18788 55972
rect 18508 53900 18564 53956
rect 18172 51548 18228 51604
rect 18284 52780 18340 52836
rect 17724 50540 17780 50596
rect 17500 49532 17556 49588
rect 17836 49756 17892 49812
rect 17836 49420 17892 49476
rect 17388 48412 17444 48468
rect 16492 45836 16548 45892
rect 16156 43538 16212 43540
rect 16156 43486 16158 43538
rect 16158 43486 16210 43538
rect 16210 43486 16212 43538
rect 16156 43484 16212 43486
rect 16268 44828 16324 44884
rect 15484 42194 15540 42196
rect 15484 42142 15486 42194
rect 15486 42142 15538 42194
rect 15538 42142 15540 42194
rect 15484 42140 15540 42142
rect 15932 42252 15988 42308
rect 15372 41356 15428 41412
rect 15708 41020 15764 41076
rect 15372 40572 15428 40628
rect 15596 40348 15652 40404
rect 15932 40348 15988 40404
rect 15708 40178 15764 40180
rect 15708 40126 15710 40178
rect 15710 40126 15762 40178
rect 15762 40126 15764 40178
rect 15708 40124 15764 40126
rect 15932 38780 15988 38836
rect 15260 38220 15316 38276
rect 15372 37490 15428 37492
rect 15372 37438 15374 37490
rect 15374 37438 15426 37490
rect 15426 37438 15428 37490
rect 15372 37436 15428 37438
rect 15148 36594 15204 36596
rect 15148 36542 15150 36594
rect 15150 36542 15202 36594
rect 15202 36542 15204 36594
rect 15148 36540 15204 36542
rect 15372 35420 15428 35476
rect 15148 34636 15204 34692
rect 15596 37826 15652 37828
rect 15596 37774 15598 37826
rect 15598 37774 15650 37826
rect 15650 37774 15652 37826
rect 15596 37772 15652 37774
rect 15932 38162 15988 38164
rect 15932 38110 15934 38162
rect 15934 38110 15986 38162
rect 15986 38110 15988 38162
rect 15932 38108 15988 38110
rect 15820 38050 15876 38052
rect 15820 37998 15822 38050
rect 15822 37998 15874 38050
rect 15874 37998 15876 38050
rect 15820 37996 15876 37998
rect 15932 37826 15988 37828
rect 15932 37774 15934 37826
rect 15934 37774 15986 37826
rect 15986 37774 15988 37826
rect 15932 37772 15988 37774
rect 16380 44156 16436 44212
rect 16380 43036 16436 43092
rect 16380 41132 16436 41188
rect 16716 45052 16772 45108
rect 16940 45666 16996 45668
rect 16940 45614 16942 45666
rect 16942 45614 16994 45666
rect 16994 45614 16996 45666
rect 16940 45612 16996 45614
rect 16828 44994 16884 44996
rect 16828 44942 16830 44994
rect 16830 44942 16882 44994
rect 16882 44942 16884 44994
rect 16828 44940 16884 44942
rect 17052 44828 17108 44884
rect 17164 47180 17220 47236
rect 16716 44044 16772 44100
rect 16716 43036 16772 43092
rect 17052 44210 17108 44212
rect 17052 44158 17054 44210
rect 17054 44158 17106 44210
rect 17106 44158 17108 44210
rect 17052 44156 17108 44158
rect 16828 43372 16884 43428
rect 16716 42530 16772 42532
rect 16716 42478 16718 42530
rect 16718 42478 16770 42530
rect 16770 42478 16772 42530
rect 16716 42476 16772 42478
rect 16940 43596 16996 43652
rect 16940 42140 16996 42196
rect 16940 41916 16996 41972
rect 16380 40684 16436 40740
rect 16492 40796 16548 40852
rect 16156 39452 16212 39508
rect 16268 40460 16324 40516
rect 16492 40460 16548 40516
rect 16380 38556 16436 38612
rect 16492 38780 16548 38836
rect 16156 37660 16212 37716
rect 17052 40962 17108 40964
rect 17052 40910 17054 40962
rect 17054 40910 17106 40962
rect 17106 40910 17108 40962
rect 17052 40908 17108 40910
rect 16828 40460 16884 40516
rect 16828 38722 16884 38724
rect 16828 38670 16830 38722
rect 16830 38670 16882 38722
rect 16882 38670 16884 38722
rect 16828 38668 16884 38670
rect 16828 38444 16884 38500
rect 16380 38162 16436 38164
rect 16380 38110 16382 38162
rect 16382 38110 16434 38162
rect 16434 38110 16436 38162
rect 16380 38108 16436 38110
rect 15596 35698 15652 35700
rect 15596 35646 15598 35698
rect 15598 35646 15650 35698
rect 15650 35646 15652 35698
rect 15596 35644 15652 35646
rect 15820 35586 15876 35588
rect 15820 35534 15822 35586
rect 15822 35534 15874 35586
rect 15874 35534 15876 35586
rect 15820 35532 15876 35534
rect 15932 35420 15988 35476
rect 14812 32844 14868 32900
rect 14700 32450 14756 32452
rect 14700 32398 14702 32450
rect 14702 32398 14754 32450
rect 14754 32398 14756 32450
rect 14700 32396 14756 32398
rect 15148 32562 15204 32564
rect 15148 32510 15150 32562
rect 15150 32510 15202 32562
rect 15202 32510 15204 32562
rect 15148 32508 15204 32510
rect 15260 31666 15316 31668
rect 15260 31614 15262 31666
rect 15262 31614 15314 31666
rect 15314 31614 15316 31666
rect 15260 31612 15316 31614
rect 15148 29820 15204 29876
rect 14700 29426 14756 29428
rect 14700 29374 14702 29426
rect 14702 29374 14754 29426
rect 14754 29374 14756 29426
rect 14700 29372 14756 29374
rect 13132 22428 13188 22484
rect 13132 20748 13188 20804
rect 12572 17388 12628 17444
rect 12236 16716 12292 16772
rect 12124 16156 12180 16212
rect 12908 16210 12964 16212
rect 12908 16158 12910 16210
rect 12910 16158 12962 16210
rect 12962 16158 12964 16210
rect 12908 16156 12964 16158
rect 12012 16098 12068 16100
rect 12012 16046 12014 16098
rect 12014 16046 12066 16098
rect 12066 16046 12068 16098
rect 12012 16044 12068 16046
rect 11788 15986 11844 15988
rect 11788 15934 11790 15986
rect 11790 15934 11842 15986
rect 11842 15934 11844 15986
rect 11788 15932 11844 15934
rect 11676 15260 11732 15316
rect 11340 12348 11396 12404
rect 10780 11676 10836 11732
rect 11004 11788 11060 11844
rect 10780 10834 10836 10836
rect 10780 10782 10782 10834
rect 10782 10782 10834 10834
rect 10834 10782 10836 10834
rect 10780 10780 10836 10782
rect 10668 10668 10724 10724
rect 10444 10332 10500 10388
rect 11004 10556 11060 10612
rect 10668 9884 10724 9940
rect 12236 15874 12292 15876
rect 12236 15822 12238 15874
rect 12238 15822 12290 15874
rect 12290 15822 12292 15874
rect 12236 15820 12292 15822
rect 12684 15596 12740 15652
rect 12124 15372 12180 15428
rect 12236 12402 12292 12404
rect 12236 12350 12238 12402
rect 12238 12350 12290 12402
rect 12290 12350 12292 12402
rect 12236 12348 12292 12350
rect 11676 11676 11732 11732
rect 12012 12290 12068 12292
rect 12012 12238 12014 12290
rect 12014 12238 12066 12290
rect 12066 12238 12068 12290
rect 12012 12236 12068 12238
rect 11788 11452 11844 11508
rect 12124 11676 12180 11732
rect 12348 11564 12404 11620
rect 13132 15314 13188 15316
rect 13132 15262 13134 15314
rect 13134 15262 13186 15314
rect 13186 15262 13188 15314
rect 13132 15260 13188 15262
rect 13468 23154 13524 23156
rect 13468 23102 13470 23154
rect 13470 23102 13522 23154
rect 13522 23102 13524 23154
rect 13468 23100 13524 23102
rect 15036 26908 15092 26964
rect 13804 22540 13860 22596
rect 13468 21532 13524 21588
rect 14140 21586 14196 21588
rect 14140 21534 14142 21586
rect 14142 21534 14194 21586
rect 14194 21534 14196 21586
rect 14140 21532 14196 21534
rect 13692 21196 13748 21252
rect 13692 20860 13748 20916
rect 14812 26290 14868 26292
rect 14812 26238 14814 26290
rect 14814 26238 14866 26290
rect 14866 26238 14868 26290
rect 14812 26236 14868 26238
rect 15148 23436 15204 23492
rect 14924 22370 14980 22372
rect 14924 22318 14926 22370
rect 14926 22318 14978 22370
rect 14978 22318 14980 22370
rect 14924 22316 14980 22318
rect 15148 22316 15204 22372
rect 14252 19346 14308 19348
rect 14252 19294 14254 19346
rect 14254 19294 14306 19346
rect 14306 19294 14308 19346
rect 14252 19292 14308 19294
rect 13468 19234 13524 19236
rect 13468 19182 13470 19234
rect 13470 19182 13522 19234
rect 13522 19182 13524 19234
rect 13468 19180 13524 19182
rect 15596 32732 15652 32788
rect 15596 32396 15652 32452
rect 15820 34690 15876 34692
rect 15820 34638 15822 34690
rect 15822 34638 15874 34690
rect 15874 34638 15876 34690
rect 15820 34636 15876 34638
rect 16156 33964 16212 34020
rect 16044 33852 16100 33908
rect 15820 33628 15876 33684
rect 15820 31612 15876 31668
rect 15820 30940 15876 30996
rect 15484 29538 15540 29540
rect 15484 29486 15486 29538
rect 15486 29486 15538 29538
rect 15538 29486 15540 29538
rect 15484 29484 15540 29486
rect 16604 37772 16660 37828
rect 16716 37660 16772 37716
rect 16604 37490 16660 37492
rect 16604 37438 16606 37490
rect 16606 37438 16658 37490
rect 16658 37438 16660 37490
rect 16604 37436 16660 37438
rect 16828 37436 16884 37492
rect 16828 36540 16884 36596
rect 16828 32844 16884 32900
rect 15932 29820 15988 29876
rect 16156 28476 16212 28532
rect 16268 28028 16324 28084
rect 16380 27804 16436 27860
rect 16268 27074 16324 27076
rect 16268 27022 16270 27074
rect 16270 27022 16322 27074
rect 16322 27022 16324 27074
rect 16268 27020 16324 27022
rect 15596 26962 15652 26964
rect 15596 26910 15598 26962
rect 15598 26910 15650 26962
rect 15650 26910 15652 26962
rect 15596 26908 15652 26910
rect 15820 26290 15876 26292
rect 15820 26238 15822 26290
rect 15822 26238 15874 26290
rect 15874 26238 15876 26290
rect 15820 26236 15876 26238
rect 16604 29650 16660 29652
rect 16604 29598 16606 29650
rect 16606 29598 16658 29650
rect 16658 29598 16660 29650
rect 16604 29596 16660 29598
rect 17052 37100 17108 37156
rect 17052 35644 17108 35700
rect 17052 29372 17108 29428
rect 17052 28476 17108 28532
rect 16828 27356 16884 27412
rect 17388 45500 17444 45556
rect 17500 46172 17556 46228
rect 17612 45724 17668 45780
rect 17500 44940 17556 44996
rect 17388 44380 17444 44436
rect 18844 53004 18900 53060
rect 19180 53900 19236 53956
rect 18956 52780 19012 52836
rect 19404 53058 19460 53060
rect 19404 53006 19406 53058
rect 19406 53006 19458 53058
rect 19458 53006 19460 53058
rect 19404 53004 19460 53006
rect 18396 51324 18452 51380
rect 18620 51436 18676 51492
rect 18284 50988 18340 51044
rect 18620 50988 18676 51044
rect 18620 50764 18676 50820
rect 18508 50316 18564 50372
rect 18620 49922 18676 49924
rect 18620 49870 18622 49922
rect 18622 49870 18674 49922
rect 18674 49870 18676 49922
rect 18620 49868 18676 49870
rect 18620 49026 18676 49028
rect 18620 48974 18622 49026
rect 18622 48974 18674 49026
rect 18674 48974 18676 49026
rect 18620 48972 18676 48974
rect 18732 46732 18788 46788
rect 18396 46508 18452 46564
rect 18172 46284 18228 46340
rect 18284 46450 18340 46452
rect 18284 46398 18286 46450
rect 18286 46398 18338 46450
rect 18338 46398 18340 46450
rect 18284 46396 18340 46398
rect 17724 44156 17780 44212
rect 17836 44044 17892 44100
rect 18060 41916 18116 41972
rect 17836 41020 17892 41076
rect 17612 40460 17668 40516
rect 17500 40348 17556 40404
rect 17276 40236 17332 40292
rect 17388 40124 17444 40180
rect 17612 38668 17668 38724
rect 17388 37826 17444 37828
rect 17388 37774 17390 37826
rect 17390 37774 17442 37826
rect 17442 37774 17444 37826
rect 17388 37772 17444 37774
rect 17276 36764 17332 36820
rect 17276 36594 17332 36596
rect 17276 36542 17278 36594
rect 17278 36542 17330 36594
rect 17330 36542 17332 36594
rect 17276 36540 17332 36542
rect 17500 35810 17556 35812
rect 17500 35758 17502 35810
rect 17502 35758 17554 35810
rect 17554 35758 17556 35810
rect 17500 35756 17556 35758
rect 17388 35586 17444 35588
rect 17388 35534 17390 35586
rect 17390 35534 17442 35586
rect 17442 35534 17444 35586
rect 17388 35532 17444 35534
rect 17724 37154 17780 37156
rect 17724 37102 17726 37154
rect 17726 37102 17778 37154
rect 17778 37102 17780 37154
rect 17724 37100 17780 37102
rect 17836 36764 17892 36820
rect 17836 36540 17892 36596
rect 17948 35698 18004 35700
rect 17948 35646 17950 35698
rect 17950 35646 18002 35698
rect 18002 35646 18004 35698
rect 17948 35644 18004 35646
rect 18172 40460 18228 40516
rect 18060 35420 18116 35476
rect 17724 35084 17780 35140
rect 18396 45724 18452 45780
rect 18508 44828 18564 44884
rect 18732 44380 18788 44436
rect 19836 62746 19892 62748
rect 19836 62694 19838 62746
rect 19838 62694 19890 62746
rect 19890 62694 19892 62746
rect 19836 62692 19892 62694
rect 19940 62746 19996 62748
rect 19940 62694 19942 62746
rect 19942 62694 19994 62746
rect 19994 62694 19996 62746
rect 19940 62692 19996 62694
rect 20044 62746 20100 62748
rect 20044 62694 20046 62746
rect 20046 62694 20098 62746
rect 20098 62694 20100 62746
rect 20044 62692 20100 62694
rect 20076 62466 20132 62468
rect 20076 62414 20078 62466
rect 20078 62414 20130 62466
rect 20130 62414 20132 62466
rect 20076 62412 20132 62414
rect 20076 61346 20132 61348
rect 20076 61294 20078 61346
rect 20078 61294 20130 61346
rect 20130 61294 20132 61346
rect 20076 61292 20132 61294
rect 19836 61178 19892 61180
rect 19836 61126 19838 61178
rect 19838 61126 19890 61178
rect 19890 61126 19892 61178
rect 19836 61124 19892 61126
rect 19940 61178 19996 61180
rect 19940 61126 19942 61178
rect 19942 61126 19994 61178
rect 19994 61126 19996 61178
rect 19940 61124 19996 61126
rect 20044 61178 20100 61180
rect 20044 61126 20046 61178
rect 20046 61126 20098 61178
rect 20098 61126 20100 61178
rect 20044 61124 20100 61126
rect 19836 59610 19892 59612
rect 19836 59558 19838 59610
rect 19838 59558 19890 59610
rect 19890 59558 19892 59610
rect 19836 59556 19892 59558
rect 19940 59610 19996 59612
rect 19940 59558 19942 59610
rect 19942 59558 19994 59610
rect 19994 59558 19996 59610
rect 19940 59556 19996 59558
rect 20044 59610 20100 59612
rect 20044 59558 20046 59610
rect 20046 59558 20098 59610
rect 20098 59558 20100 59610
rect 20044 59556 20100 59558
rect 20300 58492 20356 58548
rect 21420 67900 21476 67956
rect 21644 67676 21700 67732
rect 21532 67618 21588 67620
rect 21532 67566 21534 67618
rect 21534 67566 21586 67618
rect 21586 67566 21588 67618
rect 21532 67564 21588 67566
rect 21420 66386 21476 66388
rect 21420 66334 21422 66386
rect 21422 66334 21474 66386
rect 21474 66334 21476 66386
rect 21420 66332 21476 66334
rect 20524 65996 20580 66052
rect 21196 65490 21252 65492
rect 21196 65438 21198 65490
rect 21198 65438 21250 65490
rect 21250 65438 21252 65490
rect 21196 65436 21252 65438
rect 21308 65324 21364 65380
rect 20748 64706 20804 64708
rect 20748 64654 20750 64706
rect 20750 64654 20802 64706
rect 20802 64654 20804 64706
rect 20748 64652 20804 64654
rect 22204 73948 22260 74004
rect 22540 74284 22596 74340
rect 23436 78706 23492 78708
rect 23436 78654 23438 78706
rect 23438 78654 23490 78706
rect 23490 78654 23492 78706
rect 23436 78652 23492 78654
rect 22764 78594 22820 78596
rect 22764 78542 22766 78594
rect 22766 78542 22818 78594
rect 22818 78542 22820 78594
rect 22764 78540 22820 78542
rect 23660 82124 23716 82180
rect 23884 84530 23940 84532
rect 23884 84478 23886 84530
rect 23886 84478 23938 84530
rect 23938 84478 23940 84530
rect 23884 84476 23940 84478
rect 24108 88060 24164 88116
rect 25228 89068 25284 89124
rect 25116 88732 25172 88788
rect 24556 87836 24612 87892
rect 24780 87948 24836 88004
rect 24556 87554 24612 87556
rect 24556 87502 24558 87554
rect 24558 87502 24610 87554
rect 24610 87502 24612 87554
rect 24556 87500 24612 87502
rect 24668 87442 24724 87444
rect 24668 87390 24670 87442
rect 24670 87390 24722 87442
rect 24722 87390 24724 87442
rect 24668 87388 24724 87390
rect 24668 86882 24724 86884
rect 24668 86830 24670 86882
rect 24670 86830 24722 86882
rect 24722 86830 24724 86882
rect 24668 86828 24724 86830
rect 24108 86380 24164 86436
rect 24332 86156 24388 86212
rect 24892 86604 24948 86660
rect 24220 84588 24276 84644
rect 24444 84306 24500 84308
rect 24444 84254 24446 84306
rect 24446 84254 24498 84306
rect 24498 84254 24500 84306
rect 24444 84252 24500 84254
rect 24108 82348 24164 82404
rect 24220 84140 24276 84196
rect 24108 82124 24164 82180
rect 23772 80444 23828 80500
rect 23996 81228 24052 81284
rect 23660 80332 23716 80388
rect 23660 79436 23716 79492
rect 23884 79602 23940 79604
rect 23884 79550 23886 79602
rect 23886 79550 23938 79602
rect 23938 79550 23940 79602
rect 23884 79548 23940 79550
rect 24108 80444 24164 80500
rect 23884 78876 23940 78932
rect 23996 78818 24052 78820
rect 23996 78766 23998 78818
rect 23998 78766 24050 78818
rect 24050 78766 24052 78818
rect 23996 78764 24052 78766
rect 23772 77868 23828 77924
rect 22876 75068 22932 75124
rect 22540 72716 22596 72772
rect 22316 70194 22372 70196
rect 22316 70142 22318 70194
rect 22318 70142 22370 70194
rect 22370 70142 22372 70194
rect 22316 70140 22372 70142
rect 22988 74898 23044 74900
rect 22988 74846 22990 74898
rect 22990 74846 23042 74898
rect 23042 74846 23044 74898
rect 22988 74844 23044 74846
rect 23100 74060 23156 74116
rect 24108 76524 24164 76580
rect 25004 87836 25060 87892
rect 24668 86380 24724 86436
rect 24892 86044 24948 86100
rect 25116 86940 25172 86996
rect 25452 90466 25508 90468
rect 25452 90414 25454 90466
rect 25454 90414 25506 90466
rect 25506 90414 25508 90466
rect 25452 90412 25508 90414
rect 25116 86716 25172 86772
rect 26124 91868 26180 91924
rect 25788 88844 25844 88900
rect 25564 88002 25620 88004
rect 25564 87950 25566 88002
rect 25566 87950 25618 88002
rect 25618 87950 25620 88002
rect 25564 87948 25620 87950
rect 25452 87612 25508 87668
rect 25340 87500 25396 87556
rect 25228 85874 25284 85876
rect 25228 85822 25230 85874
rect 25230 85822 25282 85874
rect 25282 85822 25284 85874
rect 25228 85820 25284 85822
rect 25228 82738 25284 82740
rect 25228 82686 25230 82738
rect 25230 82686 25282 82738
rect 25282 82686 25284 82738
rect 25228 82684 25284 82686
rect 24892 82012 24948 82068
rect 25004 81900 25060 81956
rect 24780 80668 24836 80724
rect 24892 81676 24948 81732
rect 24332 78988 24388 79044
rect 25004 81228 25060 81284
rect 25004 79436 25060 79492
rect 24332 78594 24388 78596
rect 24332 78542 24334 78594
rect 24334 78542 24386 78594
rect 24386 78542 24388 78594
rect 24332 78540 24388 78542
rect 24220 76412 24276 76468
rect 24780 78540 24836 78596
rect 25900 88732 25956 88788
rect 26124 89570 26180 89572
rect 26124 89518 26126 89570
rect 26126 89518 26178 89570
rect 26178 89518 26180 89570
rect 26124 89516 26180 89518
rect 26236 89404 26292 89460
rect 26236 87612 26292 87668
rect 26124 86604 26180 86660
rect 25452 82460 25508 82516
rect 25900 85596 25956 85652
rect 25676 84530 25732 84532
rect 25676 84478 25678 84530
rect 25678 84478 25730 84530
rect 25730 84478 25732 84530
rect 25676 84476 25732 84478
rect 25788 84194 25844 84196
rect 25788 84142 25790 84194
rect 25790 84142 25842 84194
rect 25842 84142 25844 84194
rect 25788 84140 25844 84142
rect 25900 83132 25956 83188
rect 25900 82908 25956 82964
rect 25788 82348 25844 82404
rect 25452 81788 25508 81844
rect 25452 81282 25508 81284
rect 25452 81230 25454 81282
rect 25454 81230 25506 81282
rect 25506 81230 25508 81282
rect 25452 81228 25508 81230
rect 25900 82236 25956 82292
rect 25676 80892 25732 80948
rect 25452 80668 25508 80724
rect 25900 80668 25956 80724
rect 26236 84700 26292 84756
rect 26236 84476 26292 84532
rect 26236 83244 26292 83300
rect 26796 97356 26852 97412
rect 28476 97356 28532 97412
rect 26460 95788 26516 95844
rect 27356 95842 27412 95844
rect 27356 95790 27358 95842
rect 27358 95790 27410 95842
rect 27410 95790 27412 95842
rect 27356 95788 27412 95790
rect 27356 94556 27412 94612
rect 27804 95228 27860 95284
rect 27468 93884 27524 93940
rect 26684 92818 26740 92820
rect 26684 92766 26686 92818
rect 26686 92766 26738 92818
rect 26738 92766 26740 92818
rect 26684 92764 26740 92766
rect 27468 92818 27524 92820
rect 27468 92766 27470 92818
rect 27470 92766 27522 92818
rect 27522 92766 27524 92818
rect 27468 92764 27524 92766
rect 26460 92428 26516 92484
rect 27356 92146 27412 92148
rect 27356 92094 27358 92146
rect 27358 92094 27410 92146
rect 27410 92094 27412 92146
rect 27356 92092 27412 92094
rect 26572 87388 26628 87444
rect 26908 89068 26964 89124
rect 27020 87948 27076 88004
rect 27356 88620 27412 88676
rect 27356 87836 27412 87892
rect 27468 88956 27524 89012
rect 27244 87554 27300 87556
rect 27244 87502 27246 87554
rect 27246 87502 27298 87554
rect 27298 87502 27300 87554
rect 27244 87500 27300 87502
rect 27132 87164 27188 87220
rect 26908 86546 26964 86548
rect 26908 86494 26910 86546
rect 26910 86494 26962 86546
rect 26962 86494 26964 86546
rect 26908 86492 26964 86494
rect 26908 84306 26964 84308
rect 26908 84254 26910 84306
rect 26910 84254 26962 84306
rect 26962 84254 26964 84306
rect 26908 84252 26964 84254
rect 27356 85596 27412 85652
rect 27468 84924 27524 84980
rect 27356 84476 27412 84532
rect 27132 82908 27188 82964
rect 26460 82850 26516 82852
rect 26460 82798 26462 82850
rect 26462 82798 26514 82850
rect 26514 82798 26516 82850
rect 26460 82796 26516 82798
rect 26348 81900 26404 81956
rect 26572 82684 26628 82740
rect 26684 82124 26740 82180
rect 27020 82572 27076 82628
rect 26908 82460 26964 82516
rect 27132 82460 27188 82516
rect 27356 84252 27412 84308
rect 27468 84194 27524 84196
rect 27468 84142 27470 84194
rect 27470 84142 27522 84194
rect 27522 84142 27524 84194
rect 27468 84140 27524 84142
rect 27356 82572 27412 82628
rect 27244 82348 27300 82404
rect 27356 82178 27412 82180
rect 27356 82126 27358 82178
rect 27358 82126 27410 82178
rect 27410 82126 27412 82178
rect 27356 82124 27412 82126
rect 26908 81842 26964 81844
rect 26908 81790 26910 81842
rect 26910 81790 26962 81842
rect 26962 81790 26964 81842
rect 26908 81788 26964 81790
rect 27132 81676 27188 81732
rect 26012 80556 26068 80612
rect 26348 80556 26404 80612
rect 24556 76636 24612 76692
rect 23772 75010 23828 75012
rect 23772 74958 23774 75010
rect 23774 74958 23826 75010
rect 23826 74958 23828 75010
rect 23772 74956 23828 74958
rect 23884 74898 23940 74900
rect 23884 74846 23886 74898
rect 23886 74846 23938 74898
rect 23938 74846 23940 74898
rect 23884 74844 23940 74846
rect 23548 72716 23604 72772
rect 23996 72156 24052 72212
rect 24668 76412 24724 76468
rect 24556 75852 24612 75908
rect 24332 74956 24388 75012
rect 24444 75628 24500 75684
rect 24332 73388 24388 73444
rect 22876 71596 22932 71652
rect 25228 77532 25284 77588
rect 25788 80444 25844 80500
rect 25564 78988 25620 79044
rect 25788 78540 25844 78596
rect 25788 78092 25844 78148
rect 25564 77644 25620 77700
rect 25340 76690 25396 76692
rect 25340 76638 25342 76690
rect 25342 76638 25394 76690
rect 25394 76638 25396 76690
rect 25340 76636 25396 76638
rect 25228 75122 25284 75124
rect 25228 75070 25230 75122
rect 25230 75070 25282 75122
rect 25282 75070 25284 75122
rect 25228 75068 25284 75070
rect 25340 74956 25396 75012
rect 24668 73164 24724 73220
rect 24780 72716 24836 72772
rect 25228 74844 25284 74900
rect 25228 72604 25284 72660
rect 25004 72156 25060 72212
rect 24668 71650 24724 71652
rect 24668 71598 24670 71650
rect 24670 71598 24722 71650
rect 24722 71598 24724 71650
rect 24668 71596 24724 71598
rect 24332 70924 24388 70980
rect 22428 67900 22484 67956
rect 22316 67116 22372 67172
rect 22092 66668 22148 66724
rect 22316 66332 22372 66388
rect 21644 64594 21700 64596
rect 21644 64542 21646 64594
rect 21646 64542 21698 64594
rect 21698 64542 21700 64594
rect 21644 64540 21700 64542
rect 21532 64482 21588 64484
rect 21532 64430 21534 64482
rect 21534 64430 21586 64482
rect 21586 64430 21588 64482
rect 21532 64428 21588 64430
rect 20860 63980 20916 64036
rect 21196 63922 21252 63924
rect 21196 63870 21198 63922
rect 21198 63870 21250 63922
rect 21250 63870 21252 63922
rect 21196 63868 21252 63870
rect 21084 62354 21140 62356
rect 21084 62302 21086 62354
rect 21086 62302 21138 62354
rect 21138 62302 21140 62354
rect 21084 62300 21140 62302
rect 19836 58042 19892 58044
rect 19836 57990 19838 58042
rect 19838 57990 19890 58042
rect 19890 57990 19892 58042
rect 19836 57988 19892 57990
rect 19940 58042 19996 58044
rect 19940 57990 19942 58042
rect 19942 57990 19994 58042
rect 19994 57990 19996 58042
rect 19940 57988 19996 57990
rect 20044 58042 20100 58044
rect 20044 57990 20046 58042
rect 20046 57990 20098 58042
rect 20098 57990 20100 58042
rect 20044 57988 20100 57990
rect 20188 57762 20244 57764
rect 20188 57710 20190 57762
rect 20190 57710 20242 57762
rect 20242 57710 20244 57762
rect 20188 57708 20244 57710
rect 19964 57650 20020 57652
rect 19964 57598 19966 57650
rect 19966 57598 20018 57650
rect 20018 57598 20020 57650
rect 19964 57596 20020 57598
rect 19836 56474 19892 56476
rect 19836 56422 19838 56474
rect 19838 56422 19890 56474
rect 19890 56422 19892 56474
rect 19836 56420 19892 56422
rect 19940 56474 19996 56476
rect 19940 56422 19942 56474
rect 19942 56422 19994 56474
rect 19994 56422 19996 56474
rect 19940 56420 19996 56422
rect 20044 56474 20100 56476
rect 20044 56422 20046 56474
rect 20046 56422 20098 56474
rect 20098 56422 20100 56474
rect 20044 56420 20100 56422
rect 19740 56252 19796 56308
rect 19740 55410 19796 55412
rect 19740 55358 19742 55410
rect 19742 55358 19794 55410
rect 19794 55358 19796 55410
rect 19740 55356 19796 55358
rect 19836 54906 19892 54908
rect 19836 54854 19838 54906
rect 19838 54854 19890 54906
rect 19890 54854 19892 54906
rect 19836 54852 19892 54854
rect 19940 54906 19996 54908
rect 19940 54854 19942 54906
rect 19942 54854 19994 54906
rect 19994 54854 19996 54906
rect 19940 54852 19996 54854
rect 20044 54906 20100 54908
rect 20044 54854 20046 54906
rect 20046 54854 20098 54906
rect 20098 54854 20100 54906
rect 20044 54852 20100 54854
rect 19836 53338 19892 53340
rect 19836 53286 19838 53338
rect 19838 53286 19890 53338
rect 19890 53286 19892 53338
rect 19836 53284 19892 53286
rect 19940 53338 19996 53340
rect 19940 53286 19942 53338
rect 19942 53286 19994 53338
rect 19994 53286 19996 53338
rect 19940 53284 19996 53286
rect 20044 53338 20100 53340
rect 20044 53286 20046 53338
rect 20046 53286 20098 53338
rect 20098 53286 20100 53338
rect 20044 53284 20100 53286
rect 20748 60674 20804 60676
rect 20748 60622 20750 60674
rect 20750 60622 20802 60674
rect 20802 60622 20804 60674
rect 20748 60620 20804 60622
rect 21196 62188 21252 62244
rect 21420 63138 21476 63140
rect 21420 63086 21422 63138
rect 21422 63086 21474 63138
rect 21474 63086 21476 63138
rect 21420 63084 21476 63086
rect 21420 62914 21476 62916
rect 21420 62862 21422 62914
rect 21422 62862 21474 62914
rect 21474 62862 21476 62914
rect 21420 62860 21476 62862
rect 21980 65212 22036 65268
rect 22316 65324 22372 65380
rect 25564 76466 25620 76468
rect 25564 76414 25566 76466
rect 25566 76414 25618 76466
rect 25618 76414 25620 76466
rect 25564 76412 25620 76414
rect 26124 79548 26180 79604
rect 26012 78706 26068 78708
rect 26012 78654 26014 78706
rect 26014 78654 26066 78706
rect 26066 78654 26068 78706
rect 26012 78652 26068 78654
rect 26124 78146 26180 78148
rect 26124 78094 26126 78146
rect 26126 78094 26178 78146
rect 26178 78094 26180 78146
rect 26124 78092 26180 78094
rect 26012 76300 26068 76356
rect 25676 75068 25732 75124
rect 25788 75292 25844 75348
rect 25564 72716 25620 72772
rect 26348 78034 26404 78036
rect 26348 77982 26350 78034
rect 26350 77982 26402 78034
rect 26402 77982 26404 78034
rect 26348 77980 26404 77982
rect 26572 80780 26628 80836
rect 26684 81058 26740 81060
rect 26684 81006 26686 81058
rect 26686 81006 26738 81058
rect 26738 81006 26740 81058
rect 26684 81004 26740 81006
rect 26908 79548 26964 79604
rect 27132 81170 27188 81172
rect 27132 81118 27134 81170
rect 27134 81118 27186 81170
rect 27186 81118 27188 81170
rect 27132 81116 27188 81118
rect 27468 81452 27524 81508
rect 27244 79490 27300 79492
rect 27244 79438 27246 79490
rect 27246 79438 27298 79490
rect 27298 79438 27300 79490
rect 27244 79436 27300 79438
rect 27132 79100 27188 79156
rect 29148 95282 29204 95284
rect 29148 95230 29150 95282
rect 29150 95230 29202 95282
rect 29202 95230 29204 95282
rect 29148 95228 29204 95230
rect 30156 96066 30212 96068
rect 30156 96014 30158 96066
rect 30158 96014 30210 96066
rect 30210 96014 30212 96066
rect 30156 96012 30212 96014
rect 29596 95228 29652 95284
rect 30156 95228 30212 95284
rect 32284 96850 32340 96852
rect 32284 96798 32286 96850
rect 32286 96798 32338 96850
rect 32338 96798 32340 96850
rect 32284 96796 32340 96798
rect 32956 96796 33012 96852
rect 31276 96012 31332 96068
rect 30940 95676 30996 95732
rect 30492 93884 30548 93940
rect 35196 98026 35252 98028
rect 35196 97974 35198 98026
rect 35198 97974 35250 98026
rect 35250 97974 35252 98026
rect 35196 97972 35252 97974
rect 35300 98026 35356 98028
rect 35300 97974 35302 98026
rect 35302 97974 35354 98026
rect 35354 97974 35356 98026
rect 35300 97972 35356 97974
rect 35404 98026 35460 98028
rect 35404 97974 35406 98026
rect 35406 97974 35458 98026
rect 35458 97974 35460 98026
rect 35404 97972 35460 97974
rect 33404 95900 33460 95956
rect 35196 96850 35252 96852
rect 35196 96798 35198 96850
rect 35198 96798 35250 96850
rect 35250 96798 35252 96850
rect 35196 96796 35252 96798
rect 35196 96458 35252 96460
rect 35196 96406 35198 96458
rect 35198 96406 35250 96458
rect 35250 96406 35252 96458
rect 35196 96404 35252 96406
rect 35300 96458 35356 96460
rect 35300 96406 35302 96458
rect 35302 96406 35354 96458
rect 35354 96406 35356 96458
rect 35300 96404 35356 96406
rect 35404 96458 35460 96460
rect 35404 96406 35406 96458
rect 35406 96406 35458 96458
rect 35458 96406 35460 96458
rect 35404 96404 35460 96406
rect 35868 96124 35924 96180
rect 33180 95788 33236 95844
rect 33068 95282 33124 95284
rect 33068 95230 33070 95282
rect 33070 95230 33122 95282
rect 33122 95230 33124 95282
rect 33068 95228 33124 95230
rect 30940 93100 30996 93156
rect 35196 95842 35252 95844
rect 35196 95790 35198 95842
rect 35198 95790 35250 95842
rect 35250 95790 35252 95842
rect 35196 95788 35252 95790
rect 34076 95116 34132 95172
rect 35644 95282 35700 95284
rect 35644 95230 35646 95282
rect 35646 95230 35698 95282
rect 35698 95230 35700 95282
rect 35644 95228 35700 95230
rect 36428 95116 36484 95172
rect 35196 95058 35252 95060
rect 35196 95006 35198 95058
rect 35198 95006 35250 95058
rect 35250 95006 35252 95058
rect 35196 95004 35252 95006
rect 31500 93100 31556 93156
rect 31836 93996 31892 94052
rect 30156 92930 30212 92932
rect 30156 92878 30158 92930
rect 30158 92878 30210 92930
rect 30210 92878 30212 92930
rect 30156 92876 30212 92878
rect 32844 93996 32900 94052
rect 29260 92764 29316 92820
rect 31836 92764 31892 92820
rect 32508 92988 32564 93044
rect 32732 92930 32788 92932
rect 32732 92878 32734 92930
rect 32734 92878 32786 92930
rect 32786 92878 32788 92930
rect 32732 92876 32788 92878
rect 32508 92652 32564 92708
rect 28364 91980 28420 92036
rect 33180 92764 33236 92820
rect 33180 91308 33236 91364
rect 33852 92876 33908 92932
rect 37772 95058 37828 95060
rect 37772 95006 37774 95058
rect 37774 95006 37826 95058
rect 37826 95006 37828 95058
rect 37772 95004 37828 95006
rect 35196 94890 35252 94892
rect 35196 94838 35198 94890
rect 35198 94838 35250 94890
rect 35250 94838 35252 94890
rect 35196 94836 35252 94838
rect 35300 94890 35356 94892
rect 35300 94838 35302 94890
rect 35302 94838 35354 94890
rect 35354 94838 35356 94890
rect 35300 94836 35356 94838
rect 35404 94890 35460 94892
rect 35404 94838 35406 94890
rect 35406 94838 35458 94890
rect 35458 94838 35460 94890
rect 35404 94836 35460 94838
rect 34076 92706 34132 92708
rect 34076 92654 34078 92706
rect 34078 92654 34130 92706
rect 34130 92654 34132 92706
rect 34076 92652 34132 92654
rect 35196 93322 35252 93324
rect 35196 93270 35198 93322
rect 35198 93270 35250 93322
rect 35250 93270 35252 93322
rect 35196 93268 35252 93270
rect 35300 93322 35356 93324
rect 35300 93270 35302 93322
rect 35302 93270 35354 93322
rect 35354 93270 35356 93322
rect 35300 93268 35356 93270
rect 35404 93322 35460 93324
rect 35404 93270 35406 93322
rect 35406 93270 35458 93322
rect 35458 93270 35460 93322
rect 35404 93268 35460 93270
rect 35084 92652 35140 92708
rect 37660 92034 37716 92036
rect 37660 91982 37662 92034
rect 37662 91982 37714 92034
rect 37714 91982 37716 92034
rect 37660 91980 37716 91982
rect 35196 91754 35252 91756
rect 35196 91702 35198 91754
rect 35198 91702 35250 91754
rect 35250 91702 35252 91754
rect 35196 91700 35252 91702
rect 35300 91754 35356 91756
rect 35300 91702 35302 91754
rect 35302 91702 35354 91754
rect 35354 91702 35356 91754
rect 35300 91700 35356 91702
rect 35404 91754 35460 91756
rect 35404 91702 35406 91754
rect 35406 91702 35458 91754
rect 35458 91702 35460 91754
rect 35404 91700 35460 91702
rect 34524 91362 34580 91364
rect 34524 91310 34526 91362
rect 34526 91310 34578 91362
rect 34578 91310 34580 91362
rect 34524 91308 34580 91310
rect 28252 90466 28308 90468
rect 28252 90414 28254 90466
rect 28254 90414 28306 90466
rect 28306 90414 28308 90466
rect 28252 90412 28308 90414
rect 28028 89068 28084 89124
rect 29708 90690 29764 90692
rect 29708 90638 29710 90690
rect 29710 90638 29762 90690
rect 29762 90638 29764 90690
rect 29708 90636 29764 90638
rect 30156 90690 30212 90692
rect 30156 90638 30158 90690
rect 30158 90638 30210 90690
rect 30210 90638 30212 90690
rect 30156 90636 30212 90638
rect 35084 90636 35140 90692
rect 27692 88844 27748 88900
rect 27804 88114 27860 88116
rect 27804 88062 27806 88114
rect 27806 88062 27858 88114
rect 27858 88062 27860 88114
rect 27804 88060 27860 88062
rect 29260 89068 29316 89124
rect 30156 88898 30212 88900
rect 30156 88846 30158 88898
rect 30158 88846 30210 88898
rect 30210 88846 30212 88898
rect 30156 88844 30212 88846
rect 28588 88226 28644 88228
rect 28588 88174 28590 88226
rect 28590 88174 28642 88226
rect 28642 88174 28644 88226
rect 28588 88172 28644 88174
rect 29260 88226 29316 88228
rect 29260 88174 29262 88226
rect 29262 88174 29314 88226
rect 29314 88174 29316 88226
rect 29260 88172 29316 88174
rect 28028 86940 28084 86996
rect 29148 87948 29204 88004
rect 27692 86492 27748 86548
rect 27916 86434 27972 86436
rect 27916 86382 27918 86434
rect 27918 86382 27970 86434
rect 27970 86382 27972 86434
rect 27916 86380 27972 86382
rect 28924 85708 28980 85764
rect 28476 85596 28532 85652
rect 28028 84476 28084 84532
rect 27804 83692 27860 83748
rect 27692 82236 27748 82292
rect 27804 82012 27860 82068
rect 29484 87836 29540 87892
rect 29148 85148 29204 85204
rect 29596 86770 29652 86772
rect 29596 86718 29598 86770
rect 29598 86718 29650 86770
rect 29650 86718 29652 86770
rect 29596 86716 29652 86718
rect 29932 85820 29988 85876
rect 31052 88172 31108 88228
rect 32060 87612 32116 87668
rect 32508 88172 32564 88228
rect 30380 87388 30436 87444
rect 30828 86716 30884 86772
rect 30716 85708 30772 85764
rect 31052 87442 31108 87444
rect 31052 87390 31054 87442
rect 31054 87390 31106 87442
rect 31106 87390 31108 87442
rect 31052 87388 31108 87390
rect 32060 87442 32116 87444
rect 32060 87390 32062 87442
rect 32062 87390 32114 87442
rect 32114 87390 32116 87442
rect 32060 87388 32116 87390
rect 31164 85874 31220 85876
rect 31164 85822 31166 85874
rect 31166 85822 31218 85874
rect 31218 85822 31220 85874
rect 31164 85820 31220 85822
rect 28476 84364 28532 84420
rect 28476 84028 28532 84084
rect 30156 84700 30212 84756
rect 29372 84588 29428 84644
rect 28364 83580 28420 83636
rect 28364 83244 28420 83300
rect 28028 82460 28084 82516
rect 27692 81282 27748 81284
rect 27692 81230 27694 81282
rect 27694 81230 27746 81282
rect 27746 81230 27748 81282
rect 27692 81228 27748 81230
rect 28140 81452 28196 81508
rect 27692 79660 27748 79716
rect 27692 79324 27748 79380
rect 27580 78988 27636 79044
rect 27020 78764 27076 78820
rect 27132 78876 27188 78932
rect 27244 78818 27300 78820
rect 27244 78766 27246 78818
rect 27246 78766 27298 78818
rect 27298 78766 27300 78818
rect 27244 78764 27300 78766
rect 26684 78540 26740 78596
rect 27020 77644 27076 77700
rect 27244 77810 27300 77812
rect 27244 77758 27246 77810
rect 27246 77758 27298 77810
rect 27298 77758 27300 77810
rect 27244 77756 27300 77758
rect 26684 77532 26740 77588
rect 27020 77420 27076 77476
rect 26348 76860 26404 76916
rect 28588 81788 28644 81844
rect 28364 81676 28420 81732
rect 29260 83746 29316 83748
rect 29260 83694 29262 83746
rect 29262 83694 29314 83746
rect 29314 83694 29316 83746
rect 29260 83692 29316 83694
rect 29708 84418 29764 84420
rect 29708 84366 29710 84418
rect 29710 84366 29762 84418
rect 29762 84366 29764 84418
rect 29708 84364 29764 84366
rect 29596 83410 29652 83412
rect 29596 83358 29598 83410
rect 29598 83358 29650 83410
rect 29650 83358 29652 83410
rect 29596 83356 29652 83358
rect 29036 82962 29092 82964
rect 29036 82910 29038 82962
rect 29038 82910 29090 82962
rect 29090 82910 29092 82962
rect 29036 82908 29092 82910
rect 29148 82796 29204 82852
rect 28924 82572 28980 82628
rect 28812 82124 28868 82180
rect 27916 78876 27972 78932
rect 28140 78876 28196 78932
rect 28028 78764 28084 78820
rect 27468 78594 27524 78596
rect 27468 78542 27470 78594
rect 27470 78542 27522 78594
rect 27522 78542 27524 78594
rect 27468 78540 27524 78542
rect 28476 81170 28532 81172
rect 28476 81118 28478 81170
rect 28478 81118 28530 81170
rect 28530 81118 28532 81170
rect 28476 81116 28532 81118
rect 28476 80892 28532 80948
rect 28252 78540 28308 78596
rect 28364 78818 28420 78820
rect 28364 78766 28366 78818
rect 28366 78766 28418 78818
rect 28418 78766 28420 78818
rect 28364 78764 28420 78766
rect 28028 77922 28084 77924
rect 28028 77870 28030 77922
rect 28030 77870 28082 77922
rect 28082 77870 28084 77922
rect 28028 77868 28084 77870
rect 26796 76636 26852 76692
rect 26236 75292 26292 75348
rect 26348 75852 26404 75908
rect 26236 73218 26292 73220
rect 26236 73166 26238 73218
rect 26238 73166 26290 73218
rect 26290 73166 26292 73218
rect 26236 73164 26292 73166
rect 26124 73052 26180 73108
rect 26684 75852 26740 75908
rect 26796 76188 26852 76244
rect 26460 74844 26516 74900
rect 27356 76972 27412 77028
rect 27804 76748 27860 76804
rect 27244 76578 27300 76580
rect 27244 76526 27246 76578
rect 27246 76526 27298 76578
rect 27298 76526 27300 76578
rect 27244 76524 27300 76526
rect 27468 76524 27524 76580
rect 27356 76466 27412 76468
rect 27356 76414 27358 76466
rect 27358 76414 27410 76466
rect 27410 76414 27412 76466
rect 27356 76412 27412 76414
rect 27132 76300 27188 76356
rect 29372 82738 29428 82740
rect 29372 82686 29374 82738
rect 29374 82686 29426 82738
rect 29426 82686 29428 82738
rect 29372 82684 29428 82686
rect 30044 83298 30100 83300
rect 30044 83246 30046 83298
rect 30046 83246 30098 83298
rect 30098 83246 30100 83298
rect 30044 83244 30100 83246
rect 30156 83020 30212 83076
rect 29708 81676 29764 81732
rect 29820 82348 29876 82404
rect 29260 81058 29316 81060
rect 29260 81006 29262 81058
rect 29262 81006 29314 81058
rect 29314 81006 29316 81058
rect 29260 81004 29316 81006
rect 29596 81228 29652 81284
rect 28700 78764 28756 78820
rect 29372 79436 29428 79492
rect 29148 78930 29204 78932
rect 29148 78878 29150 78930
rect 29150 78878 29202 78930
rect 29202 78878 29204 78930
rect 29148 78876 29204 78878
rect 28476 78034 28532 78036
rect 28476 77982 28478 78034
rect 28478 77982 28530 78034
rect 28530 77982 28532 78034
rect 28476 77980 28532 77982
rect 28812 78204 28868 78260
rect 29148 78540 29204 78596
rect 29260 78258 29316 78260
rect 29260 78206 29262 78258
rect 29262 78206 29314 78258
rect 29314 78206 29316 78258
rect 29260 78204 29316 78206
rect 29708 78930 29764 78932
rect 29708 78878 29710 78930
rect 29710 78878 29762 78930
rect 29762 78878 29764 78930
rect 29708 78876 29764 78878
rect 29484 78818 29540 78820
rect 29484 78766 29486 78818
rect 29486 78766 29538 78818
rect 29538 78766 29540 78818
rect 29484 78764 29540 78766
rect 27916 76300 27972 76356
rect 27804 75740 27860 75796
rect 27580 75628 27636 75684
rect 27804 75292 27860 75348
rect 27020 74844 27076 74900
rect 27132 75010 27188 75012
rect 27132 74958 27134 75010
rect 27134 74958 27186 75010
rect 27186 74958 27188 75010
rect 27132 74956 27188 74958
rect 26908 73052 26964 73108
rect 26796 72380 26852 72436
rect 25564 70978 25620 70980
rect 25564 70926 25566 70978
rect 25566 70926 25618 70978
rect 25618 70926 25620 70978
rect 25564 70924 25620 70926
rect 25340 70418 25396 70420
rect 25340 70366 25342 70418
rect 25342 70366 25394 70418
rect 25394 70366 25396 70418
rect 25340 70364 25396 70366
rect 23212 66892 23268 66948
rect 22876 65212 22932 65268
rect 22540 64594 22596 64596
rect 22540 64542 22542 64594
rect 22542 64542 22594 64594
rect 22594 64542 22596 64594
rect 22540 64540 22596 64542
rect 21868 64034 21924 64036
rect 21868 63982 21870 64034
rect 21870 63982 21922 64034
rect 21922 63982 21924 64034
rect 21868 63980 21924 63982
rect 22876 63084 22932 63140
rect 22204 62972 22260 63028
rect 21420 61682 21476 61684
rect 21420 61630 21422 61682
rect 21422 61630 21474 61682
rect 21474 61630 21476 61682
rect 21420 61628 21476 61630
rect 21196 60786 21252 60788
rect 21196 60734 21198 60786
rect 21198 60734 21250 60786
rect 21250 60734 21252 60786
rect 21196 60732 21252 60734
rect 21084 60396 21140 60452
rect 20636 60284 20692 60340
rect 21756 61628 21812 61684
rect 21644 60396 21700 60452
rect 20412 53730 20468 53732
rect 20412 53678 20414 53730
rect 20414 53678 20466 53730
rect 20466 53678 20468 53730
rect 20412 53676 20468 53678
rect 20300 53564 20356 53620
rect 19964 52444 20020 52500
rect 20076 52162 20132 52164
rect 20076 52110 20078 52162
rect 20078 52110 20130 52162
rect 20130 52110 20132 52162
rect 20076 52108 20132 52110
rect 19964 51996 20020 52052
rect 18844 51884 18900 51940
rect 19836 51770 19892 51772
rect 19180 51660 19236 51716
rect 19628 51660 19684 51716
rect 19836 51718 19838 51770
rect 19838 51718 19890 51770
rect 19890 51718 19892 51770
rect 19836 51716 19892 51718
rect 19940 51770 19996 51772
rect 19940 51718 19942 51770
rect 19942 51718 19994 51770
rect 19994 51718 19996 51770
rect 19940 51716 19996 51718
rect 20044 51770 20100 51772
rect 20044 51718 20046 51770
rect 20046 51718 20098 51770
rect 20098 51718 20100 51770
rect 20044 51716 20100 51718
rect 19516 51548 19572 51604
rect 19180 51100 19236 51156
rect 19404 51324 19460 51380
rect 19516 50482 19572 50484
rect 19516 50430 19518 50482
rect 19518 50430 19570 50482
rect 19570 50430 19572 50482
rect 19516 50428 19572 50430
rect 19404 50034 19460 50036
rect 19404 49982 19406 50034
rect 19406 49982 19458 50034
rect 19458 49982 19460 50034
rect 19404 49980 19460 49982
rect 18508 41020 18564 41076
rect 18508 40684 18564 40740
rect 18508 40460 18564 40516
rect 19068 47180 19124 47236
rect 19068 45948 19124 46004
rect 19068 45724 19124 45780
rect 19404 49196 19460 49252
rect 19404 48524 19460 48580
rect 19516 46674 19572 46676
rect 19516 46622 19518 46674
rect 19518 46622 19570 46674
rect 19570 46622 19572 46674
rect 19516 46620 19572 46622
rect 19404 46284 19460 46340
rect 19404 45388 19460 45444
rect 18396 39058 18452 39060
rect 18396 39006 18398 39058
rect 18398 39006 18450 39058
rect 18450 39006 18452 39058
rect 18396 39004 18452 39006
rect 18284 38444 18340 38500
rect 18284 37490 18340 37492
rect 18284 37438 18286 37490
rect 18286 37438 18338 37490
rect 18338 37438 18340 37490
rect 18284 37436 18340 37438
rect 18620 38780 18676 38836
rect 19068 43596 19124 43652
rect 19068 43148 19124 43204
rect 18732 37436 18788 37492
rect 18508 36594 18564 36596
rect 18508 36542 18510 36594
rect 18510 36542 18562 36594
rect 18562 36542 18564 36594
rect 18508 36540 18564 36542
rect 18620 37324 18676 37380
rect 18620 35644 18676 35700
rect 18732 35586 18788 35588
rect 18732 35534 18734 35586
rect 18734 35534 18786 35586
rect 18786 35534 18788 35586
rect 18732 35532 18788 35534
rect 18396 35474 18452 35476
rect 18396 35422 18398 35474
rect 18398 35422 18450 35474
rect 18450 35422 18452 35474
rect 18396 35420 18452 35422
rect 18172 34972 18228 35028
rect 18284 35308 18340 35364
rect 17388 34524 17444 34580
rect 17500 34860 17556 34916
rect 17388 33516 17444 33572
rect 18172 34802 18228 34804
rect 18172 34750 18174 34802
rect 18174 34750 18226 34802
rect 18226 34750 18228 34802
rect 18172 34748 18228 34750
rect 18060 34300 18116 34356
rect 17612 33852 17668 33908
rect 17948 33964 18004 34020
rect 17836 33516 17892 33572
rect 17276 32732 17332 32788
rect 17612 33404 17668 33460
rect 17500 32844 17556 32900
rect 17836 32844 17892 32900
rect 17612 32284 17668 32340
rect 18060 32338 18116 32340
rect 18060 32286 18062 32338
rect 18062 32286 18114 32338
rect 18114 32286 18116 32338
rect 18060 32284 18116 32286
rect 18060 30716 18116 30772
rect 17388 29596 17444 29652
rect 17948 28476 18004 28532
rect 17612 28082 17668 28084
rect 17612 28030 17614 28082
rect 17614 28030 17666 28082
rect 17666 28030 17668 28082
rect 17612 28028 17668 28030
rect 17836 28140 17892 28196
rect 17724 27970 17780 27972
rect 17724 27918 17726 27970
rect 17726 27918 17778 27970
rect 17778 27918 17780 27970
rect 17724 27916 17780 27918
rect 17388 27858 17444 27860
rect 17388 27806 17390 27858
rect 17390 27806 17442 27858
rect 17442 27806 17444 27858
rect 17388 27804 17444 27806
rect 17500 27356 17556 27412
rect 16716 26796 16772 26852
rect 16940 27074 16996 27076
rect 16940 27022 16942 27074
rect 16942 27022 16994 27074
rect 16994 27022 16996 27074
rect 16940 27020 16996 27022
rect 16604 26460 16660 26516
rect 15484 26012 15540 26068
rect 16156 26066 16212 26068
rect 16156 26014 16158 26066
rect 16158 26014 16210 26066
rect 16210 26014 16212 26066
rect 16156 26012 16212 26014
rect 15484 25340 15540 25396
rect 15484 23884 15540 23940
rect 15820 23660 15876 23716
rect 15484 22316 15540 22372
rect 15708 22146 15764 22148
rect 15708 22094 15710 22146
rect 15710 22094 15762 22146
rect 15762 22094 15764 22146
rect 15708 22092 15764 22094
rect 16268 23548 16324 23604
rect 16716 23660 16772 23716
rect 17164 26908 17220 26964
rect 17052 26012 17108 26068
rect 17276 26684 17332 26740
rect 16716 23212 16772 23268
rect 15484 21196 15540 21252
rect 15372 18284 15428 18340
rect 13356 17500 13412 17556
rect 13468 17442 13524 17444
rect 13468 17390 13470 17442
rect 13470 17390 13522 17442
rect 13522 17390 13524 17442
rect 13468 17388 13524 17390
rect 13804 16210 13860 16212
rect 13804 16158 13806 16210
rect 13806 16158 13858 16210
rect 13858 16158 13860 16210
rect 13804 16156 13860 16158
rect 14700 16828 14756 16884
rect 16828 22988 16884 23044
rect 16156 22316 16212 22372
rect 16380 21756 16436 21812
rect 15596 16882 15652 16884
rect 15596 16830 15598 16882
rect 15598 16830 15650 16882
rect 15650 16830 15652 16882
rect 15596 16828 15652 16830
rect 14700 16492 14756 16548
rect 14476 16098 14532 16100
rect 14476 16046 14478 16098
rect 14478 16046 14530 16098
rect 14530 16046 14532 16098
rect 14476 16044 14532 16046
rect 14252 15932 14308 15988
rect 13356 12236 13412 12292
rect 13804 12402 13860 12404
rect 13804 12350 13806 12402
rect 13806 12350 13858 12402
rect 13858 12350 13860 12402
rect 13804 12348 13860 12350
rect 12908 11506 12964 11508
rect 12908 11454 12910 11506
rect 12910 11454 12962 11506
rect 12962 11454 12964 11506
rect 12908 11452 12964 11454
rect 12124 11116 12180 11172
rect 11788 10834 11844 10836
rect 11788 10782 11790 10834
rect 11790 10782 11842 10834
rect 11842 10782 11844 10834
rect 11788 10780 11844 10782
rect 11564 9938 11620 9940
rect 11564 9886 11566 9938
rect 11566 9886 11618 9938
rect 11618 9886 11620 9938
rect 11564 9884 11620 9886
rect 10780 9212 10836 9268
rect 10332 7084 10388 7140
rect 10668 7698 10724 7700
rect 10668 7646 10670 7698
rect 10670 7646 10722 7698
rect 10722 7646 10724 7698
rect 10668 7644 10724 7646
rect 10444 6860 10500 6916
rect 10444 6690 10500 6692
rect 10444 6638 10446 6690
rect 10446 6638 10498 6690
rect 10498 6638 10500 6690
rect 10444 6636 10500 6638
rect 10780 6914 10836 6916
rect 10780 6862 10782 6914
rect 10782 6862 10834 6914
rect 10834 6862 10836 6914
rect 10780 6860 10836 6862
rect 11116 7644 11172 7700
rect 10892 6748 10948 6804
rect 10668 6524 10724 6580
rect 9324 5516 9380 5572
rect 8316 3554 8372 3556
rect 8316 3502 8318 3554
rect 8318 3502 8370 3554
rect 8370 3502 8372 3554
rect 8316 3500 8372 3502
rect 8764 3500 8820 3556
rect 6748 1762 6804 1764
rect 6748 1710 6750 1762
rect 6750 1710 6802 1762
rect 6802 1710 6804 1762
rect 6748 1708 6804 1710
rect 9772 4562 9828 4564
rect 9772 4510 9774 4562
rect 9774 4510 9826 4562
rect 9826 4510 9828 4562
rect 9772 4508 9828 4510
rect 10780 4508 10836 4564
rect 10108 4338 10164 4340
rect 10108 4286 10110 4338
rect 10110 4286 10162 4338
rect 10162 4286 10164 4338
rect 10108 4284 10164 4286
rect 9100 3388 9156 3444
rect 9772 2658 9828 2660
rect 9772 2606 9774 2658
rect 9774 2606 9826 2658
rect 9826 2606 9828 2658
rect 9772 2604 9828 2606
rect 11452 6860 11508 6916
rect 12124 6914 12180 6916
rect 12124 6862 12126 6914
rect 12126 6862 12178 6914
rect 12178 6862 12180 6914
rect 12124 6860 12180 6862
rect 12460 11170 12516 11172
rect 12460 11118 12462 11170
rect 12462 11118 12514 11170
rect 12514 11118 12516 11170
rect 12460 11116 12516 11118
rect 14588 15148 14644 15204
rect 14476 14252 14532 14308
rect 14364 12124 14420 12180
rect 13356 11116 13412 11172
rect 13468 7644 13524 7700
rect 14476 11116 14532 11172
rect 14476 7698 14532 7700
rect 14476 7646 14478 7698
rect 14478 7646 14530 7698
rect 14530 7646 14532 7698
rect 14476 7644 14532 7646
rect 13692 6860 13748 6916
rect 14364 6914 14420 6916
rect 14364 6862 14366 6914
rect 14366 6862 14418 6914
rect 14418 6862 14420 6914
rect 14364 6860 14420 6862
rect 15148 16044 15204 16100
rect 16828 22092 16884 22148
rect 16716 21756 16772 21812
rect 16268 17106 16324 17108
rect 16268 17054 16270 17106
rect 16270 17054 16322 17106
rect 16322 17054 16324 17106
rect 16268 17052 16324 17054
rect 16828 19234 16884 19236
rect 16828 19182 16830 19234
rect 16830 19182 16882 19234
rect 16882 19182 16884 19234
rect 16828 19180 16884 19182
rect 17388 26514 17444 26516
rect 17388 26462 17390 26514
rect 17390 26462 17442 26514
rect 17442 26462 17444 26514
rect 17388 26460 17444 26462
rect 18396 34076 18452 34132
rect 17724 26066 17780 26068
rect 17724 26014 17726 26066
rect 17726 26014 17778 26066
rect 17778 26014 17780 26066
rect 17724 26012 17780 26014
rect 18396 30156 18452 30212
rect 18956 38722 19012 38724
rect 18956 38670 18958 38722
rect 18958 38670 19010 38722
rect 19010 38670 19012 38722
rect 18956 38668 19012 38670
rect 19180 41970 19236 41972
rect 19180 41918 19182 41970
rect 19182 41918 19234 41970
rect 19234 41918 19236 41970
rect 19180 41916 19236 41918
rect 19180 41020 19236 41076
rect 19180 40796 19236 40852
rect 19180 39004 19236 39060
rect 19180 38834 19236 38836
rect 19180 38782 19182 38834
rect 19182 38782 19234 38834
rect 19234 38782 19236 38834
rect 19180 38780 19236 38782
rect 19516 42140 19572 42196
rect 19516 41970 19572 41972
rect 19516 41918 19518 41970
rect 19518 41918 19570 41970
rect 19570 41918 19572 41970
rect 19516 41916 19572 41918
rect 19516 41020 19572 41076
rect 19516 39452 19572 39508
rect 19516 38780 19572 38836
rect 19404 38444 19460 38500
rect 19292 35586 19348 35588
rect 19292 35534 19294 35586
rect 19294 35534 19346 35586
rect 19346 35534 19348 35586
rect 19292 35532 19348 35534
rect 18956 34972 19012 35028
rect 18620 34524 18676 34580
rect 18844 34690 18900 34692
rect 18844 34638 18846 34690
rect 18846 34638 18898 34690
rect 18898 34638 18900 34690
rect 18844 34636 18900 34638
rect 19180 34524 19236 34580
rect 18956 34300 19012 34356
rect 18844 34130 18900 34132
rect 18844 34078 18846 34130
rect 18846 34078 18898 34130
rect 18898 34078 18900 34130
rect 18844 34076 18900 34078
rect 18844 30322 18900 30324
rect 18844 30270 18846 30322
rect 18846 30270 18898 30322
rect 18898 30270 18900 30322
rect 18844 30268 18900 30270
rect 18508 29708 18564 29764
rect 18396 28700 18452 28756
rect 18732 29596 18788 29652
rect 18620 28642 18676 28644
rect 18620 28590 18622 28642
rect 18622 28590 18674 28642
rect 18674 28590 18676 28642
rect 18620 28588 18676 28590
rect 18508 28082 18564 28084
rect 18508 28030 18510 28082
rect 18510 28030 18562 28082
rect 18562 28030 18564 28082
rect 18508 28028 18564 28030
rect 18284 23548 18340 23604
rect 18172 23436 18228 23492
rect 17388 23212 17444 23268
rect 17948 23212 18004 23268
rect 17612 23042 17668 23044
rect 17612 22990 17614 23042
rect 17614 22990 17666 23042
rect 17666 22990 17668 23042
rect 17612 22988 17668 22990
rect 18172 23042 18228 23044
rect 18172 22990 18174 23042
rect 18174 22990 18226 23042
rect 18226 22990 18228 23042
rect 18172 22988 18228 22990
rect 17388 22316 17444 22372
rect 18620 27804 18676 27860
rect 18508 23324 18564 23380
rect 18508 22540 18564 22596
rect 18508 22258 18564 22260
rect 18508 22206 18510 22258
rect 18510 22206 18562 22258
rect 18562 22206 18564 22258
rect 18508 22204 18564 22206
rect 17388 21420 17444 21476
rect 17052 19180 17108 19236
rect 17388 20802 17444 20804
rect 17388 20750 17390 20802
rect 17390 20750 17442 20802
rect 17442 20750 17444 20802
rect 17388 20748 17444 20750
rect 17276 19346 17332 19348
rect 17276 19294 17278 19346
rect 17278 19294 17330 19346
rect 17330 19294 17332 19346
rect 17276 19292 17332 19294
rect 17276 19068 17332 19124
rect 16940 18172 16996 18228
rect 16716 16940 16772 16996
rect 16380 16770 16436 16772
rect 16380 16718 16382 16770
rect 16382 16718 16434 16770
rect 16434 16718 16436 16770
rect 16380 16716 16436 16718
rect 16156 16492 16212 16548
rect 16940 17948 16996 18004
rect 15820 15596 15876 15652
rect 14924 15260 14980 15316
rect 16044 15202 16100 15204
rect 16044 15150 16046 15202
rect 16046 15150 16098 15202
rect 16098 15150 16100 15202
rect 16044 15148 16100 15150
rect 16492 15538 16548 15540
rect 16492 15486 16494 15538
rect 16494 15486 16546 15538
rect 16546 15486 16548 15538
rect 16492 15484 16548 15486
rect 16492 15260 16548 15316
rect 15148 14306 15204 14308
rect 15148 14254 15150 14306
rect 15150 14254 15202 14306
rect 15202 14254 15204 14306
rect 15148 14252 15204 14254
rect 15148 13580 15204 13636
rect 16156 13020 16212 13076
rect 15484 12402 15540 12404
rect 15484 12350 15486 12402
rect 15486 12350 15538 12402
rect 15538 12350 15540 12402
rect 15484 12348 15540 12350
rect 15932 12348 15988 12404
rect 14812 12124 14868 12180
rect 16492 12348 16548 12404
rect 16604 12460 16660 12516
rect 15932 12178 15988 12180
rect 15932 12126 15934 12178
rect 15934 12126 15986 12178
rect 15986 12126 15988 12178
rect 15932 12124 15988 12126
rect 16268 12178 16324 12180
rect 16268 12126 16270 12178
rect 16270 12126 16322 12178
rect 16322 12126 16324 12178
rect 16268 12124 16324 12126
rect 15708 11228 15764 11284
rect 15148 11170 15204 11172
rect 15148 11118 15150 11170
rect 15150 11118 15202 11170
rect 15202 11118 15204 11170
rect 15148 11116 15204 11118
rect 15820 10780 15876 10836
rect 16156 10834 16212 10836
rect 16156 10782 16158 10834
rect 16158 10782 16210 10834
rect 16210 10782 16212 10834
rect 16156 10780 16212 10782
rect 15820 10444 15876 10500
rect 16604 11282 16660 11284
rect 16604 11230 16606 11282
rect 16606 11230 16658 11282
rect 16658 11230 16660 11282
rect 16604 11228 16660 11230
rect 16604 10780 16660 10836
rect 16380 9938 16436 9940
rect 16380 9886 16382 9938
rect 16382 9886 16434 9938
rect 16434 9886 16436 9938
rect 16380 9884 16436 9886
rect 15932 8034 15988 8036
rect 15932 7982 15934 8034
rect 15934 7982 15986 8034
rect 15986 7982 15988 8034
rect 15932 7980 15988 7982
rect 16940 17052 16996 17108
rect 17052 13074 17108 13076
rect 17052 13022 17054 13074
rect 17054 13022 17106 13074
rect 17106 13022 17108 13074
rect 17052 13020 17108 13022
rect 17388 17948 17444 18004
rect 17724 21420 17780 21476
rect 18844 23884 18900 23940
rect 18844 23714 18900 23716
rect 18844 23662 18846 23714
rect 18846 23662 18898 23714
rect 18898 23662 18900 23714
rect 18844 23660 18900 23662
rect 18284 20748 18340 20804
rect 18060 18226 18116 18228
rect 18060 18174 18062 18226
rect 18062 18174 18114 18226
rect 18114 18174 18116 18226
rect 18060 18172 18116 18174
rect 17500 17106 17556 17108
rect 17500 17054 17502 17106
rect 17502 17054 17554 17106
rect 17554 17054 17556 17106
rect 17500 17052 17556 17054
rect 17612 16940 17668 16996
rect 17388 16716 17444 16772
rect 17948 16994 18004 16996
rect 17948 16942 17950 16994
rect 17950 16942 18002 16994
rect 18002 16942 18004 16994
rect 17948 16940 18004 16942
rect 18284 16492 18340 16548
rect 18732 16716 18788 16772
rect 17836 16268 17892 16324
rect 18732 15484 18788 15540
rect 17836 15426 17892 15428
rect 17836 15374 17838 15426
rect 17838 15374 17890 15426
rect 17890 15374 17892 15426
rect 17836 15372 17892 15374
rect 18172 15260 18228 15316
rect 18284 15202 18340 15204
rect 18284 15150 18286 15202
rect 18286 15150 18338 15202
rect 18338 15150 18340 15202
rect 18284 15148 18340 15150
rect 19292 34300 19348 34356
rect 19180 32172 19236 32228
rect 19516 37490 19572 37492
rect 19516 37438 19518 37490
rect 19518 37438 19570 37490
rect 19570 37438 19572 37490
rect 19516 37436 19572 37438
rect 20636 57596 20692 57652
rect 20860 55356 20916 55412
rect 20748 53900 20804 53956
rect 20636 53676 20692 53732
rect 20524 53004 20580 53060
rect 20300 52050 20356 52052
rect 20300 51998 20302 52050
rect 20302 51998 20354 52050
rect 20354 51998 20356 52050
rect 20300 51996 20356 51998
rect 20636 52946 20692 52948
rect 20636 52894 20638 52946
rect 20638 52894 20690 52946
rect 20690 52894 20692 52946
rect 20636 52892 20692 52894
rect 20748 52780 20804 52836
rect 20860 52162 20916 52164
rect 20860 52110 20862 52162
rect 20862 52110 20914 52162
rect 20914 52110 20916 52162
rect 20860 52108 20916 52110
rect 20524 51436 20580 51492
rect 20076 50428 20132 50484
rect 19836 50202 19892 50204
rect 19836 50150 19838 50202
rect 19838 50150 19890 50202
rect 19890 50150 19892 50202
rect 19836 50148 19892 50150
rect 19940 50202 19996 50204
rect 19940 50150 19942 50202
rect 19942 50150 19994 50202
rect 19994 50150 19996 50202
rect 19940 50148 19996 50150
rect 20044 50202 20100 50204
rect 20044 50150 20046 50202
rect 20046 50150 20098 50202
rect 20098 50150 20100 50202
rect 20044 50148 20100 50150
rect 20412 50092 20468 50148
rect 20636 50540 20692 50596
rect 20188 49810 20244 49812
rect 20188 49758 20190 49810
rect 20190 49758 20242 49810
rect 20242 49758 20244 49810
rect 20188 49756 20244 49758
rect 19836 48634 19892 48636
rect 19836 48582 19838 48634
rect 19838 48582 19890 48634
rect 19890 48582 19892 48634
rect 19836 48580 19892 48582
rect 19940 48634 19996 48636
rect 19940 48582 19942 48634
rect 19942 48582 19994 48634
rect 19994 48582 19996 48634
rect 19940 48580 19996 48582
rect 20044 48634 20100 48636
rect 20044 48582 20046 48634
rect 20046 48582 20098 48634
rect 20098 48582 20100 48634
rect 20044 48580 20100 48582
rect 20076 47234 20132 47236
rect 20076 47182 20078 47234
rect 20078 47182 20130 47234
rect 20130 47182 20132 47234
rect 20076 47180 20132 47182
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 19964 46786 20020 46788
rect 19964 46734 19966 46786
rect 19966 46734 20018 46786
rect 20018 46734 20020 46786
rect 19964 46732 20020 46734
rect 19852 45778 19908 45780
rect 19852 45726 19854 45778
rect 19854 45726 19906 45778
rect 19906 45726 19908 45778
rect 19852 45724 19908 45726
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 20300 44434 20356 44436
rect 20300 44382 20302 44434
rect 20302 44382 20354 44434
rect 20354 44382 20356 44434
rect 20300 44380 20356 44382
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 19852 43372 19908 43428
rect 20524 49532 20580 49588
rect 20860 49980 20916 50036
rect 20748 49922 20804 49924
rect 20748 49870 20750 49922
rect 20750 49870 20802 49922
rect 20802 49870 20804 49922
rect 20748 49868 20804 49870
rect 20524 48188 20580 48244
rect 20524 45890 20580 45892
rect 20524 45838 20526 45890
rect 20526 45838 20578 45890
rect 20578 45838 20580 45890
rect 20524 45836 20580 45838
rect 20412 43820 20468 43876
rect 20860 47068 20916 47124
rect 20860 46508 20916 46564
rect 20748 44828 20804 44884
rect 20412 43148 20468 43204
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 20076 42028 20132 42084
rect 20076 40908 20132 40964
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 19964 36988 20020 37044
rect 19628 36428 19684 36484
rect 19628 36204 19684 36260
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19964 35868 20020 35924
rect 20076 35532 20132 35588
rect 19628 35308 19684 35364
rect 19628 34748 19684 34804
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19516 33852 19572 33908
rect 19852 33964 19908 34020
rect 19740 33516 19796 33572
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19628 32172 19684 32228
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19516 31052 19572 31108
rect 19404 30434 19460 30436
rect 19404 30382 19406 30434
rect 19406 30382 19458 30434
rect 19458 30382 19460 30434
rect 19404 30380 19460 30382
rect 19180 30322 19236 30324
rect 19180 30270 19182 30322
rect 19182 30270 19234 30322
rect 19234 30270 19236 30322
rect 19180 30268 19236 30270
rect 19628 30380 19684 30436
rect 19852 30994 19908 30996
rect 19852 30942 19854 30994
rect 19854 30942 19906 30994
rect 19906 30942 19908 30994
rect 19852 30940 19908 30942
rect 19964 30828 20020 30884
rect 19068 29820 19124 29876
rect 19068 29372 19124 29428
rect 19964 30156 20020 30212
rect 19068 25340 19124 25396
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 20748 42866 20804 42868
rect 20748 42814 20750 42866
rect 20750 42814 20802 42866
rect 20802 42814 20804 42866
rect 20748 42812 20804 42814
rect 20636 42364 20692 42420
rect 20300 41916 20356 41972
rect 20748 41916 20804 41972
rect 20412 40514 20468 40516
rect 20412 40462 20414 40514
rect 20414 40462 20466 40514
rect 20466 40462 20468 40514
rect 20412 40460 20468 40462
rect 20636 41580 20692 41636
rect 20860 40908 20916 40964
rect 20300 38668 20356 38724
rect 20412 39004 20468 39060
rect 20300 37212 20356 37268
rect 20524 37884 20580 37940
rect 20748 37996 20804 38052
rect 20524 36652 20580 36708
rect 20300 29932 20356 29988
rect 20300 29484 20356 29540
rect 20188 28530 20244 28532
rect 20188 28478 20190 28530
rect 20190 28478 20242 28530
rect 20242 28478 20244 28530
rect 20188 28476 20244 28478
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 20076 27858 20132 27860
rect 20076 27806 20078 27858
rect 20078 27806 20130 27858
rect 20130 27806 20132 27858
rect 20076 27804 20132 27806
rect 20300 27074 20356 27076
rect 20300 27022 20302 27074
rect 20302 27022 20354 27074
rect 20354 27022 20356 27074
rect 20300 27020 20356 27022
rect 19068 23378 19124 23380
rect 19068 23326 19070 23378
rect 19070 23326 19122 23378
rect 19122 23326 19124 23378
rect 19068 23324 19124 23326
rect 19180 22370 19236 22372
rect 19180 22318 19182 22370
rect 19182 22318 19234 22370
rect 19234 22318 19236 22370
rect 19180 22316 19236 22318
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19628 25228 19684 25284
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 20524 28476 20580 28532
rect 21532 59388 21588 59444
rect 21420 58434 21476 58436
rect 21420 58382 21422 58434
rect 21422 58382 21474 58434
rect 21474 58382 21476 58434
rect 21420 58380 21476 58382
rect 21420 55074 21476 55076
rect 21420 55022 21422 55074
rect 21422 55022 21474 55074
rect 21474 55022 21476 55074
rect 21420 55020 21476 55022
rect 21308 52946 21364 52948
rect 21308 52894 21310 52946
rect 21310 52894 21362 52946
rect 21362 52894 21364 52946
rect 21308 52892 21364 52894
rect 21084 52108 21140 52164
rect 21084 49644 21140 49700
rect 21084 46732 21140 46788
rect 21084 45724 21140 45780
rect 21868 57484 21924 57540
rect 22092 57036 22148 57092
rect 22092 55410 22148 55412
rect 22092 55358 22094 55410
rect 22094 55358 22146 55410
rect 22146 55358 22148 55410
rect 22092 55356 22148 55358
rect 22092 55132 22148 55188
rect 21868 55020 21924 55076
rect 23212 65490 23268 65492
rect 23212 65438 23214 65490
rect 23214 65438 23266 65490
rect 23266 65438 23268 65490
rect 23212 65436 23268 65438
rect 23212 64316 23268 64372
rect 23324 63980 23380 64036
rect 23548 63922 23604 63924
rect 23548 63870 23550 63922
rect 23550 63870 23602 63922
rect 23602 63870 23604 63922
rect 23548 63868 23604 63870
rect 23996 65490 24052 65492
rect 23996 65438 23998 65490
rect 23998 65438 24050 65490
rect 24050 65438 24052 65490
rect 23996 65436 24052 65438
rect 24220 65378 24276 65380
rect 24220 65326 24222 65378
rect 24222 65326 24274 65378
rect 24274 65326 24276 65378
rect 24220 65324 24276 65326
rect 24108 65212 24164 65268
rect 24108 64706 24164 64708
rect 24108 64654 24110 64706
rect 24110 64654 24162 64706
rect 24162 64654 24164 64706
rect 24108 64652 24164 64654
rect 23884 64540 23940 64596
rect 23772 64316 23828 64372
rect 24332 64316 24388 64372
rect 23884 63868 23940 63924
rect 23100 62972 23156 63028
rect 23100 62578 23156 62580
rect 23100 62526 23102 62578
rect 23102 62526 23154 62578
rect 23154 62526 23156 62578
rect 23100 62524 23156 62526
rect 22316 62188 22372 62244
rect 22652 61292 22708 61348
rect 22540 60956 22596 61012
rect 22316 57596 22372 57652
rect 22428 60620 22484 60676
rect 21532 54460 21588 54516
rect 21644 53954 21700 53956
rect 21644 53902 21646 53954
rect 21646 53902 21698 53954
rect 21698 53902 21700 53954
rect 21644 53900 21700 53902
rect 21868 53618 21924 53620
rect 21868 53566 21870 53618
rect 21870 53566 21922 53618
rect 21922 53566 21924 53618
rect 21868 53564 21924 53566
rect 23212 62188 23268 62244
rect 22988 61292 23044 61348
rect 23100 61964 23156 62020
rect 23100 60956 23156 61012
rect 22764 60786 22820 60788
rect 22764 60734 22766 60786
rect 22766 60734 22818 60786
rect 22818 60734 22820 60786
rect 22764 60732 22820 60734
rect 23660 63756 23716 63812
rect 23212 59106 23268 59108
rect 23212 59054 23214 59106
rect 23214 59054 23266 59106
rect 23266 59054 23268 59106
rect 23212 59052 23268 59054
rect 24220 63922 24276 63924
rect 24220 63870 24222 63922
rect 24222 63870 24274 63922
rect 24274 63870 24276 63922
rect 24220 63868 24276 63870
rect 24332 63756 24388 63812
rect 26012 71596 26068 71652
rect 25900 70476 25956 70532
rect 26460 70588 26516 70644
rect 27580 73500 27636 73556
rect 27804 74060 27860 74116
rect 29260 77250 29316 77252
rect 29260 77198 29262 77250
rect 29262 77198 29314 77250
rect 29314 77198 29316 77250
rect 29260 77196 29316 77198
rect 28364 76748 28420 76804
rect 28588 76972 28644 77028
rect 29708 77196 29764 77252
rect 29708 77026 29764 77028
rect 29708 76974 29710 77026
rect 29710 76974 29762 77026
rect 29762 76974 29764 77026
rect 29708 76972 29764 76974
rect 28252 76242 28308 76244
rect 28252 76190 28254 76242
rect 28254 76190 28306 76242
rect 28306 76190 28308 76242
rect 28252 76188 28308 76190
rect 28700 75852 28756 75908
rect 28364 75516 28420 75572
rect 27804 73052 27860 73108
rect 28476 74732 28532 74788
rect 28364 74114 28420 74116
rect 28364 74062 28366 74114
rect 28366 74062 28418 74114
rect 28418 74062 28420 74114
rect 28364 74060 28420 74062
rect 27804 72546 27860 72548
rect 27804 72494 27806 72546
rect 27806 72494 27858 72546
rect 27858 72494 27860 72546
rect 27804 72492 27860 72494
rect 27132 70588 27188 70644
rect 25788 70252 25844 70308
rect 26796 69916 26852 69972
rect 27692 70700 27748 70756
rect 27468 70476 27524 70532
rect 27356 69916 27412 69972
rect 26124 69356 26180 69412
rect 26684 69410 26740 69412
rect 26684 69358 26686 69410
rect 26686 69358 26738 69410
rect 26738 69358 26740 69410
rect 26684 69356 26740 69358
rect 27468 69244 27524 69300
rect 28140 73612 28196 73668
rect 28028 73052 28084 73108
rect 28364 73330 28420 73332
rect 28364 73278 28366 73330
rect 28366 73278 28418 73330
rect 28418 73278 28420 73330
rect 28364 73276 28420 73278
rect 28252 73164 28308 73220
rect 28140 72380 28196 72436
rect 28028 70924 28084 70980
rect 28140 71596 28196 71652
rect 27804 70364 27860 70420
rect 28252 70924 28308 70980
rect 27916 69468 27972 69524
rect 27916 69298 27972 69300
rect 27916 69246 27918 69298
rect 27918 69246 27970 69298
rect 27970 69246 27972 69298
rect 27916 69244 27972 69246
rect 27692 68124 27748 68180
rect 24780 66556 24836 66612
rect 24668 65378 24724 65380
rect 24668 65326 24670 65378
rect 24670 65326 24722 65378
rect 24722 65326 24724 65378
rect 24668 65324 24724 65326
rect 24668 64594 24724 64596
rect 24668 64542 24670 64594
rect 24670 64542 24722 64594
rect 24722 64542 24724 64594
rect 24668 64540 24724 64542
rect 24668 63980 24724 64036
rect 24556 63138 24612 63140
rect 24556 63086 24558 63138
rect 24558 63086 24610 63138
rect 24610 63086 24612 63138
rect 24556 63084 24612 63086
rect 24332 62972 24388 63028
rect 23212 57650 23268 57652
rect 23212 57598 23214 57650
rect 23214 57598 23266 57650
rect 23266 57598 23268 57650
rect 23212 57596 23268 57598
rect 22764 57538 22820 57540
rect 22764 57486 22766 57538
rect 22766 57486 22818 57538
rect 22818 57486 22820 57538
rect 22764 57484 22820 57486
rect 23884 61346 23940 61348
rect 23884 61294 23886 61346
rect 23886 61294 23938 61346
rect 23938 61294 23940 61346
rect 23884 61292 23940 61294
rect 23660 61010 23716 61012
rect 23660 60958 23662 61010
rect 23662 60958 23714 61010
rect 23714 60958 23716 61010
rect 23660 60956 23716 60958
rect 23884 60002 23940 60004
rect 23884 59950 23886 60002
rect 23886 59950 23938 60002
rect 23938 59950 23940 60002
rect 23884 59948 23940 59950
rect 24220 60732 24276 60788
rect 24668 60732 24724 60788
rect 24668 59948 24724 60004
rect 23660 59052 23716 59108
rect 23548 57036 23604 57092
rect 22540 55410 22596 55412
rect 22540 55358 22542 55410
rect 22542 55358 22594 55410
rect 22594 55358 22596 55410
rect 22540 55356 22596 55358
rect 21980 53452 22036 53508
rect 21644 52780 21700 52836
rect 21420 52220 21476 52276
rect 21532 52668 21588 52724
rect 21308 52162 21364 52164
rect 21308 52110 21310 52162
rect 21310 52110 21362 52162
rect 21362 52110 21364 52162
rect 21308 52108 21364 52110
rect 21532 50876 21588 50932
rect 21420 49308 21476 49364
rect 21756 51996 21812 52052
rect 22092 52274 22148 52276
rect 22092 52222 22094 52274
rect 22094 52222 22146 52274
rect 22146 52222 22148 52274
rect 22092 52220 22148 52222
rect 23324 55356 23380 55412
rect 23436 54402 23492 54404
rect 23436 54350 23438 54402
rect 23438 54350 23490 54402
rect 23490 54350 23492 54402
rect 23436 54348 23492 54350
rect 23100 54236 23156 54292
rect 22316 53506 22372 53508
rect 22316 53454 22318 53506
rect 22318 53454 22370 53506
rect 22370 53454 22372 53506
rect 22316 53452 22372 53454
rect 22316 52332 22372 52388
rect 22204 51884 22260 51940
rect 22428 51324 22484 51380
rect 22540 50876 22596 50932
rect 22204 50764 22260 50820
rect 21980 50652 22036 50708
rect 21756 50594 21812 50596
rect 21756 50542 21758 50594
rect 21758 50542 21810 50594
rect 21810 50542 21812 50594
rect 21756 50540 21812 50542
rect 22764 52892 22820 52948
rect 22988 51378 23044 51380
rect 22988 51326 22990 51378
rect 22990 51326 23042 51378
rect 23042 51326 23044 51378
rect 22988 51324 23044 51326
rect 22316 48972 22372 49028
rect 21644 48748 21700 48804
rect 21980 48524 22036 48580
rect 21868 48242 21924 48244
rect 21868 48190 21870 48242
rect 21870 48190 21922 48242
rect 21922 48190 21924 48242
rect 21868 48188 21924 48190
rect 21532 47068 21588 47124
rect 21532 45052 21588 45108
rect 21308 44882 21364 44884
rect 21308 44830 21310 44882
rect 21310 44830 21362 44882
rect 21362 44830 21364 44882
rect 21308 44828 21364 44830
rect 21196 44604 21252 44660
rect 21532 44492 21588 44548
rect 21644 45164 21700 45220
rect 21308 44322 21364 44324
rect 21308 44270 21310 44322
rect 21310 44270 21362 44322
rect 21362 44270 21364 44322
rect 21308 44268 21364 44270
rect 21196 43820 21252 43876
rect 21308 42812 21364 42868
rect 21644 43484 21700 43540
rect 21756 46620 21812 46676
rect 22316 48524 22372 48580
rect 22092 48188 22148 48244
rect 22204 47068 22260 47124
rect 22092 46620 22148 46676
rect 21980 45836 22036 45892
rect 22092 45724 22148 45780
rect 21868 44380 21924 44436
rect 21980 45276 22036 45332
rect 21868 43314 21924 43316
rect 21868 43262 21870 43314
rect 21870 43262 21922 43314
rect 21922 43262 21924 43314
rect 21868 43260 21924 43262
rect 21868 42140 21924 42196
rect 21532 42028 21588 42084
rect 22204 45276 22260 45332
rect 22204 43484 22260 43540
rect 21644 41692 21700 41748
rect 21532 41244 21588 41300
rect 22092 41468 22148 41524
rect 21308 41186 21364 41188
rect 21308 41134 21310 41186
rect 21310 41134 21362 41186
rect 21362 41134 21364 41186
rect 21308 41132 21364 41134
rect 21868 41132 21924 41188
rect 21756 40348 21812 40404
rect 21644 39506 21700 39508
rect 21644 39454 21646 39506
rect 21646 39454 21698 39506
rect 21698 39454 21700 39506
rect 21644 39452 21700 39454
rect 21644 38668 21700 38724
rect 21644 37938 21700 37940
rect 21644 37886 21646 37938
rect 21646 37886 21698 37938
rect 21698 37886 21700 37938
rect 21644 37884 21700 37886
rect 21868 37938 21924 37940
rect 21868 37886 21870 37938
rect 21870 37886 21922 37938
rect 21922 37886 21924 37938
rect 21868 37884 21924 37886
rect 21756 37324 21812 37380
rect 21084 37212 21140 37268
rect 20860 35922 20916 35924
rect 20860 35870 20862 35922
rect 20862 35870 20914 35922
rect 20914 35870 20916 35922
rect 20860 35868 20916 35870
rect 21084 37042 21140 37044
rect 21084 36990 21086 37042
rect 21086 36990 21138 37042
rect 21138 36990 21140 37042
rect 21084 36988 21140 36990
rect 21532 36258 21588 36260
rect 21532 36206 21534 36258
rect 21534 36206 21586 36258
rect 21586 36206 21588 36258
rect 21532 36204 21588 36206
rect 20748 33516 20804 33572
rect 21868 33516 21924 33572
rect 21420 31836 21476 31892
rect 21308 31724 21364 31780
rect 21196 29426 21252 29428
rect 21196 29374 21198 29426
rect 21198 29374 21250 29426
rect 21250 29374 21252 29426
rect 21196 29372 21252 29374
rect 22092 40684 22148 40740
rect 24220 55020 24276 55076
rect 23548 54236 23604 54292
rect 24220 54290 24276 54292
rect 24220 54238 24222 54290
rect 24222 54238 24274 54290
rect 24274 54238 24276 54290
rect 24220 54236 24276 54238
rect 23436 53506 23492 53508
rect 23436 53454 23438 53506
rect 23438 53454 23490 53506
rect 23490 53454 23492 53506
rect 23436 53452 23492 53454
rect 23660 53116 23716 53172
rect 23436 52444 23492 52500
rect 23436 51884 23492 51940
rect 23548 51490 23604 51492
rect 23548 51438 23550 51490
rect 23550 51438 23602 51490
rect 23602 51438 23604 51490
rect 23548 51436 23604 51438
rect 23436 50428 23492 50484
rect 23100 50092 23156 50148
rect 22988 49698 23044 49700
rect 22988 49646 22990 49698
rect 22990 49646 23042 49698
rect 23042 49646 23044 49698
rect 22988 49644 23044 49646
rect 22652 48748 22708 48804
rect 23100 48914 23156 48916
rect 23100 48862 23102 48914
rect 23102 48862 23154 48914
rect 23154 48862 23156 48914
rect 23100 48860 23156 48862
rect 22764 48636 22820 48692
rect 22652 48242 22708 48244
rect 22652 48190 22654 48242
rect 22654 48190 22706 48242
rect 22706 48190 22708 48242
rect 22652 48188 22708 48190
rect 22540 44434 22596 44436
rect 22540 44382 22542 44434
rect 22542 44382 22594 44434
rect 22594 44382 22596 44434
rect 22540 44380 22596 44382
rect 22988 48412 23044 48468
rect 22876 45836 22932 45892
rect 22764 45778 22820 45780
rect 22764 45726 22766 45778
rect 22766 45726 22818 45778
rect 22818 45726 22820 45778
rect 22764 45724 22820 45726
rect 22652 43596 22708 43652
rect 22876 45500 22932 45556
rect 22540 43538 22596 43540
rect 22540 43486 22542 43538
rect 22542 43486 22594 43538
rect 22594 43486 22596 43538
rect 22540 43484 22596 43486
rect 22540 43036 22596 43092
rect 22428 41916 22484 41972
rect 22316 41132 22372 41188
rect 22316 40962 22372 40964
rect 22316 40910 22318 40962
rect 22318 40910 22370 40962
rect 22370 40910 22372 40962
rect 22316 40908 22372 40910
rect 22652 41580 22708 41636
rect 22428 40796 22484 40852
rect 22652 41410 22708 41412
rect 22652 41358 22654 41410
rect 22654 41358 22706 41410
rect 22706 41358 22708 41410
rect 22652 41356 22708 41358
rect 22652 40460 22708 40516
rect 22540 40290 22596 40292
rect 22540 40238 22542 40290
rect 22542 40238 22594 40290
rect 22594 40238 22596 40290
rect 22540 40236 22596 40238
rect 22204 40012 22260 40068
rect 23324 49922 23380 49924
rect 23324 49870 23326 49922
rect 23326 49870 23378 49922
rect 23378 49870 23380 49922
rect 23324 49868 23380 49870
rect 23548 49868 23604 49924
rect 23212 45388 23268 45444
rect 23324 46732 23380 46788
rect 23100 45276 23156 45332
rect 23884 52668 23940 52724
rect 23660 48636 23716 48692
rect 23772 52556 23828 52612
rect 23660 48300 23716 48356
rect 23660 47292 23716 47348
rect 23660 46786 23716 46788
rect 23660 46734 23662 46786
rect 23662 46734 23714 46786
rect 23714 46734 23716 46786
rect 23660 46732 23716 46734
rect 22876 44268 22932 44324
rect 23212 43708 23268 43764
rect 23212 43036 23268 43092
rect 23660 45948 23716 46004
rect 23436 45106 23492 45108
rect 23436 45054 23438 45106
rect 23438 45054 23490 45106
rect 23490 45054 23492 45106
rect 23436 45052 23492 45054
rect 23996 52108 24052 52164
rect 23996 50594 24052 50596
rect 23996 50542 23998 50594
rect 23998 50542 24050 50594
rect 24050 50542 24052 50594
rect 23996 50540 24052 50542
rect 23884 48242 23940 48244
rect 23884 48190 23886 48242
rect 23886 48190 23938 48242
rect 23938 48190 23940 48242
rect 23884 48188 23940 48190
rect 23884 45778 23940 45780
rect 23884 45726 23886 45778
rect 23886 45726 23938 45778
rect 23938 45726 23940 45778
rect 23884 45724 23940 45726
rect 23772 45164 23828 45220
rect 23660 45106 23716 45108
rect 23660 45054 23662 45106
rect 23662 45054 23714 45106
rect 23714 45054 23716 45106
rect 23660 45052 23716 45054
rect 23548 44492 23604 44548
rect 23772 43820 23828 43876
rect 23660 43650 23716 43652
rect 23660 43598 23662 43650
rect 23662 43598 23714 43650
rect 23714 43598 23716 43650
rect 23660 43596 23716 43598
rect 24220 49756 24276 49812
rect 24108 48860 24164 48916
rect 24220 46956 24276 47012
rect 24108 46620 24164 46676
rect 24220 45500 24276 45556
rect 24220 44882 24276 44884
rect 24220 44830 24222 44882
rect 24222 44830 24274 44882
rect 24274 44830 24276 44882
rect 24220 44828 24276 44830
rect 24108 44380 24164 44436
rect 24668 58434 24724 58436
rect 24668 58382 24670 58434
rect 24670 58382 24722 58434
rect 24722 58382 24724 58434
rect 24668 58380 24724 58382
rect 24556 56924 24612 56980
rect 24668 56812 24724 56868
rect 24556 55186 24612 55188
rect 24556 55134 24558 55186
rect 24558 55134 24610 55186
rect 24610 55134 24612 55186
rect 24556 55132 24612 55134
rect 24444 54402 24500 54404
rect 24444 54350 24446 54402
rect 24446 54350 24498 54402
rect 24498 54350 24500 54402
rect 24444 54348 24500 54350
rect 24668 52162 24724 52164
rect 24668 52110 24670 52162
rect 24670 52110 24722 52162
rect 24722 52110 24724 52162
rect 24668 52108 24724 52110
rect 24444 45836 24500 45892
rect 24556 50372 24612 50428
rect 24668 49308 24724 49364
rect 24668 48524 24724 48580
rect 26012 66668 26068 66724
rect 26012 66386 26068 66388
rect 26012 66334 26014 66386
rect 26014 66334 26066 66386
rect 26066 66334 26068 66386
rect 26012 66332 26068 66334
rect 27020 66332 27076 66388
rect 26348 66108 26404 66164
rect 24892 65436 24948 65492
rect 25228 65490 25284 65492
rect 25228 65438 25230 65490
rect 25230 65438 25282 65490
rect 25282 65438 25284 65490
rect 25228 65436 25284 65438
rect 25116 65324 25172 65380
rect 24892 65212 24948 65268
rect 25564 65324 25620 65380
rect 25340 65212 25396 65268
rect 26236 65378 26292 65380
rect 26236 65326 26238 65378
rect 26238 65326 26290 65378
rect 26290 65326 26292 65378
rect 26236 65324 26292 65326
rect 26684 65378 26740 65380
rect 26684 65326 26686 65378
rect 26686 65326 26738 65378
rect 26738 65326 26740 65378
rect 26684 65324 26740 65326
rect 25564 64092 25620 64148
rect 26236 64316 26292 64372
rect 26908 64482 26964 64484
rect 26908 64430 26910 64482
rect 26910 64430 26962 64482
rect 26962 64430 26964 64482
rect 26908 64428 26964 64430
rect 26460 63756 26516 63812
rect 25788 62972 25844 63028
rect 26684 63644 26740 63700
rect 28140 70418 28196 70420
rect 28140 70366 28142 70418
rect 28142 70366 28194 70418
rect 28194 70366 28196 70418
rect 28140 70364 28196 70366
rect 28140 70140 28196 70196
rect 29596 76466 29652 76468
rect 29596 76414 29598 76466
rect 29598 76414 29650 76466
rect 29650 76414 29652 76466
rect 29596 76412 29652 76414
rect 29148 75964 29204 76020
rect 29708 76188 29764 76244
rect 29260 75794 29316 75796
rect 29260 75742 29262 75794
rect 29262 75742 29314 75794
rect 29314 75742 29316 75794
rect 29260 75740 29316 75742
rect 29036 73330 29092 73332
rect 29036 73278 29038 73330
rect 29038 73278 29090 73330
rect 29090 73278 29092 73330
rect 29036 73276 29092 73278
rect 28924 71148 28980 71204
rect 29596 74844 29652 74900
rect 29260 74786 29316 74788
rect 29260 74734 29262 74786
rect 29262 74734 29314 74786
rect 29314 74734 29316 74786
rect 29260 74732 29316 74734
rect 29260 74060 29316 74116
rect 29260 73612 29316 73668
rect 29260 73052 29316 73108
rect 29932 80946 29988 80948
rect 29932 80894 29934 80946
rect 29934 80894 29986 80946
rect 29986 80894 29988 80946
rect 29932 80892 29988 80894
rect 30604 84588 30660 84644
rect 30492 83634 30548 83636
rect 30492 83582 30494 83634
rect 30494 83582 30546 83634
rect 30546 83582 30548 83634
rect 30492 83580 30548 83582
rect 30604 83132 30660 83188
rect 30380 82236 30436 82292
rect 30380 81340 30436 81396
rect 30268 79436 30324 79492
rect 30828 85202 30884 85204
rect 30828 85150 30830 85202
rect 30830 85150 30882 85202
rect 30882 85150 30884 85202
rect 30828 85148 30884 85150
rect 31052 84588 31108 84644
rect 30940 83298 30996 83300
rect 30940 83246 30942 83298
rect 30942 83246 30994 83298
rect 30994 83246 30996 83298
rect 30940 83244 30996 83246
rect 31276 85090 31332 85092
rect 31276 85038 31278 85090
rect 31278 85038 31330 85090
rect 31330 85038 31332 85090
rect 31276 85036 31332 85038
rect 31836 85708 31892 85764
rect 31948 85260 32004 85316
rect 35196 90186 35252 90188
rect 35196 90134 35198 90186
rect 35198 90134 35250 90186
rect 35250 90134 35252 90186
rect 35196 90132 35252 90134
rect 35300 90186 35356 90188
rect 35300 90134 35302 90186
rect 35302 90134 35354 90186
rect 35354 90134 35356 90186
rect 35300 90132 35356 90134
rect 35404 90186 35460 90188
rect 35404 90134 35406 90186
rect 35406 90134 35458 90186
rect 35458 90134 35460 90186
rect 35404 90132 35460 90134
rect 38220 91980 38276 92036
rect 38220 91420 38276 91476
rect 35196 88618 35252 88620
rect 35196 88566 35198 88618
rect 35198 88566 35250 88618
rect 35250 88566 35252 88618
rect 35196 88564 35252 88566
rect 35300 88618 35356 88620
rect 35300 88566 35302 88618
rect 35302 88566 35354 88618
rect 35354 88566 35356 88618
rect 35300 88564 35356 88566
rect 35404 88618 35460 88620
rect 35404 88566 35406 88618
rect 35406 88566 35458 88618
rect 35458 88566 35460 88618
rect 35404 88564 35460 88566
rect 35084 88002 35140 88004
rect 35084 87950 35086 88002
rect 35086 87950 35138 88002
rect 35138 87950 35140 88002
rect 35084 87948 35140 87950
rect 35532 88002 35588 88004
rect 35532 87950 35534 88002
rect 35534 87950 35586 88002
rect 35586 87950 35588 88002
rect 35532 87948 35588 87950
rect 32956 87442 33012 87444
rect 32956 87390 32958 87442
rect 32958 87390 33010 87442
rect 33010 87390 33012 87442
rect 32956 87388 33012 87390
rect 32508 85762 32564 85764
rect 32508 85710 32510 85762
rect 32510 85710 32562 85762
rect 32562 85710 32564 85762
rect 32508 85708 32564 85710
rect 32844 86044 32900 86100
rect 32508 85314 32564 85316
rect 32508 85262 32510 85314
rect 32510 85262 32562 85314
rect 32562 85262 32564 85314
rect 32508 85260 32564 85262
rect 33516 87330 33572 87332
rect 33516 87278 33518 87330
rect 33518 87278 33570 87330
rect 33570 87278 33572 87330
rect 33516 87276 33572 87278
rect 33628 86044 33684 86100
rect 32060 85036 32116 85092
rect 31500 84812 31556 84868
rect 31388 83410 31444 83412
rect 31388 83358 31390 83410
rect 31390 83358 31442 83410
rect 31442 83358 31444 83410
rect 31388 83356 31444 83358
rect 33292 85260 33348 85316
rect 33628 85036 33684 85092
rect 33852 85484 33908 85540
rect 32732 84866 32788 84868
rect 32732 84814 32734 84866
rect 32734 84814 32786 84866
rect 32786 84814 32788 84866
rect 32732 84812 32788 84814
rect 34972 87276 35028 87332
rect 35196 87050 35252 87052
rect 35196 86998 35198 87050
rect 35198 86998 35250 87050
rect 35250 86998 35252 87050
rect 35196 86996 35252 86998
rect 35300 87050 35356 87052
rect 35300 86998 35302 87050
rect 35302 86998 35354 87050
rect 35354 86998 35356 87050
rect 35300 86996 35356 86998
rect 35404 87050 35460 87052
rect 35404 86998 35406 87050
rect 35406 86998 35458 87050
rect 35458 86998 35460 87050
rect 35404 86996 35460 86998
rect 34524 85484 34580 85540
rect 34748 85148 34804 85204
rect 34412 85090 34468 85092
rect 34412 85038 34414 85090
rect 34414 85038 34466 85090
rect 34466 85038 34468 85090
rect 34412 85036 34468 85038
rect 35196 85482 35252 85484
rect 35196 85430 35198 85482
rect 35198 85430 35250 85482
rect 35250 85430 35252 85482
rect 35196 85428 35252 85430
rect 35300 85482 35356 85484
rect 35300 85430 35302 85482
rect 35302 85430 35354 85482
rect 35354 85430 35356 85482
rect 35300 85428 35356 85430
rect 35404 85482 35460 85484
rect 35404 85430 35406 85482
rect 35406 85430 35458 85482
rect 35458 85430 35460 85482
rect 35404 85428 35460 85430
rect 35084 85036 35140 85092
rect 33964 84700 34020 84756
rect 31948 84028 32004 84084
rect 31612 82626 31668 82628
rect 31612 82574 31614 82626
rect 31614 82574 31666 82626
rect 31666 82574 31668 82626
rect 31612 82572 31668 82574
rect 31276 81730 31332 81732
rect 31276 81678 31278 81730
rect 31278 81678 31330 81730
rect 31330 81678 31332 81730
rect 31276 81676 31332 81678
rect 30492 79212 30548 79268
rect 30044 78764 30100 78820
rect 30492 78764 30548 78820
rect 30604 78876 30660 78932
rect 33180 82626 33236 82628
rect 33180 82574 33182 82626
rect 33182 82574 33234 82626
rect 33234 82574 33236 82626
rect 33180 82572 33236 82574
rect 31612 81394 31668 81396
rect 31612 81342 31614 81394
rect 31614 81342 31666 81394
rect 31666 81342 31668 81394
rect 31612 81340 31668 81342
rect 30156 78540 30212 78596
rect 30492 78594 30548 78596
rect 30492 78542 30494 78594
rect 30494 78542 30546 78594
rect 30546 78542 30548 78594
rect 30492 78540 30548 78542
rect 32956 81954 33012 81956
rect 32956 81902 32958 81954
rect 32958 81902 33010 81954
rect 33010 81902 33012 81954
rect 32956 81900 33012 81902
rect 34524 84028 34580 84084
rect 34972 84812 35028 84868
rect 34748 84476 34804 84532
rect 33852 82348 33908 82404
rect 34188 81900 34244 81956
rect 30940 79378 30996 79380
rect 30940 79326 30942 79378
rect 30942 79326 30994 79378
rect 30994 79326 30996 79378
rect 30940 79324 30996 79326
rect 31500 78652 31556 78708
rect 30268 77644 30324 77700
rect 30380 77980 30436 78036
rect 30380 76972 30436 77028
rect 30156 76748 30212 76804
rect 29820 75516 29876 75572
rect 29820 74226 29876 74228
rect 29820 74174 29822 74226
rect 29822 74174 29874 74226
rect 29874 74174 29876 74226
rect 29820 74172 29876 74174
rect 29820 73442 29876 73444
rect 29820 73390 29822 73442
rect 29822 73390 29874 73442
rect 29874 73390 29876 73442
rect 29820 73388 29876 73390
rect 29820 72658 29876 72660
rect 29820 72606 29822 72658
rect 29822 72606 29874 72658
rect 29874 72606 29876 72658
rect 29820 72604 29876 72606
rect 29372 71484 29428 71540
rect 29372 70978 29428 70980
rect 29372 70926 29374 70978
rect 29374 70926 29426 70978
rect 29426 70926 29428 70978
rect 29372 70924 29428 70926
rect 29148 70364 29204 70420
rect 28476 69916 28532 69972
rect 28364 69580 28420 69636
rect 29260 69692 29316 69748
rect 30156 75740 30212 75796
rect 30044 75458 30100 75460
rect 30044 75406 30046 75458
rect 30046 75406 30098 75458
rect 30098 75406 30100 75458
rect 30044 75404 30100 75406
rect 30492 76578 30548 76580
rect 30492 76526 30494 76578
rect 30494 76526 30546 76578
rect 30546 76526 30548 76578
rect 30492 76524 30548 76526
rect 30380 76188 30436 76244
rect 30716 76188 30772 76244
rect 30828 77756 30884 77812
rect 32396 78930 32452 78932
rect 32396 78878 32398 78930
rect 32398 78878 32450 78930
rect 32450 78878 32452 78930
rect 32396 78876 32452 78878
rect 31724 78316 31780 78372
rect 31836 78540 31892 78596
rect 31052 77532 31108 77588
rect 31276 78034 31332 78036
rect 31276 77982 31278 78034
rect 31278 77982 31330 78034
rect 31330 77982 31332 78034
rect 31276 77980 31332 77982
rect 31500 78034 31556 78036
rect 31500 77982 31502 78034
rect 31502 77982 31554 78034
rect 31554 77982 31556 78034
rect 31500 77980 31556 77982
rect 32060 78652 32116 78708
rect 30940 77420 30996 77476
rect 31164 77308 31220 77364
rect 31164 76860 31220 76916
rect 31276 76972 31332 77028
rect 30380 75740 30436 75796
rect 31052 75964 31108 76020
rect 30604 75682 30660 75684
rect 30604 75630 30606 75682
rect 30606 75630 30658 75682
rect 30658 75630 30660 75682
rect 30604 75628 30660 75630
rect 30940 75570 30996 75572
rect 30940 75518 30942 75570
rect 30942 75518 30994 75570
rect 30994 75518 30996 75570
rect 30940 75516 30996 75518
rect 31612 77532 31668 77588
rect 31500 77138 31556 77140
rect 31500 77086 31502 77138
rect 31502 77086 31554 77138
rect 31554 77086 31556 77138
rect 31500 77084 31556 77086
rect 31724 76748 31780 76804
rect 32732 78540 32788 78596
rect 32396 78316 32452 78372
rect 32172 78258 32228 78260
rect 32172 78206 32174 78258
rect 32174 78206 32226 78258
rect 32226 78206 32228 78258
rect 32172 78204 32228 78206
rect 32060 77420 32116 77476
rect 32396 77308 32452 77364
rect 32172 77250 32228 77252
rect 32172 77198 32174 77250
rect 32174 77198 32226 77250
rect 32226 77198 32228 77250
rect 32172 77196 32228 77198
rect 32060 76860 32116 76916
rect 32396 76860 32452 76916
rect 32508 76748 32564 76804
rect 32844 77980 32900 78036
rect 35420 84700 35476 84756
rect 35308 84476 35364 84532
rect 36204 87948 36260 88004
rect 35980 85148 36036 85204
rect 35868 85090 35924 85092
rect 35868 85038 35870 85090
rect 35870 85038 35922 85090
rect 35922 85038 35924 85090
rect 35868 85036 35924 85038
rect 34860 83522 34916 83524
rect 34860 83470 34862 83522
rect 34862 83470 34914 83522
rect 34914 83470 34916 83522
rect 34860 83468 34916 83470
rect 34636 83298 34692 83300
rect 34636 83246 34638 83298
rect 34638 83246 34690 83298
rect 34690 83246 34692 83298
rect 34636 83244 34692 83246
rect 35196 83914 35252 83916
rect 35196 83862 35198 83914
rect 35198 83862 35250 83914
rect 35250 83862 35252 83914
rect 35196 83860 35252 83862
rect 35300 83914 35356 83916
rect 35300 83862 35302 83914
rect 35302 83862 35354 83914
rect 35354 83862 35356 83914
rect 35300 83860 35356 83862
rect 35404 83914 35460 83916
rect 35404 83862 35406 83914
rect 35406 83862 35458 83914
rect 35458 83862 35460 83914
rect 35404 83860 35460 83862
rect 35644 83916 35700 83972
rect 36092 83692 36148 83748
rect 35980 83522 36036 83524
rect 35980 83470 35982 83522
rect 35982 83470 36034 83522
rect 36034 83470 36036 83522
rect 35980 83468 36036 83470
rect 36204 83410 36260 83412
rect 36204 83358 36206 83410
rect 36206 83358 36258 83410
rect 36258 83358 36260 83410
rect 36204 83356 36260 83358
rect 36876 85148 36932 85204
rect 38332 84924 38388 84980
rect 37660 84866 37716 84868
rect 37660 84814 37662 84866
rect 37662 84814 37714 84866
rect 37714 84814 37716 84866
rect 37660 84812 37716 84814
rect 36540 84588 36596 84644
rect 36428 84476 36484 84532
rect 37100 84476 37156 84532
rect 37212 84028 37268 84084
rect 37100 83746 37156 83748
rect 37100 83694 37102 83746
rect 37102 83694 37154 83746
rect 37154 83694 37156 83746
rect 37100 83692 37156 83694
rect 36988 83410 37044 83412
rect 36988 83358 36990 83410
rect 36990 83358 37042 83410
rect 37042 83358 37044 83410
rect 36988 83356 37044 83358
rect 37660 83916 37716 83972
rect 37548 83298 37604 83300
rect 37548 83246 37550 83298
rect 37550 83246 37602 83298
rect 37602 83246 37604 83298
rect 37548 83244 37604 83246
rect 34524 82572 34580 82628
rect 38108 84028 38164 84084
rect 38220 83916 38276 83972
rect 34636 82348 34692 82404
rect 35196 82346 35252 82348
rect 35196 82294 35198 82346
rect 35198 82294 35250 82346
rect 35250 82294 35252 82346
rect 35196 82292 35252 82294
rect 35300 82346 35356 82348
rect 35300 82294 35302 82346
rect 35302 82294 35354 82346
rect 35354 82294 35356 82346
rect 35300 82292 35356 82294
rect 35404 82346 35460 82348
rect 35404 82294 35406 82346
rect 35406 82294 35458 82346
rect 35458 82294 35460 82346
rect 35404 82292 35460 82294
rect 35196 81954 35252 81956
rect 35196 81902 35198 81954
rect 35198 81902 35250 81954
rect 35250 81902 35252 81954
rect 35196 81900 35252 81902
rect 36204 81954 36260 81956
rect 36204 81902 36206 81954
rect 36206 81902 36258 81954
rect 36258 81902 36260 81954
rect 36204 81900 36260 81902
rect 37884 81900 37940 81956
rect 34412 81676 34468 81732
rect 35308 81730 35364 81732
rect 35308 81678 35310 81730
rect 35310 81678 35362 81730
rect 35362 81678 35364 81730
rect 35308 81676 35364 81678
rect 34188 80668 34244 80724
rect 35196 80778 35252 80780
rect 35196 80726 35198 80778
rect 35198 80726 35250 80778
rect 35250 80726 35252 80778
rect 35196 80724 35252 80726
rect 35300 80778 35356 80780
rect 35300 80726 35302 80778
rect 35302 80726 35354 80778
rect 35354 80726 35356 80778
rect 35300 80724 35356 80726
rect 35404 80778 35460 80780
rect 35404 80726 35406 80778
rect 35406 80726 35458 80778
rect 35458 80726 35460 80778
rect 35404 80724 35460 80726
rect 33292 78930 33348 78932
rect 33292 78878 33294 78930
rect 33294 78878 33346 78930
rect 33346 78878 33348 78930
rect 33292 78876 33348 78878
rect 35196 79210 35252 79212
rect 35196 79158 35198 79210
rect 35198 79158 35250 79210
rect 35250 79158 35252 79210
rect 35196 79156 35252 79158
rect 35300 79210 35356 79212
rect 35300 79158 35302 79210
rect 35302 79158 35354 79210
rect 35354 79158 35356 79210
rect 35300 79156 35356 79158
rect 35404 79210 35460 79212
rect 35404 79158 35406 79210
rect 35406 79158 35458 79210
rect 35458 79158 35460 79210
rect 35404 79156 35460 79158
rect 34412 77980 34468 78036
rect 34076 77922 34132 77924
rect 34076 77870 34078 77922
rect 34078 77870 34130 77922
rect 34130 77870 34132 77922
rect 34076 77868 34132 77870
rect 33180 77644 33236 77700
rect 33068 77420 33124 77476
rect 34860 78594 34916 78596
rect 34860 78542 34862 78594
rect 34862 78542 34914 78594
rect 34914 78542 34916 78594
rect 34860 78540 34916 78542
rect 35308 78258 35364 78260
rect 35308 78206 35310 78258
rect 35310 78206 35362 78258
rect 35362 78206 35364 78258
rect 35308 78204 35364 78206
rect 34636 78146 34692 78148
rect 34636 78094 34638 78146
rect 34638 78094 34690 78146
rect 34690 78094 34692 78146
rect 34636 78092 34692 78094
rect 35084 78034 35140 78036
rect 35084 77982 35086 78034
rect 35086 77982 35138 78034
rect 35138 77982 35140 78034
rect 35084 77980 35140 77982
rect 35532 78034 35588 78036
rect 35532 77982 35534 78034
rect 35534 77982 35586 78034
rect 35586 77982 35588 78034
rect 35532 77980 35588 77982
rect 35084 77756 35140 77812
rect 34524 77532 34580 77588
rect 34412 77196 34468 77252
rect 33292 77138 33348 77140
rect 33292 77086 33294 77138
rect 33294 77086 33346 77138
rect 33346 77086 33348 77138
rect 33292 77084 33348 77086
rect 33180 76860 33236 76916
rect 34188 77138 34244 77140
rect 34188 77086 34190 77138
rect 34190 77086 34242 77138
rect 34242 77086 34244 77138
rect 34188 77084 34244 77086
rect 34300 77026 34356 77028
rect 34300 76974 34302 77026
rect 34302 76974 34354 77026
rect 34354 76974 34356 77026
rect 34300 76972 34356 76974
rect 33628 76860 33684 76916
rect 32956 76524 33012 76580
rect 32284 75740 32340 75796
rect 33516 76466 33572 76468
rect 33516 76414 33518 76466
rect 33518 76414 33570 76466
rect 33570 76414 33572 76466
rect 33516 76412 33572 76414
rect 31948 75682 32004 75684
rect 31948 75630 31950 75682
rect 31950 75630 32002 75682
rect 32002 75630 32004 75682
rect 31948 75628 32004 75630
rect 30492 75180 30548 75236
rect 30604 74898 30660 74900
rect 30604 74846 30606 74898
rect 30606 74846 30658 74898
rect 30658 74846 30660 74898
rect 30604 74844 30660 74846
rect 30268 74226 30324 74228
rect 30268 74174 30270 74226
rect 30270 74174 30322 74226
rect 30322 74174 30324 74226
rect 30268 74172 30324 74174
rect 29820 70588 29876 70644
rect 29932 71036 29988 71092
rect 29708 70140 29764 70196
rect 28252 69244 28308 69300
rect 28476 68460 28532 68516
rect 28588 67900 28644 67956
rect 29596 69580 29652 69636
rect 29372 69468 29428 69524
rect 29148 69410 29204 69412
rect 29148 69358 29150 69410
rect 29150 69358 29202 69410
rect 29202 69358 29204 69410
rect 29148 69356 29204 69358
rect 29036 68514 29092 68516
rect 29036 68462 29038 68514
rect 29038 68462 29090 68514
rect 29090 68462 29092 68514
rect 29036 68460 29092 68462
rect 29260 68460 29316 68516
rect 29708 68460 29764 68516
rect 29596 68236 29652 68292
rect 29596 67116 29652 67172
rect 29148 67058 29204 67060
rect 29148 67006 29150 67058
rect 29150 67006 29202 67058
rect 29202 67006 29204 67058
rect 29148 67004 29204 67006
rect 29484 66780 29540 66836
rect 29708 68124 29764 68180
rect 30268 71484 30324 71540
rect 30268 70812 30324 70868
rect 30716 74226 30772 74228
rect 30716 74174 30718 74226
rect 30718 74174 30770 74226
rect 30770 74174 30772 74226
rect 30716 74172 30772 74174
rect 30492 73554 30548 73556
rect 30492 73502 30494 73554
rect 30494 73502 30546 73554
rect 30546 73502 30548 73554
rect 30492 73500 30548 73502
rect 30380 70588 30436 70644
rect 29820 67900 29876 67956
rect 30044 68684 30100 68740
rect 30044 68514 30100 68516
rect 30044 68462 30046 68514
rect 30046 68462 30098 68514
rect 30098 68462 30100 68514
rect 30044 68460 30100 68462
rect 30604 70924 30660 70980
rect 30716 70812 30772 70868
rect 31612 75404 31668 75460
rect 31500 74172 31556 74228
rect 31500 73948 31556 74004
rect 31052 73442 31108 73444
rect 31052 73390 31054 73442
rect 31054 73390 31106 73442
rect 31106 73390 31108 73442
rect 31052 73388 31108 73390
rect 31276 72546 31332 72548
rect 31276 72494 31278 72546
rect 31278 72494 31330 72546
rect 31330 72494 31332 72546
rect 31276 72492 31332 72494
rect 30492 69468 30548 69524
rect 30716 70140 30772 70196
rect 30380 68908 30436 68964
rect 31052 70866 31108 70868
rect 31052 70814 31054 70866
rect 31054 70814 31106 70866
rect 31106 70814 31108 70866
rect 31052 70812 31108 70814
rect 31052 70588 31108 70644
rect 30044 66946 30100 66948
rect 30044 66894 30046 66946
rect 30046 66894 30098 66946
rect 30098 66894 30100 66946
rect 30044 66892 30100 66894
rect 28812 65996 28868 66052
rect 28588 64930 28644 64932
rect 28588 64878 28590 64930
rect 28590 64878 28642 64930
rect 28642 64878 28644 64930
rect 28588 64876 28644 64878
rect 27804 64594 27860 64596
rect 27804 64542 27806 64594
rect 27806 64542 27858 64594
rect 27858 64542 27860 64594
rect 27804 64540 27860 64542
rect 30716 68572 30772 68628
rect 30492 67170 30548 67172
rect 30492 67118 30494 67170
rect 30494 67118 30546 67170
rect 30546 67118 30548 67170
rect 30492 67116 30548 67118
rect 29708 65996 29764 66052
rect 29484 64876 29540 64932
rect 29596 65436 29652 65492
rect 29260 64594 29316 64596
rect 29260 64542 29262 64594
rect 29262 64542 29314 64594
rect 29314 64542 29316 64594
rect 29260 64540 29316 64542
rect 29484 64482 29540 64484
rect 29484 64430 29486 64482
rect 29486 64430 29538 64482
rect 29538 64430 29540 64482
rect 29484 64428 29540 64430
rect 28140 64092 28196 64148
rect 27132 64034 27188 64036
rect 27132 63982 27134 64034
rect 27134 63982 27186 64034
rect 27186 63982 27188 64034
rect 27132 63980 27188 63982
rect 27804 63980 27860 64036
rect 27356 63756 27412 63812
rect 27020 63084 27076 63140
rect 26684 62524 26740 62580
rect 28812 64092 28868 64148
rect 29148 64092 29204 64148
rect 29484 64092 29540 64148
rect 29260 64034 29316 64036
rect 29260 63982 29262 64034
rect 29262 63982 29314 64034
rect 29314 63982 29316 64034
rect 29260 63980 29316 63982
rect 30380 65996 30436 66052
rect 30044 64482 30100 64484
rect 30044 64430 30046 64482
rect 30046 64430 30098 64482
rect 30098 64430 30100 64482
rect 30044 64428 30100 64430
rect 28924 63922 28980 63924
rect 28924 63870 28926 63922
rect 28926 63870 28978 63922
rect 28978 63870 28980 63922
rect 28924 63868 28980 63870
rect 28252 63644 28308 63700
rect 27692 60956 27748 61012
rect 24892 58380 24948 58436
rect 24892 57036 24948 57092
rect 24892 56252 24948 56308
rect 27468 60786 27524 60788
rect 27468 60734 27470 60786
rect 27470 60734 27522 60786
rect 27522 60734 27524 60786
rect 27468 60732 27524 60734
rect 25676 60002 25732 60004
rect 25676 59950 25678 60002
rect 25678 59950 25730 60002
rect 25730 59950 25732 60002
rect 25676 59948 25732 59950
rect 26012 59948 26068 60004
rect 25676 59164 25732 59220
rect 25340 56306 25396 56308
rect 25340 56254 25342 56306
rect 25342 56254 25394 56306
rect 25394 56254 25396 56306
rect 25340 56252 25396 56254
rect 25004 55020 25060 55076
rect 24892 49138 24948 49140
rect 24892 49086 24894 49138
rect 24894 49086 24946 49138
rect 24946 49086 24948 49138
rect 24892 49084 24948 49086
rect 25116 51884 25172 51940
rect 25340 51996 25396 52052
rect 26348 60002 26404 60004
rect 26348 59950 26350 60002
rect 26350 59950 26402 60002
rect 26402 59950 26404 60002
rect 26348 59948 26404 59950
rect 27692 59890 27748 59892
rect 27692 59838 27694 59890
rect 27694 59838 27746 59890
rect 27746 59838 27748 59890
rect 27692 59836 27748 59838
rect 27804 63138 27860 63140
rect 27804 63086 27806 63138
rect 27806 63086 27858 63138
rect 27858 63086 27860 63138
rect 27804 63084 27860 63086
rect 28476 62972 28532 63028
rect 29484 63644 29540 63700
rect 29260 63026 29316 63028
rect 29260 62974 29262 63026
rect 29262 62974 29314 63026
rect 29314 62974 29316 63026
rect 29260 62972 29316 62974
rect 29596 63026 29652 63028
rect 29596 62974 29598 63026
rect 29598 62974 29650 63026
rect 29650 62974 29652 63026
rect 29596 62972 29652 62974
rect 29932 63922 29988 63924
rect 29932 63870 29934 63922
rect 29934 63870 29986 63922
rect 29986 63870 29988 63922
rect 29932 63868 29988 63870
rect 29484 62354 29540 62356
rect 29484 62302 29486 62354
rect 29486 62302 29538 62354
rect 29538 62302 29540 62354
rect 29484 62300 29540 62302
rect 28588 61964 28644 62020
rect 26012 53900 26068 53956
rect 26348 59052 26404 59108
rect 25900 53340 25956 53396
rect 25228 49810 25284 49812
rect 25228 49758 25230 49810
rect 25230 49758 25282 49810
rect 25282 49758 25284 49810
rect 25228 49756 25284 49758
rect 25340 49308 25396 49364
rect 25228 48748 25284 48804
rect 25564 49308 25620 49364
rect 26124 51212 26180 51268
rect 26124 50652 26180 50708
rect 25900 49084 25956 49140
rect 25788 48636 25844 48692
rect 24668 46674 24724 46676
rect 24668 46622 24670 46674
rect 24670 46622 24722 46674
rect 24722 46622 24724 46674
rect 24668 46620 24724 46622
rect 23436 43484 23492 43540
rect 22988 41468 23044 41524
rect 22876 41298 22932 41300
rect 22876 41246 22878 41298
rect 22878 41246 22930 41298
rect 22930 41246 22932 41298
rect 22876 41244 22932 41246
rect 22876 40908 22932 40964
rect 22988 40460 23044 40516
rect 22204 39394 22260 39396
rect 22204 39342 22206 39394
rect 22206 39342 22258 39394
rect 22258 39342 22260 39394
rect 22204 39340 22260 39342
rect 22092 39004 22148 39060
rect 22204 38780 22260 38836
rect 23324 41692 23380 41748
rect 23772 42476 23828 42532
rect 23548 42252 23604 42308
rect 24108 43484 24164 43540
rect 25228 46844 25284 46900
rect 26124 48130 26180 48132
rect 26124 48078 26126 48130
rect 26126 48078 26178 48130
rect 26178 48078 26180 48130
rect 26124 48076 26180 48078
rect 25340 46732 25396 46788
rect 25564 46562 25620 46564
rect 25564 46510 25566 46562
rect 25566 46510 25618 46562
rect 25618 46510 25620 46562
rect 25564 46508 25620 46510
rect 25452 46060 25508 46116
rect 25676 45836 25732 45892
rect 26236 46284 26292 46340
rect 25788 45948 25844 46004
rect 24780 45164 24836 45220
rect 24668 45052 24724 45108
rect 24892 44828 24948 44884
rect 23996 41916 24052 41972
rect 23548 41692 23604 41748
rect 23212 41132 23268 41188
rect 22764 38780 22820 38836
rect 22652 38556 22708 38612
rect 22316 38444 22372 38500
rect 22540 38332 22596 38388
rect 22428 37378 22484 37380
rect 22428 37326 22430 37378
rect 22430 37326 22482 37378
rect 22482 37326 22484 37378
rect 22428 37324 22484 37326
rect 22428 36316 22484 36372
rect 22204 36258 22260 36260
rect 22204 36206 22206 36258
rect 22206 36206 22258 36258
rect 22258 36206 22260 36258
rect 22204 36204 22260 36206
rect 22204 35980 22260 36036
rect 22316 35308 22372 35364
rect 22428 33628 22484 33684
rect 21980 31724 22036 31780
rect 22428 29932 22484 29988
rect 21756 29426 21812 29428
rect 21756 29374 21758 29426
rect 21758 29374 21810 29426
rect 21810 29374 21812 29426
rect 21756 29372 21812 29374
rect 21644 28140 21700 28196
rect 18956 18396 19012 18452
rect 19628 23884 19684 23940
rect 19628 23548 19684 23604
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19964 22540 20020 22596
rect 19628 22258 19684 22260
rect 19628 22206 19630 22258
rect 19630 22206 19682 22258
rect 19682 22206 19684 22258
rect 19628 22204 19684 22206
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 19516 21756 19572 21812
rect 19068 16770 19124 16772
rect 19068 16718 19070 16770
rect 19070 16718 19122 16770
rect 19122 16718 19124 16770
rect 19068 16716 19124 16718
rect 19068 16492 19124 16548
rect 18956 15596 19012 15652
rect 17948 13634 18004 13636
rect 17948 13582 17950 13634
rect 17950 13582 18002 13634
rect 18002 13582 18004 13634
rect 17948 13580 18004 13582
rect 18284 13074 18340 13076
rect 18284 13022 18286 13074
rect 18286 13022 18338 13074
rect 18338 13022 18340 13074
rect 18284 13020 18340 13022
rect 17388 12460 17444 12516
rect 17500 12178 17556 12180
rect 17500 12126 17502 12178
rect 17502 12126 17554 12178
rect 17554 12126 17556 12178
rect 17500 12124 17556 12126
rect 17388 11900 17444 11956
rect 17836 11900 17892 11956
rect 18060 12178 18116 12180
rect 18060 12126 18062 12178
rect 18062 12126 18114 12178
rect 18114 12126 18116 12178
rect 18060 12124 18116 12126
rect 17948 11788 18004 11844
rect 17724 10780 17780 10836
rect 17836 11452 17892 11508
rect 16828 10444 16884 10500
rect 17500 10498 17556 10500
rect 17500 10446 17502 10498
rect 17502 10446 17554 10498
rect 17554 10446 17556 10498
rect 17500 10444 17556 10446
rect 17164 9884 17220 9940
rect 17724 9996 17780 10052
rect 17500 9772 17556 9828
rect 18620 13634 18676 13636
rect 18620 13582 18622 13634
rect 18622 13582 18674 13634
rect 18674 13582 18676 13634
rect 18620 13580 18676 13582
rect 18620 13132 18676 13188
rect 18956 15036 19012 15092
rect 18844 13020 18900 13076
rect 18956 12348 19012 12404
rect 19404 15986 19460 15988
rect 19404 15934 19406 15986
rect 19406 15934 19458 15986
rect 19458 15934 19460 15986
rect 19404 15932 19460 15934
rect 19292 15596 19348 15652
rect 19292 15426 19348 15428
rect 19292 15374 19294 15426
rect 19294 15374 19346 15426
rect 19346 15374 19348 15426
rect 19292 15372 19348 15374
rect 19404 15202 19460 15204
rect 19404 15150 19406 15202
rect 19406 15150 19458 15202
rect 19458 15150 19460 15202
rect 19404 15148 19460 15150
rect 19180 15036 19236 15092
rect 19180 12348 19236 12404
rect 19068 12290 19124 12292
rect 19068 12238 19070 12290
rect 19070 12238 19122 12290
rect 19122 12238 19124 12290
rect 19068 12236 19124 12238
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 20076 18620 20132 18676
rect 19964 18396 20020 18452
rect 19740 18284 19796 18340
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19628 16268 19684 16324
rect 20412 23660 20468 23716
rect 20300 23324 20356 23380
rect 22764 37436 22820 37492
rect 23100 38162 23156 38164
rect 23100 38110 23102 38162
rect 23102 38110 23154 38162
rect 23154 38110 23156 38162
rect 23100 38108 23156 38110
rect 23100 37884 23156 37940
rect 22988 36428 23044 36484
rect 22988 36204 23044 36260
rect 22988 34076 23044 34132
rect 23884 41468 23940 41524
rect 23436 40290 23492 40292
rect 23436 40238 23438 40290
rect 23438 40238 23490 40290
rect 23490 40238 23492 40290
rect 23436 40236 23492 40238
rect 23324 38946 23380 38948
rect 23324 38894 23326 38946
rect 23326 38894 23378 38946
rect 23378 38894 23380 38946
rect 23324 38892 23380 38894
rect 23436 38332 23492 38388
rect 23324 33628 23380 33684
rect 23772 41074 23828 41076
rect 23772 41022 23774 41074
rect 23774 41022 23826 41074
rect 23826 41022 23828 41074
rect 23772 41020 23828 41022
rect 23884 40684 23940 40740
rect 23660 40348 23716 40404
rect 24108 41244 24164 41300
rect 24332 42252 24388 42308
rect 24668 42588 24724 42644
rect 24332 42028 24388 42084
rect 24220 41580 24276 41636
rect 24108 41020 24164 41076
rect 24444 41132 24500 41188
rect 24220 40796 24276 40852
rect 24220 40626 24276 40628
rect 24220 40574 24222 40626
rect 24222 40574 24274 40626
rect 24274 40574 24276 40626
rect 24220 40572 24276 40574
rect 25564 44156 25620 44212
rect 26012 45218 26068 45220
rect 26012 45166 26014 45218
rect 26014 45166 26066 45218
rect 26066 45166 26068 45218
rect 26012 45164 26068 45166
rect 25788 44828 25844 44884
rect 25564 43820 25620 43876
rect 25564 43426 25620 43428
rect 25564 43374 25566 43426
rect 25566 43374 25618 43426
rect 25618 43374 25620 43426
rect 25564 43372 25620 43374
rect 25004 41916 25060 41972
rect 24780 41468 24836 41524
rect 24668 40626 24724 40628
rect 24668 40574 24670 40626
rect 24670 40574 24722 40626
rect 24722 40574 24724 40626
rect 24668 40572 24724 40574
rect 23996 39900 24052 39956
rect 24668 39900 24724 39956
rect 24108 39842 24164 39844
rect 24108 39790 24110 39842
rect 24110 39790 24162 39842
rect 24162 39790 24164 39842
rect 24108 39788 24164 39790
rect 23660 39676 23716 39732
rect 23660 38108 23716 38164
rect 24108 39340 24164 39396
rect 24444 39730 24500 39732
rect 24444 39678 24446 39730
rect 24446 39678 24498 39730
rect 24498 39678 24500 39730
rect 24444 39676 24500 39678
rect 24444 39340 24500 39396
rect 24444 39004 24500 39060
rect 23996 37436 24052 37492
rect 24108 38108 24164 38164
rect 23548 36258 23604 36260
rect 23548 36206 23550 36258
rect 23550 36206 23602 36258
rect 23602 36206 23604 36258
rect 23548 36204 23604 36206
rect 23548 34130 23604 34132
rect 23548 34078 23550 34130
rect 23550 34078 23602 34130
rect 23602 34078 23604 34130
rect 23548 34076 23604 34078
rect 23996 36482 24052 36484
rect 23996 36430 23998 36482
rect 23998 36430 24050 36482
rect 24050 36430 24052 36482
rect 23996 36428 24052 36430
rect 23548 33628 23604 33684
rect 23772 35308 23828 35364
rect 24892 39506 24948 39508
rect 24892 39454 24894 39506
rect 24894 39454 24946 39506
rect 24946 39454 24948 39506
rect 24892 39452 24948 39454
rect 28476 61516 28532 61572
rect 28252 60898 28308 60900
rect 28252 60846 28254 60898
rect 28254 60846 28306 60898
rect 28306 60846 28308 60898
rect 28252 60844 28308 60846
rect 27916 60786 27972 60788
rect 27916 60734 27918 60786
rect 27918 60734 27970 60786
rect 27970 60734 27972 60786
rect 27916 60732 27972 60734
rect 28364 60732 28420 60788
rect 29260 61852 29316 61908
rect 29820 62578 29876 62580
rect 29820 62526 29822 62578
rect 29822 62526 29874 62578
rect 29874 62526 29876 62578
rect 29820 62524 29876 62526
rect 29932 61964 29988 62020
rect 29148 61404 29204 61460
rect 27692 58322 27748 58324
rect 27692 58270 27694 58322
rect 27694 58270 27746 58322
rect 27746 58270 27748 58322
rect 27692 58268 27748 58270
rect 26684 57036 26740 57092
rect 27468 56978 27524 56980
rect 27468 56926 27470 56978
rect 27470 56926 27522 56978
rect 27522 56926 27524 56978
rect 27468 56924 27524 56926
rect 26796 53900 26852 53956
rect 26796 53340 26852 53396
rect 28028 58210 28084 58212
rect 28028 58158 28030 58210
rect 28030 58158 28082 58210
rect 28082 58158 28084 58210
rect 28028 58156 28084 58158
rect 28028 57596 28084 57652
rect 28700 59778 28756 59780
rect 28700 59726 28702 59778
rect 28702 59726 28754 59778
rect 28754 59726 28756 59778
rect 28700 59724 28756 59726
rect 28252 58268 28308 58324
rect 28140 57036 28196 57092
rect 28140 56252 28196 56308
rect 27020 54236 27076 54292
rect 27692 54290 27748 54292
rect 27692 54238 27694 54290
rect 27694 54238 27746 54290
rect 27746 54238 27748 54290
rect 27692 54236 27748 54238
rect 27356 53900 27412 53956
rect 27692 51324 27748 51380
rect 27692 50706 27748 50708
rect 27692 50654 27694 50706
rect 27694 50654 27746 50706
rect 27746 50654 27748 50706
rect 27692 50652 27748 50654
rect 27244 50594 27300 50596
rect 27244 50542 27246 50594
rect 27246 50542 27298 50594
rect 27298 50542 27300 50594
rect 27244 50540 27300 50542
rect 26908 49810 26964 49812
rect 26908 49758 26910 49810
rect 26910 49758 26962 49810
rect 26962 49758 26964 49810
rect 26908 49756 26964 49758
rect 26460 48524 26516 48580
rect 26460 47852 26516 47908
rect 27244 49868 27300 49924
rect 27356 49644 27412 49700
rect 26796 48524 26852 48580
rect 26684 46732 26740 46788
rect 26796 48076 26852 48132
rect 27020 49308 27076 49364
rect 27692 49698 27748 49700
rect 27692 49646 27694 49698
rect 27694 49646 27746 49698
rect 27746 49646 27748 49698
rect 27692 49644 27748 49646
rect 27692 49420 27748 49476
rect 27468 48188 27524 48244
rect 27692 48636 27748 48692
rect 26908 47180 26964 47236
rect 26572 46450 26628 46452
rect 26572 46398 26574 46450
rect 26574 46398 26626 46450
rect 26626 46398 26628 46450
rect 26572 46396 26628 46398
rect 26348 45164 26404 45220
rect 25788 42642 25844 42644
rect 25788 42590 25790 42642
rect 25790 42590 25842 42642
rect 25842 42590 25844 42642
rect 25788 42588 25844 42590
rect 26348 43596 26404 43652
rect 25340 42476 25396 42532
rect 25228 41970 25284 41972
rect 25228 41918 25230 41970
rect 25230 41918 25282 41970
rect 25282 41918 25284 41970
rect 25228 41916 25284 41918
rect 25116 39676 25172 39732
rect 24668 37436 24724 37492
rect 24556 37100 24612 37156
rect 24332 36370 24388 36372
rect 24332 36318 24334 36370
rect 24334 36318 24386 36370
rect 24386 36318 24388 36370
rect 24332 36316 24388 36318
rect 24220 35980 24276 36036
rect 23996 33628 24052 33684
rect 23436 31890 23492 31892
rect 23436 31838 23438 31890
rect 23438 31838 23490 31890
rect 23490 31838 23492 31890
rect 23436 31836 23492 31838
rect 23324 31164 23380 31220
rect 22876 30380 22932 30436
rect 22764 30156 22820 30212
rect 23436 30380 23492 30436
rect 23436 30156 23492 30212
rect 20748 24556 20804 24612
rect 20412 22370 20468 22372
rect 20412 22318 20414 22370
rect 20414 22318 20466 22370
rect 20466 22318 20468 22370
rect 20412 22316 20468 22318
rect 22652 26460 22708 26516
rect 22092 24610 22148 24612
rect 22092 24558 22094 24610
rect 22094 24558 22146 24610
rect 22146 24558 22148 24610
rect 22092 24556 22148 24558
rect 21980 24108 22036 24164
rect 21532 22482 21588 22484
rect 21532 22430 21534 22482
rect 21534 22430 21586 22482
rect 21586 22430 21588 22482
rect 21532 22428 21588 22430
rect 22204 22482 22260 22484
rect 22204 22430 22206 22482
rect 22206 22430 22258 22482
rect 22258 22430 22260 22482
rect 22204 22428 22260 22430
rect 20524 21644 20580 21700
rect 21532 21644 21588 21700
rect 21980 21698 22036 21700
rect 21980 21646 21982 21698
rect 21982 21646 22034 21698
rect 22034 21646 22036 21698
rect 21980 21644 22036 21646
rect 22428 21420 22484 21476
rect 20636 18620 20692 18676
rect 21084 18732 21140 18788
rect 20412 18450 20468 18452
rect 20412 18398 20414 18450
rect 20414 18398 20466 18450
rect 20466 18398 20468 18450
rect 20412 18396 20468 18398
rect 19740 16156 19796 16212
rect 20748 17666 20804 17668
rect 20748 17614 20750 17666
rect 20750 17614 20802 17666
rect 20802 17614 20804 17666
rect 20748 17612 20804 17614
rect 20524 16044 20580 16100
rect 20412 15874 20468 15876
rect 20412 15822 20414 15874
rect 20414 15822 20466 15874
rect 20466 15822 20468 15874
rect 20412 15820 20468 15822
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 19740 15036 19796 15092
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 18956 11900 19012 11956
rect 19292 11788 19348 11844
rect 19628 11900 19684 11956
rect 19740 11788 19796 11844
rect 19740 11564 19796 11620
rect 19852 11452 19908 11508
rect 19964 11282 20020 11284
rect 19964 11230 19966 11282
rect 19966 11230 20018 11282
rect 20018 11230 20020 11282
rect 19964 11228 20020 11230
rect 20300 15372 20356 15428
rect 20860 15148 20916 15204
rect 20188 12012 20244 12068
rect 20412 11676 20468 11732
rect 20188 11564 20244 11620
rect 20188 11394 20244 11396
rect 20188 11342 20190 11394
rect 20190 11342 20242 11394
rect 20242 11342 20244 11394
rect 20188 11340 20244 11342
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 18284 10780 18340 10836
rect 19068 10668 19124 10724
rect 18508 10610 18564 10612
rect 18508 10558 18510 10610
rect 18510 10558 18562 10610
rect 18562 10558 18564 10610
rect 18508 10556 18564 10558
rect 17388 9602 17444 9604
rect 17388 9550 17390 9602
rect 17390 9550 17442 9602
rect 17442 9550 17444 9602
rect 17388 9548 17444 9550
rect 16604 8818 16660 8820
rect 16604 8766 16606 8818
rect 16606 8766 16658 8818
rect 16658 8766 16660 8818
rect 16604 8764 16660 8766
rect 16604 7980 16660 8036
rect 15708 7196 15764 7252
rect 13020 6076 13076 6132
rect 15148 6636 15204 6692
rect 14924 5068 14980 5124
rect 19740 10722 19796 10724
rect 19740 10670 19742 10722
rect 19742 10670 19794 10722
rect 19794 10670 19796 10722
rect 19740 10668 19796 10670
rect 19180 10556 19236 10612
rect 18620 9884 18676 9940
rect 18956 10444 19012 10500
rect 18172 9548 18228 9604
rect 18396 9772 18452 9828
rect 16380 6636 16436 6692
rect 16268 6130 16324 6132
rect 16268 6078 16270 6130
rect 16270 6078 16322 6130
rect 16322 6078 16324 6130
rect 16268 6076 16324 6078
rect 15708 5122 15764 5124
rect 15708 5070 15710 5122
rect 15710 5070 15762 5122
rect 15762 5070 15764 5122
rect 15708 5068 15764 5070
rect 12908 4396 12964 4452
rect 10556 4284 10612 4340
rect 10556 4060 10612 4116
rect 10332 3554 10388 3556
rect 10332 3502 10334 3554
rect 10334 3502 10386 3554
rect 10386 3502 10388 3554
rect 10332 3500 10388 3502
rect 9996 3276 10052 3332
rect 10444 2604 10500 2660
rect 10556 2492 10612 2548
rect 14140 4396 14196 4452
rect 14028 4284 14084 4340
rect 16380 4956 16436 5012
rect 16828 5068 16884 5124
rect 17724 5068 17780 5124
rect 19068 7362 19124 7364
rect 19068 7310 19070 7362
rect 19070 7310 19122 7362
rect 19122 7310 19124 7362
rect 19068 7308 19124 7310
rect 18284 6690 18340 6692
rect 18284 6638 18286 6690
rect 18286 6638 18338 6690
rect 18338 6638 18340 6690
rect 18284 6636 18340 6638
rect 18956 5906 19012 5908
rect 18956 5854 18958 5906
rect 18958 5854 19010 5906
rect 19010 5854 19012 5906
rect 18956 5852 19012 5854
rect 19628 10610 19684 10612
rect 19628 10558 19630 10610
rect 19630 10558 19682 10610
rect 19682 10558 19684 10610
rect 19628 10556 19684 10558
rect 19292 10108 19348 10164
rect 11116 3276 11172 3332
rect 10892 2828 10948 2884
rect 11116 2604 11172 2660
rect 11564 2882 11620 2884
rect 11564 2830 11566 2882
rect 11566 2830 11618 2882
rect 11618 2830 11620 2882
rect 11564 2828 11620 2830
rect 11564 2156 11620 2212
rect 11900 2716 11956 2772
rect 12684 2770 12740 2772
rect 12684 2718 12686 2770
rect 12686 2718 12738 2770
rect 12738 2718 12740 2770
rect 12684 2716 12740 2718
rect 14476 4172 14532 4228
rect 12908 2604 12964 2660
rect 13468 3276 13524 3332
rect 13244 2210 13300 2212
rect 13244 2158 13246 2210
rect 13246 2158 13298 2210
rect 13298 2158 13300 2210
rect 13244 2156 13300 2158
rect 14252 2828 14308 2884
rect 19852 10444 19908 10500
rect 20188 10444 20244 10500
rect 20748 11564 20804 11620
rect 20524 11116 20580 11172
rect 20636 10834 20692 10836
rect 20636 10782 20638 10834
rect 20638 10782 20690 10834
rect 20690 10782 20692 10834
rect 20636 10780 20692 10782
rect 20524 10556 20580 10612
rect 19964 9548 20020 9604
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 19740 8764 19796 8820
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 19516 4844 19572 4900
rect 21196 19964 21252 20020
rect 23100 29932 23156 29988
rect 22876 26348 22932 26404
rect 22988 26178 23044 26180
rect 22988 26126 22990 26178
rect 22990 26126 23042 26178
rect 23042 26126 23044 26178
rect 22988 26124 23044 26126
rect 23100 25564 23156 25620
rect 23100 25340 23156 25396
rect 23436 29650 23492 29652
rect 23436 29598 23438 29650
rect 23438 29598 23490 29650
rect 23490 29598 23492 29650
rect 23436 29596 23492 29598
rect 23548 26908 23604 26964
rect 24220 31778 24276 31780
rect 24220 31726 24222 31778
rect 24222 31726 24274 31778
rect 24274 31726 24276 31778
rect 24220 31724 24276 31726
rect 24220 31218 24276 31220
rect 24220 31166 24222 31218
rect 24222 31166 24274 31218
rect 24274 31166 24276 31218
rect 24220 31164 24276 31166
rect 24108 29596 24164 29652
rect 24668 31778 24724 31780
rect 24668 31726 24670 31778
rect 24670 31726 24722 31778
rect 24722 31726 24724 31778
rect 24668 31724 24724 31726
rect 23772 28812 23828 28868
rect 24444 29260 24500 29316
rect 23996 28140 24052 28196
rect 23436 26514 23492 26516
rect 23436 26462 23438 26514
rect 23438 26462 23490 26514
rect 23490 26462 23492 26514
rect 23436 26460 23492 26462
rect 23772 26402 23828 26404
rect 23772 26350 23774 26402
rect 23774 26350 23826 26402
rect 23826 26350 23828 26402
rect 23772 26348 23828 26350
rect 23436 25228 23492 25284
rect 22764 19404 22820 19460
rect 23324 23772 23380 23828
rect 23436 23436 23492 23492
rect 24780 29260 24836 29316
rect 24668 28140 24724 28196
rect 24332 26908 24388 26964
rect 24444 26124 24500 26180
rect 24108 24892 24164 24948
rect 24220 25340 24276 25396
rect 24444 24108 24500 24164
rect 24108 23436 24164 23492
rect 23324 22428 23380 22484
rect 22652 17666 22708 17668
rect 22652 17614 22654 17666
rect 22654 17614 22706 17666
rect 22706 17614 22708 17666
rect 22652 17612 22708 17614
rect 22652 16940 22708 16996
rect 21644 16268 21700 16324
rect 21420 16098 21476 16100
rect 21420 16046 21422 16098
rect 21422 16046 21474 16098
rect 21474 16046 21476 16098
rect 21420 16044 21476 16046
rect 22092 16322 22148 16324
rect 22092 16270 22094 16322
rect 22094 16270 22146 16322
rect 22146 16270 22148 16322
rect 22092 16268 22148 16270
rect 21868 16210 21924 16212
rect 21868 16158 21870 16210
rect 21870 16158 21922 16210
rect 21922 16158 21924 16210
rect 21868 16156 21924 16158
rect 21868 15202 21924 15204
rect 21868 15150 21870 15202
rect 21870 15150 21922 15202
rect 21922 15150 21924 15202
rect 21868 15148 21924 15150
rect 21868 14530 21924 14532
rect 21868 14478 21870 14530
rect 21870 14478 21922 14530
rect 21922 14478 21924 14530
rect 21868 14476 21924 14478
rect 23324 19964 23380 20020
rect 24444 23884 24500 23940
rect 23884 20018 23940 20020
rect 23884 19966 23886 20018
rect 23886 19966 23938 20018
rect 23938 19966 23940 20018
rect 23884 19964 23940 19966
rect 24780 26290 24836 26292
rect 24780 26238 24782 26290
rect 24782 26238 24834 26290
rect 24834 26238 24836 26290
rect 24780 26236 24836 26238
rect 25676 42364 25732 42420
rect 25452 42194 25508 42196
rect 25452 42142 25454 42194
rect 25454 42142 25506 42194
rect 25506 42142 25508 42194
rect 25452 42140 25508 42142
rect 26236 42252 26292 42308
rect 26684 45836 26740 45892
rect 26572 45164 26628 45220
rect 26572 44604 26628 44660
rect 26460 43372 26516 43428
rect 26796 45778 26852 45780
rect 26796 45726 26798 45778
rect 26798 45726 26850 45778
rect 26850 45726 26852 45778
rect 26796 45724 26852 45726
rect 27244 46956 27300 47012
rect 27916 55298 27972 55300
rect 27916 55246 27918 55298
rect 27918 55246 27970 55298
rect 27970 55246 27972 55298
rect 27916 55244 27972 55246
rect 28476 55298 28532 55300
rect 28476 55246 28478 55298
rect 28478 55246 28530 55298
rect 28530 55246 28532 55298
rect 28476 55244 28532 55246
rect 28364 54684 28420 54740
rect 27916 54626 27972 54628
rect 27916 54574 27918 54626
rect 27918 54574 27970 54626
rect 27970 54574 27972 54626
rect 27916 54572 27972 54574
rect 28364 54236 28420 54292
rect 28028 52780 28084 52836
rect 28028 50540 28084 50596
rect 28252 48802 28308 48804
rect 28252 48750 28254 48802
rect 28254 48750 28306 48802
rect 28306 48750 28308 48802
rect 28252 48748 28308 48750
rect 28028 48466 28084 48468
rect 28028 48414 28030 48466
rect 28030 48414 28082 48466
rect 28082 48414 28084 48466
rect 28028 48412 28084 48414
rect 28476 53788 28532 53844
rect 28588 52834 28644 52836
rect 28588 52782 28590 52834
rect 28590 52782 28642 52834
rect 28642 52782 28644 52834
rect 28588 52780 28644 52782
rect 28476 49420 28532 49476
rect 28476 47404 28532 47460
rect 27916 46844 27972 46900
rect 28140 46562 28196 46564
rect 28140 46510 28142 46562
rect 28142 46510 28194 46562
rect 28194 46510 28196 46562
rect 28140 46508 28196 46510
rect 26908 45106 26964 45108
rect 26908 45054 26910 45106
rect 26910 45054 26962 45106
rect 26962 45054 26964 45106
rect 26908 45052 26964 45054
rect 26796 43596 26852 43652
rect 27020 43596 27076 43652
rect 26572 43484 26628 43540
rect 26348 42028 26404 42084
rect 27580 45164 27636 45220
rect 28588 48412 28644 48468
rect 28364 46396 28420 46452
rect 28588 46674 28644 46676
rect 28588 46622 28590 46674
rect 28590 46622 28642 46674
rect 28642 46622 28644 46674
rect 28588 46620 28644 46622
rect 28476 45948 28532 46004
rect 28364 45836 28420 45892
rect 28252 45388 28308 45444
rect 28588 45276 28644 45332
rect 27356 45052 27412 45108
rect 28364 45164 28420 45220
rect 27356 44380 27412 44436
rect 27580 44604 27636 44660
rect 27916 44098 27972 44100
rect 27916 44046 27918 44098
rect 27918 44046 27970 44098
rect 27970 44046 27972 44098
rect 27916 44044 27972 44046
rect 27356 43596 27412 43652
rect 27916 43596 27972 43652
rect 27132 43372 27188 43428
rect 27020 43260 27076 43316
rect 26684 43036 26740 43092
rect 26684 42364 26740 42420
rect 26236 41970 26292 41972
rect 26236 41918 26238 41970
rect 26238 41918 26290 41970
rect 26290 41918 26292 41970
rect 26236 41916 26292 41918
rect 26236 41692 26292 41748
rect 26236 41468 26292 41524
rect 25676 41186 25732 41188
rect 25676 41134 25678 41186
rect 25678 41134 25730 41186
rect 25730 41134 25732 41186
rect 25676 41132 25732 41134
rect 25900 40626 25956 40628
rect 25900 40574 25902 40626
rect 25902 40574 25954 40626
rect 25954 40574 25956 40626
rect 25900 40572 25956 40574
rect 26572 41074 26628 41076
rect 26572 41022 26574 41074
rect 26574 41022 26626 41074
rect 26626 41022 26628 41074
rect 26572 41020 26628 41022
rect 27468 43148 27524 43204
rect 27244 41916 27300 41972
rect 25676 39564 25732 39620
rect 25340 39452 25396 39508
rect 25228 37772 25284 37828
rect 26460 39618 26516 39620
rect 26460 39566 26462 39618
rect 26462 39566 26514 39618
rect 26514 39566 26516 39618
rect 26460 39564 26516 39566
rect 26012 39452 26068 39508
rect 25900 39340 25956 39396
rect 25340 37154 25396 37156
rect 25340 37102 25342 37154
rect 25342 37102 25394 37154
rect 25394 37102 25396 37154
rect 25340 37100 25396 37102
rect 25004 36204 25060 36260
rect 25228 34860 25284 34916
rect 25228 32956 25284 33012
rect 25564 34914 25620 34916
rect 25564 34862 25566 34914
rect 25566 34862 25618 34914
rect 25618 34862 25620 34914
rect 25564 34860 25620 34862
rect 25788 39004 25844 39060
rect 26460 39116 26516 39172
rect 26012 37772 26068 37828
rect 25788 37490 25844 37492
rect 25788 37438 25790 37490
rect 25790 37438 25842 37490
rect 25842 37438 25844 37490
rect 25788 37436 25844 37438
rect 25788 37100 25844 37156
rect 25676 31778 25732 31780
rect 25676 31726 25678 31778
rect 25678 31726 25730 31778
rect 25730 31726 25732 31778
rect 25676 31724 25732 31726
rect 25452 28476 25508 28532
rect 26012 36370 26068 36372
rect 26012 36318 26014 36370
rect 26014 36318 26066 36370
rect 26066 36318 26068 36370
rect 26012 36316 26068 36318
rect 26460 33068 26516 33124
rect 25900 29650 25956 29652
rect 25900 29598 25902 29650
rect 25902 29598 25954 29650
rect 25954 29598 25956 29650
rect 25900 29596 25956 29598
rect 25564 27970 25620 27972
rect 25564 27918 25566 27970
rect 25566 27918 25618 27970
rect 25618 27918 25620 27970
rect 25564 27916 25620 27918
rect 25116 25506 25172 25508
rect 25116 25454 25118 25506
rect 25118 25454 25170 25506
rect 25170 25454 25172 25506
rect 25116 25452 25172 25454
rect 25004 24108 25060 24164
rect 24668 23436 24724 23492
rect 23100 16994 23156 16996
rect 23100 16942 23102 16994
rect 23102 16942 23154 16994
rect 23154 16942 23156 16994
rect 23100 16940 23156 16942
rect 22876 16268 22932 16324
rect 22764 14476 22820 14532
rect 21196 11676 21252 11732
rect 21756 11564 21812 11620
rect 21420 11394 21476 11396
rect 21420 11342 21422 11394
rect 21422 11342 21474 11394
rect 21474 11342 21476 11394
rect 21420 11340 21476 11342
rect 21196 11116 21252 11172
rect 23884 15538 23940 15540
rect 23884 15486 23886 15538
rect 23886 15486 23938 15538
rect 23938 15486 23940 15538
rect 23884 15484 23940 15486
rect 23996 17724 24052 17780
rect 25228 23826 25284 23828
rect 25228 23774 25230 23826
rect 25230 23774 25282 23826
rect 25282 23774 25284 23826
rect 25228 23772 25284 23774
rect 25452 26850 25508 26852
rect 25452 26798 25454 26850
rect 25454 26798 25506 26850
rect 25506 26798 25508 26850
rect 25452 26796 25508 26798
rect 25676 26460 25732 26516
rect 25900 26962 25956 26964
rect 25900 26910 25902 26962
rect 25902 26910 25954 26962
rect 25954 26910 25956 26962
rect 25900 26908 25956 26910
rect 26908 40178 26964 40180
rect 26908 40126 26910 40178
rect 26910 40126 26962 40178
rect 26962 40126 26964 40178
rect 26908 40124 26964 40126
rect 28140 42754 28196 42756
rect 28140 42702 28142 42754
rect 28142 42702 28194 42754
rect 28194 42702 28196 42754
rect 28140 42700 28196 42702
rect 28476 42140 28532 42196
rect 27692 41916 27748 41972
rect 27468 41298 27524 41300
rect 27468 41246 27470 41298
rect 27470 41246 27522 41298
rect 27522 41246 27524 41298
rect 27468 41244 27524 41246
rect 27468 39506 27524 39508
rect 27468 39454 27470 39506
rect 27470 39454 27522 39506
rect 27522 39454 27524 39506
rect 27468 39452 27524 39454
rect 27132 39228 27188 39284
rect 27244 38834 27300 38836
rect 27244 38782 27246 38834
rect 27246 38782 27298 38834
rect 27298 38782 27300 38834
rect 27244 38780 27300 38782
rect 28252 41858 28308 41860
rect 28252 41806 28254 41858
rect 28254 41806 28306 41858
rect 28306 41806 28308 41858
rect 28252 41804 28308 41806
rect 28364 41356 28420 41412
rect 28140 41020 28196 41076
rect 27916 40962 27972 40964
rect 27916 40910 27918 40962
rect 27918 40910 27970 40962
rect 27970 40910 27972 40962
rect 27916 40908 27972 40910
rect 27804 40572 27860 40628
rect 28588 40236 28644 40292
rect 26908 37826 26964 37828
rect 26908 37774 26910 37826
rect 26910 37774 26962 37826
rect 26962 37774 26964 37826
rect 26908 37772 26964 37774
rect 27132 37324 27188 37380
rect 26684 35810 26740 35812
rect 26684 35758 26686 35810
rect 26686 35758 26738 35810
rect 26738 35758 26740 35810
rect 26684 35756 26740 35758
rect 26684 34860 26740 34916
rect 27020 34636 27076 34692
rect 27356 35420 27412 35476
rect 27132 33516 27188 33572
rect 27356 33180 27412 33236
rect 27132 33122 27188 33124
rect 27132 33070 27134 33122
rect 27134 33070 27186 33122
rect 27186 33070 27188 33122
rect 27132 33068 27188 33070
rect 28140 37378 28196 37380
rect 28140 37326 28142 37378
rect 28142 37326 28194 37378
rect 28194 37326 28196 37378
rect 28140 37324 28196 37326
rect 28140 35868 28196 35924
rect 28364 36204 28420 36260
rect 28252 34636 28308 34692
rect 28140 34076 28196 34132
rect 27692 33570 27748 33572
rect 27692 33518 27694 33570
rect 27694 33518 27746 33570
rect 27746 33518 27748 33570
rect 27692 33516 27748 33518
rect 28028 33346 28084 33348
rect 28028 33294 28030 33346
rect 28030 33294 28082 33346
rect 28082 33294 28084 33346
rect 28028 33292 28084 33294
rect 26908 31948 26964 32004
rect 26684 31724 26740 31780
rect 26908 31612 26964 31668
rect 26572 29484 26628 29540
rect 26348 29372 26404 29428
rect 26684 29426 26740 29428
rect 26684 29374 26686 29426
rect 26686 29374 26738 29426
rect 26738 29374 26740 29426
rect 26684 29372 26740 29374
rect 26796 29148 26852 29204
rect 26124 26684 26180 26740
rect 25452 26290 25508 26292
rect 25452 26238 25454 26290
rect 25454 26238 25506 26290
rect 25506 26238 25508 26290
rect 25452 26236 25508 26238
rect 25900 26012 25956 26068
rect 25676 25452 25732 25508
rect 26348 26348 26404 26404
rect 27244 29650 27300 29652
rect 27244 29598 27246 29650
rect 27246 29598 27298 29650
rect 27298 29598 27300 29650
rect 27244 29596 27300 29598
rect 27468 28866 27524 28868
rect 27468 28814 27470 28866
rect 27470 28814 27522 28866
rect 27522 28814 27524 28866
rect 27468 28812 27524 28814
rect 26796 28476 26852 28532
rect 27468 28140 27524 28196
rect 28476 35644 28532 35700
rect 29148 60844 29204 60900
rect 29148 59948 29204 60004
rect 30716 66162 30772 66164
rect 30716 66110 30718 66162
rect 30718 66110 30770 66162
rect 30770 66110 30772 66162
rect 30716 66108 30772 66110
rect 30940 69692 30996 69748
rect 30940 66780 30996 66836
rect 30940 66108 30996 66164
rect 30604 65490 30660 65492
rect 30604 65438 30606 65490
rect 30606 65438 30658 65490
rect 30658 65438 30660 65490
rect 30604 65436 30660 65438
rect 30940 65602 30996 65604
rect 30940 65550 30942 65602
rect 30942 65550 30994 65602
rect 30994 65550 30996 65602
rect 30940 65548 30996 65550
rect 30828 64428 30884 64484
rect 31164 70194 31220 70196
rect 31164 70142 31166 70194
rect 31166 70142 31218 70194
rect 31218 70142 31220 70194
rect 31164 70140 31220 70142
rect 31164 68908 31220 68964
rect 31836 75516 31892 75572
rect 32396 75570 32452 75572
rect 32396 75518 32398 75570
rect 32398 75518 32450 75570
rect 32450 75518 32452 75570
rect 32396 75516 32452 75518
rect 31724 75122 31780 75124
rect 31724 75070 31726 75122
rect 31726 75070 31778 75122
rect 31778 75070 31780 75122
rect 31724 75068 31780 75070
rect 31836 75180 31892 75236
rect 33292 75292 33348 75348
rect 33404 76188 33460 76244
rect 31724 70700 31780 70756
rect 32508 75122 32564 75124
rect 32508 75070 32510 75122
rect 32510 75070 32562 75122
rect 32562 75070 32564 75122
rect 32508 75068 32564 75070
rect 31948 73836 32004 73892
rect 31836 70364 31892 70420
rect 32172 72044 32228 72100
rect 31836 70194 31892 70196
rect 31836 70142 31838 70194
rect 31838 70142 31890 70194
rect 31890 70142 31892 70194
rect 31836 70140 31892 70142
rect 32396 71986 32452 71988
rect 32396 71934 32398 71986
rect 32398 71934 32450 71986
rect 32450 71934 32452 71986
rect 32396 71932 32452 71934
rect 33516 75570 33572 75572
rect 33516 75518 33518 75570
rect 33518 75518 33570 75570
rect 33570 75518 33572 75570
rect 33516 75516 33572 75518
rect 34748 77420 34804 77476
rect 35868 78594 35924 78596
rect 35868 78542 35870 78594
rect 35870 78542 35922 78594
rect 35922 78542 35924 78594
rect 35868 78540 35924 78542
rect 35756 78092 35812 78148
rect 35868 78034 35924 78036
rect 35868 77982 35870 78034
rect 35870 77982 35922 78034
rect 35922 77982 35924 78034
rect 35868 77980 35924 77982
rect 35196 77642 35252 77644
rect 35196 77590 35198 77642
rect 35198 77590 35250 77642
rect 35250 77590 35252 77642
rect 35196 77588 35252 77590
rect 35300 77642 35356 77644
rect 35300 77590 35302 77642
rect 35302 77590 35354 77642
rect 35354 77590 35356 77642
rect 35300 77588 35356 77590
rect 35404 77642 35460 77644
rect 35404 77590 35406 77642
rect 35406 77590 35458 77642
rect 35458 77590 35460 77642
rect 35404 77588 35460 77590
rect 35756 77532 35812 77588
rect 34412 76524 34468 76580
rect 35644 77362 35700 77364
rect 35644 77310 35646 77362
rect 35646 77310 35698 77362
rect 35698 77310 35700 77362
rect 35644 77308 35700 77310
rect 35420 76972 35476 77028
rect 35420 76748 35476 76804
rect 33964 76466 34020 76468
rect 33964 76414 33966 76466
rect 33966 76414 34018 76466
rect 34018 76414 34020 76466
rect 33964 76412 34020 76414
rect 34188 76242 34244 76244
rect 34188 76190 34190 76242
rect 34190 76190 34242 76242
rect 34242 76190 34244 76242
rect 34188 76188 34244 76190
rect 34524 76242 34580 76244
rect 34524 76190 34526 76242
rect 34526 76190 34578 76242
rect 34578 76190 34580 76242
rect 34524 76188 34580 76190
rect 34076 75906 34132 75908
rect 34076 75854 34078 75906
rect 34078 75854 34130 75906
rect 34130 75854 34132 75906
rect 34076 75852 34132 75854
rect 34412 75682 34468 75684
rect 34412 75630 34414 75682
rect 34414 75630 34466 75682
rect 34466 75630 34468 75682
rect 34412 75628 34468 75630
rect 33740 75458 33796 75460
rect 33740 75406 33742 75458
rect 33742 75406 33794 75458
rect 33794 75406 33796 75458
rect 33740 75404 33796 75406
rect 33964 75292 34020 75348
rect 32508 71148 32564 71204
rect 32732 74732 32788 74788
rect 32732 74060 32788 74116
rect 34076 75068 34132 75124
rect 35308 76466 35364 76468
rect 35308 76414 35310 76466
rect 35310 76414 35362 76466
rect 35362 76414 35364 76466
rect 35308 76412 35364 76414
rect 37996 78540 38052 78596
rect 37324 78204 37380 78260
rect 37100 78146 37156 78148
rect 37100 78094 37102 78146
rect 37102 78094 37154 78146
rect 37154 78094 37156 78146
rect 37100 78092 37156 78094
rect 36092 77868 36148 77924
rect 36316 77922 36372 77924
rect 36316 77870 36318 77922
rect 36318 77870 36370 77922
rect 36370 77870 36372 77922
rect 36316 77868 36372 77870
rect 36540 77810 36596 77812
rect 36540 77758 36542 77810
rect 36542 77758 36594 77810
rect 36594 77758 36596 77810
rect 36540 77756 36596 77758
rect 36204 77420 36260 77476
rect 36652 77420 36708 77476
rect 36428 77250 36484 77252
rect 36428 77198 36430 77250
rect 36430 77198 36482 77250
rect 36482 77198 36484 77250
rect 36428 77196 36484 77198
rect 35532 76188 35588 76244
rect 35196 76074 35252 76076
rect 35196 76022 35198 76074
rect 35198 76022 35250 76074
rect 35250 76022 35252 76074
rect 35196 76020 35252 76022
rect 35300 76074 35356 76076
rect 35300 76022 35302 76074
rect 35302 76022 35354 76074
rect 35354 76022 35356 76074
rect 35300 76020 35356 76022
rect 35404 76074 35460 76076
rect 35404 76022 35406 76074
rect 35406 76022 35458 76074
rect 35458 76022 35460 76074
rect 35404 76020 35460 76022
rect 34636 75404 34692 75460
rect 34636 74956 34692 75012
rect 34972 75570 35028 75572
rect 34972 75518 34974 75570
rect 34974 75518 35026 75570
rect 35026 75518 35028 75570
rect 34972 75516 35028 75518
rect 34972 74956 35028 75012
rect 35308 75404 35364 75460
rect 35196 75068 35252 75124
rect 36092 76524 36148 76580
rect 36092 75682 36148 75684
rect 36092 75630 36094 75682
rect 36094 75630 36146 75682
rect 36146 75630 36148 75682
rect 36092 75628 36148 75630
rect 36428 76748 36484 76804
rect 36316 76524 36372 76580
rect 36092 75404 36148 75460
rect 35980 75292 36036 75348
rect 35980 75068 36036 75124
rect 35756 74620 35812 74676
rect 35196 74506 35252 74508
rect 35196 74454 35198 74506
rect 35198 74454 35250 74506
rect 35250 74454 35252 74506
rect 35196 74452 35252 74454
rect 35300 74506 35356 74508
rect 35300 74454 35302 74506
rect 35302 74454 35354 74506
rect 35354 74454 35356 74506
rect 35300 74452 35356 74454
rect 35404 74506 35460 74508
rect 35404 74454 35406 74506
rect 35406 74454 35458 74506
rect 35458 74454 35460 74506
rect 35404 74452 35460 74454
rect 35308 74284 35364 74340
rect 35756 74338 35812 74340
rect 35756 74286 35758 74338
rect 35758 74286 35810 74338
rect 35810 74286 35812 74338
rect 35756 74284 35812 74286
rect 35420 74060 35476 74116
rect 36428 76412 36484 76468
rect 36316 75122 36372 75124
rect 36316 75070 36318 75122
rect 36318 75070 36370 75122
rect 36370 75070 36372 75122
rect 36316 75068 36372 75070
rect 37212 78034 37268 78036
rect 37212 77982 37214 78034
rect 37214 77982 37266 78034
rect 37266 77982 37268 78034
rect 37212 77980 37268 77982
rect 37212 77474 37268 77476
rect 37212 77422 37214 77474
rect 37214 77422 37266 77474
rect 37266 77422 37268 77474
rect 37212 77420 37268 77422
rect 36876 77196 36932 77252
rect 37884 77474 37940 77476
rect 37884 77422 37886 77474
rect 37886 77422 37938 77474
rect 37938 77422 37940 77474
rect 37884 77420 37940 77422
rect 36988 77084 37044 77140
rect 37100 77026 37156 77028
rect 37100 76974 37102 77026
rect 37102 76974 37154 77026
rect 37154 76974 37156 77026
rect 37100 76972 37156 76974
rect 37212 76748 37268 76804
rect 37436 77250 37492 77252
rect 37436 77198 37438 77250
rect 37438 77198 37490 77250
rect 37490 77198 37492 77250
rect 37436 77196 37492 77198
rect 38108 77196 38164 77252
rect 37660 76860 37716 76916
rect 37884 76578 37940 76580
rect 37884 76526 37886 76578
rect 37886 76526 37938 76578
rect 37938 76526 37940 76578
rect 37884 76524 37940 76526
rect 37100 76466 37156 76468
rect 37100 76414 37102 76466
rect 37102 76414 37154 76466
rect 37154 76414 37156 76466
rect 37100 76412 37156 76414
rect 37436 76300 37492 76356
rect 37996 75852 38052 75908
rect 37100 75794 37156 75796
rect 37100 75742 37102 75794
rect 37102 75742 37154 75794
rect 37154 75742 37156 75794
rect 37100 75740 37156 75742
rect 37212 75628 37268 75684
rect 36988 75570 37044 75572
rect 36988 75518 36990 75570
rect 36990 75518 37042 75570
rect 37042 75518 37044 75570
rect 36988 75516 37044 75518
rect 37436 75068 37492 75124
rect 36428 74620 36484 74676
rect 38220 74898 38276 74900
rect 38220 74846 38222 74898
rect 38222 74846 38274 74898
rect 38274 74846 38276 74898
rect 38220 74844 38276 74846
rect 37660 74786 37716 74788
rect 37660 74734 37662 74786
rect 37662 74734 37714 74786
rect 37714 74734 37716 74786
rect 37660 74732 37716 74734
rect 36876 74620 36932 74676
rect 36092 74060 36148 74116
rect 33628 72156 33684 72212
rect 33740 72268 33796 72324
rect 32732 70978 32788 70980
rect 32732 70926 32734 70978
rect 32734 70926 32786 70978
rect 32786 70926 32788 70978
rect 32732 70924 32788 70926
rect 32284 70812 32340 70868
rect 33852 72044 33908 72100
rect 34076 73500 34132 73556
rect 35756 73890 35812 73892
rect 35756 73838 35758 73890
rect 35758 73838 35810 73890
rect 35810 73838 35812 73890
rect 35756 73836 35812 73838
rect 35196 72938 35252 72940
rect 35196 72886 35198 72938
rect 35198 72886 35250 72938
rect 35250 72886 35252 72938
rect 35196 72884 35252 72886
rect 35300 72938 35356 72940
rect 35300 72886 35302 72938
rect 35302 72886 35354 72938
rect 35354 72886 35356 72938
rect 35300 72884 35356 72886
rect 35404 72938 35460 72940
rect 35404 72886 35406 72938
rect 35406 72886 35458 72938
rect 35458 72886 35460 72938
rect 35404 72884 35460 72886
rect 34076 72156 34132 72212
rect 33740 71932 33796 71988
rect 33292 71484 33348 71540
rect 33404 70812 33460 70868
rect 33628 71148 33684 71204
rect 34412 71874 34468 71876
rect 34412 71822 34414 71874
rect 34414 71822 34466 71874
rect 34466 71822 34468 71874
rect 34412 71820 34468 71822
rect 33068 69692 33124 69748
rect 33404 69916 33460 69972
rect 32284 69356 32340 69412
rect 31164 67116 31220 67172
rect 31164 65996 31220 66052
rect 31276 66108 31332 66164
rect 31388 65324 31444 65380
rect 30828 63644 30884 63700
rect 30492 62578 30548 62580
rect 30492 62526 30494 62578
rect 30494 62526 30546 62578
rect 30546 62526 30548 62578
rect 30492 62524 30548 62526
rect 30156 61852 30212 61908
rect 29484 60844 29540 60900
rect 29932 60002 29988 60004
rect 29932 59950 29934 60002
rect 29934 59950 29986 60002
rect 29986 59950 29988 60002
rect 29932 59948 29988 59950
rect 30268 59948 30324 60004
rect 29260 59724 29316 59780
rect 29148 56866 29204 56868
rect 29148 56814 29150 56866
rect 29150 56814 29202 56866
rect 29202 56814 29204 56866
rect 29148 56812 29204 56814
rect 28812 54514 28868 54516
rect 28812 54462 28814 54514
rect 28814 54462 28866 54514
rect 28866 54462 28868 54514
rect 28812 54460 28868 54462
rect 29148 54460 29204 54516
rect 28924 53676 28980 53732
rect 28812 48748 28868 48804
rect 28812 46508 28868 46564
rect 29148 52780 29204 52836
rect 29596 59724 29652 59780
rect 30156 59724 30212 59780
rect 29820 59442 29876 59444
rect 29820 59390 29822 59442
rect 29822 59390 29874 59442
rect 29874 59390 29876 59442
rect 29820 59388 29876 59390
rect 29484 59164 29540 59220
rect 29484 58210 29540 58212
rect 29484 58158 29486 58210
rect 29486 58158 29538 58210
rect 29538 58158 29540 58210
rect 29484 58156 29540 58158
rect 29708 57260 29764 57316
rect 29820 58268 29876 58324
rect 29372 54572 29428 54628
rect 29372 53788 29428 53844
rect 30268 58546 30324 58548
rect 30268 58494 30270 58546
rect 30270 58494 30322 58546
rect 30322 58494 30324 58546
rect 30268 58492 30324 58494
rect 30716 61852 30772 61908
rect 30492 61570 30548 61572
rect 30492 61518 30494 61570
rect 30494 61518 30546 61570
rect 30546 61518 30548 61570
rect 30492 61516 30548 61518
rect 30492 59948 30548 60004
rect 30492 59218 30548 59220
rect 30492 59166 30494 59218
rect 30494 59166 30546 59218
rect 30546 59166 30548 59218
rect 30492 59164 30548 59166
rect 30604 58492 30660 58548
rect 30380 57260 30436 57316
rect 30604 56924 30660 56980
rect 31052 61516 31108 61572
rect 30828 60786 30884 60788
rect 30828 60734 30830 60786
rect 30830 60734 30882 60786
rect 30882 60734 30884 60786
rect 30828 60732 30884 60734
rect 30940 57260 30996 57316
rect 30940 56306 30996 56308
rect 30940 56254 30942 56306
rect 30942 56254 30994 56306
rect 30994 56254 30996 56306
rect 30940 56252 30996 56254
rect 30044 54738 30100 54740
rect 30044 54686 30046 54738
rect 30046 54686 30098 54738
rect 30098 54686 30100 54738
rect 30044 54684 30100 54686
rect 30156 54402 30212 54404
rect 30156 54350 30158 54402
rect 30158 54350 30210 54402
rect 30210 54350 30212 54402
rect 30156 54348 30212 54350
rect 29484 53676 29540 53732
rect 29036 46060 29092 46116
rect 29260 48802 29316 48804
rect 29260 48750 29262 48802
rect 29262 48750 29314 48802
rect 29314 48750 29316 48802
rect 29260 48748 29316 48750
rect 30492 53676 30548 53732
rect 29372 48412 29428 48468
rect 30380 51378 30436 51380
rect 30380 51326 30382 51378
rect 30382 51326 30434 51378
rect 30434 51326 30436 51378
rect 30380 51324 30436 51326
rect 29708 49420 29764 49476
rect 29036 45724 29092 45780
rect 29036 44604 29092 44660
rect 29260 44210 29316 44212
rect 29260 44158 29262 44210
rect 29262 44158 29314 44210
rect 29314 44158 29316 44210
rect 29260 44156 29316 44158
rect 28924 42252 28980 42308
rect 28700 34524 28756 34580
rect 28588 33516 28644 33572
rect 28476 33404 28532 33460
rect 28364 33180 28420 33236
rect 29260 41692 29316 41748
rect 29148 40402 29204 40404
rect 29148 40350 29150 40402
rect 29150 40350 29202 40402
rect 29202 40350 29204 40402
rect 29148 40348 29204 40350
rect 29708 44434 29764 44436
rect 29708 44382 29710 44434
rect 29710 44382 29762 44434
rect 29762 44382 29764 44434
rect 29708 44380 29764 44382
rect 29484 43484 29540 43540
rect 29596 43426 29652 43428
rect 29596 43374 29598 43426
rect 29598 43374 29650 43426
rect 29650 43374 29652 43426
rect 29596 43372 29652 43374
rect 29484 43036 29540 43092
rect 29708 42252 29764 42308
rect 30380 50876 30436 50932
rect 30268 49420 30324 49476
rect 32060 68684 32116 68740
rect 31948 68514 32004 68516
rect 31948 68462 31950 68514
rect 31950 68462 32002 68514
rect 32002 68462 32004 68514
rect 31948 68460 32004 68462
rect 31836 68402 31892 68404
rect 31836 68350 31838 68402
rect 31838 68350 31890 68402
rect 31890 68350 31892 68402
rect 31836 68348 31892 68350
rect 32396 68460 32452 68516
rect 31724 67954 31780 67956
rect 31724 67902 31726 67954
rect 31726 67902 31778 67954
rect 31778 67902 31780 67954
rect 31724 67900 31780 67902
rect 32956 68796 33012 68852
rect 33068 68738 33124 68740
rect 33068 68686 33070 68738
rect 33070 68686 33122 68738
rect 33122 68686 33124 68738
rect 33068 68684 33124 68686
rect 33404 68124 33460 68180
rect 33068 68066 33124 68068
rect 33068 68014 33070 68066
rect 33070 68014 33122 68066
rect 33122 68014 33124 68066
rect 33068 68012 33124 68014
rect 32508 67228 32564 67284
rect 32956 67788 33012 67844
rect 31836 66162 31892 66164
rect 31836 66110 31838 66162
rect 31838 66110 31890 66162
rect 31890 66110 31892 66162
rect 31836 66108 31892 66110
rect 31612 65378 31668 65380
rect 31612 65326 31614 65378
rect 31614 65326 31666 65378
rect 31666 65326 31668 65378
rect 31612 65324 31668 65326
rect 31388 64540 31444 64596
rect 31500 62076 31556 62132
rect 31276 59836 31332 59892
rect 31276 58268 31332 58324
rect 31164 55356 31220 55412
rect 31276 54684 31332 54740
rect 34076 70418 34132 70420
rect 34076 70366 34078 70418
rect 34078 70366 34130 70418
rect 34130 70366 34132 70418
rect 34076 70364 34132 70366
rect 33740 68796 33796 68852
rect 33628 68460 33684 68516
rect 33740 67900 33796 67956
rect 32396 65212 32452 65268
rect 31948 64204 32004 64260
rect 32284 64482 32340 64484
rect 32284 64430 32286 64482
rect 32286 64430 32338 64482
rect 32338 64430 32340 64482
rect 32284 64428 32340 64430
rect 32284 64034 32340 64036
rect 32284 63982 32286 64034
rect 32286 63982 32338 64034
rect 32338 63982 32340 64034
rect 32284 63980 32340 63982
rect 32172 63308 32228 63364
rect 31724 61628 31780 61684
rect 32060 61516 32116 61572
rect 31948 61180 32004 61236
rect 32284 61740 32340 61796
rect 32284 61570 32340 61572
rect 32284 61518 32286 61570
rect 32286 61518 32338 61570
rect 32338 61518 32340 61570
rect 32284 61516 32340 61518
rect 32284 61010 32340 61012
rect 32284 60958 32286 61010
rect 32286 60958 32338 61010
rect 32338 60958 32340 61010
rect 32284 60956 32340 60958
rect 33404 67228 33460 67284
rect 33628 66332 33684 66388
rect 33292 66274 33348 66276
rect 33292 66222 33294 66274
rect 33294 66222 33346 66274
rect 33346 66222 33348 66274
rect 33292 66220 33348 66222
rect 33516 66162 33572 66164
rect 33516 66110 33518 66162
rect 33518 66110 33570 66162
rect 33570 66110 33572 66162
rect 33516 66108 33572 66110
rect 33292 65714 33348 65716
rect 33292 65662 33294 65714
rect 33294 65662 33346 65714
rect 33346 65662 33348 65714
rect 33292 65660 33348 65662
rect 33628 65548 33684 65604
rect 34636 71148 34692 71204
rect 34748 71820 34804 71876
rect 34748 70588 34804 70644
rect 34412 70194 34468 70196
rect 34412 70142 34414 70194
rect 34414 70142 34466 70194
rect 34466 70142 34468 70194
rect 34412 70140 34468 70142
rect 34300 68684 34356 68740
rect 33852 68348 33908 68404
rect 34188 68124 34244 68180
rect 34412 68066 34468 68068
rect 34412 68014 34414 68066
rect 34414 68014 34466 68066
rect 34466 68014 34468 68066
rect 34412 68012 34468 68014
rect 35644 72322 35700 72324
rect 35644 72270 35646 72322
rect 35646 72270 35698 72322
rect 35698 72270 35700 72322
rect 35644 72268 35700 72270
rect 35532 71538 35588 71540
rect 35532 71486 35534 71538
rect 35534 71486 35586 71538
rect 35586 71486 35588 71538
rect 35532 71484 35588 71486
rect 35196 71370 35252 71372
rect 35196 71318 35198 71370
rect 35198 71318 35250 71370
rect 35250 71318 35252 71370
rect 35196 71316 35252 71318
rect 35300 71370 35356 71372
rect 35300 71318 35302 71370
rect 35302 71318 35354 71370
rect 35354 71318 35356 71370
rect 35300 71316 35356 71318
rect 35404 71370 35460 71372
rect 35404 71318 35406 71370
rect 35406 71318 35458 71370
rect 35458 71318 35460 71370
rect 35404 71316 35460 71318
rect 35308 71036 35364 71092
rect 35420 70866 35476 70868
rect 35420 70814 35422 70866
rect 35422 70814 35474 70866
rect 35474 70814 35476 70866
rect 35420 70812 35476 70814
rect 35196 69802 35252 69804
rect 35196 69750 35198 69802
rect 35198 69750 35250 69802
rect 35250 69750 35252 69802
rect 35196 69748 35252 69750
rect 35300 69802 35356 69804
rect 35300 69750 35302 69802
rect 35302 69750 35354 69802
rect 35354 69750 35356 69802
rect 35300 69748 35356 69750
rect 35404 69802 35460 69804
rect 35404 69750 35406 69802
rect 35406 69750 35458 69802
rect 35458 69750 35460 69802
rect 35404 69748 35460 69750
rect 34972 68908 35028 68964
rect 35084 69356 35140 69412
rect 33404 65490 33460 65492
rect 33404 65438 33406 65490
rect 33406 65438 33458 65490
rect 33458 65438 33460 65490
rect 33404 65436 33460 65438
rect 32508 64876 32564 64932
rect 32620 64706 32676 64708
rect 32620 64654 32622 64706
rect 32622 64654 32674 64706
rect 32674 64654 32676 64706
rect 32620 64652 32676 64654
rect 32732 64316 32788 64372
rect 32508 64092 32564 64148
rect 32732 63980 32788 64036
rect 32620 63868 32676 63924
rect 32956 61964 33012 62020
rect 33180 61740 33236 61796
rect 33516 65378 33572 65380
rect 33516 65326 33518 65378
rect 33518 65326 33570 65378
rect 33570 65326 33572 65378
rect 33516 65324 33572 65326
rect 33852 65212 33908 65268
rect 33404 64876 33460 64932
rect 33292 61628 33348 61684
rect 33516 64034 33572 64036
rect 33516 63982 33518 64034
rect 33518 63982 33570 64034
rect 33570 63982 33572 64034
rect 33516 63980 33572 63982
rect 33180 61570 33236 61572
rect 33180 61518 33182 61570
rect 33182 61518 33234 61570
rect 33234 61518 33236 61570
rect 33180 61516 33236 61518
rect 33404 61404 33460 61460
rect 32844 60844 32900 60900
rect 31836 60172 31892 60228
rect 32172 60172 32228 60228
rect 32060 60114 32116 60116
rect 32060 60062 32062 60114
rect 32062 60062 32114 60114
rect 32114 60062 32116 60114
rect 32060 60060 32116 60062
rect 31724 59388 31780 59444
rect 31836 59948 31892 60004
rect 31836 58156 31892 58212
rect 33068 60226 33124 60228
rect 33068 60174 33070 60226
rect 33070 60174 33122 60226
rect 33122 60174 33124 60226
rect 33068 60172 33124 60174
rect 32956 60060 33012 60116
rect 32844 59388 32900 59444
rect 32396 59330 32452 59332
rect 32396 59278 32398 59330
rect 32398 59278 32450 59330
rect 32450 59278 32452 59330
rect 32396 59276 32452 59278
rect 32508 58716 32564 58772
rect 32956 58604 33012 58660
rect 32732 58546 32788 58548
rect 32732 58494 32734 58546
rect 32734 58494 32786 58546
rect 32786 58494 32788 58546
rect 32732 58492 32788 58494
rect 33292 60956 33348 61012
rect 34188 65490 34244 65492
rect 34188 65438 34190 65490
rect 34190 65438 34242 65490
rect 34242 65438 34244 65490
rect 34188 65436 34244 65438
rect 33852 63922 33908 63924
rect 33852 63870 33854 63922
rect 33854 63870 33906 63922
rect 33906 63870 33908 63922
rect 33852 63868 33908 63870
rect 33516 60844 33572 60900
rect 33628 61628 33684 61684
rect 33628 60732 33684 60788
rect 33740 61516 33796 61572
rect 36092 72322 36148 72324
rect 36092 72270 36094 72322
rect 36094 72270 36146 72322
rect 36146 72270 36148 72322
rect 36092 72268 36148 72270
rect 36764 72268 36820 72324
rect 36092 70140 36148 70196
rect 35868 69410 35924 69412
rect 35868 69358 35870 69410
rect 35870 69358 35922 69410
rect 35922 69358 35924 69410
rect 35868 69356 35924 69358
rect 35532 68796 35588 68852
rect 35196 68234 35252 68236
rect 35196 68182 35198 68234
rect 35198 68182 35250 68234
rect 35250 68182 35252 68234
rect 35196 68180 35252 68182
rect 35300 68234 35356 68236
rect 35300 68182 35302 68234
rect 35302 68182 35354 68234
rect 35354 68182 35356 68234
rect 35300 68180 35356 68182
rect 35404 68234 35460 68236
rect 35404 68182 35406 68234
rect 35406 68182 35458 68234
rect 35458 68182 35460 68234
rect 35404 68180 35460 68182
rect 35308 67228 35364 67284
rect 36092 67842 36148 67844
rect 36092 67790 36094 67842
rect 36094 67790 36146 67842
rect 36146 67790 36148 67842
rect 36092 67788 36148 67790
rect 36092 67618 36148 67620
rect 36092 67566 36094 67618
rect 36094 67566 36146 67618
rect 36146 67566 36148 67618
rect 36092 67564 36148 67566
rect 35196 66666 35252 66668
rect 35196 66614 35198 66666
rect 35198 66614 35250 66666
rect 35250 66614 35252 66666
rect 35196 66612 35252 66614
rect 35300 66666 35356 66668
rect 35300 66614 35302 66666
rect 35302 66614 35354 66666
rect 35354 66614 35356 66666
rect 35300 66612 35356 66614
rect 35404 66666 35460 66668
rect 35404 66614 35406 66666
rect 35406 66614 35458 66666
rect 35458 66614 35460 66666
rect 35404 66612 35460 66614
rect 34636 66386 34692 66388
rect 34636 66334 34638 66386
rect 34638 66334 34690 66386
rect 34690 66334 34692 66386
rect 34636 66332 34692 66334
rect 34748 66108 34804 66164
rect 34972 66108 35028 66164
rect 34300 64540 34356 64596
rect 34412 63980 34468 64036
rect 34636 65436 34692 65492
rect 35420 66220 35476 66276
rect 36316 71596 36372 71652
rect 36316 71036 36372 71092
rect 37212 71650 37268 71652
rect 37212 71598 37214 71650
rect 37214 71598 37266 71650
rect 37266 71598 37268 71650
rect 37212 71596 37268 71598
rect 37660 71650 37716 71652
rect 37660 71598 37662 71650
rect 37662 71598 37714 71650
rect 37714 71598 37716 71650
rect 37660 71596 37716 71598
rect 37212 70924 37268 70980
rect 38220 70588 38276 70644
rect 37324 70140 37380 70196
rect 36876 69916 36932 69972
rect 36764 67564 36820 67620
rect 37324 68908 37380 68964
rect 37884 68908 37940 68964
rect 37324 67954 37380 67956
rect 37324 67902 37326 67954
rect 37326 67902 37378 67954
rect 37378 67902 37380 67954
rect 37324 67900 37380 67902
rect 37212 67788 37268 67844
rect 36988 67228 37044 67284
rect 37436 67228 37492 67284
rect 36204 66220 36260 66276
rect 35196 65212 35252 65268
rect 35196 65098 35252 65100
rect 35196 65046 35198 65098
rect 35198 65046 35250 65098
rect 35250 65046 35252 65098
rect 35196 65044 35252 65046
rect 35300 65098 35356 65100
rect 35300 65046 35302 65098
rect 35302 65046 35354 65098
rect 35354 65046 35356 65098
rect 35300 65044 35356 65046
rect 35404 65098 35460 65100
rect 35404 65046 35406 65098
rect 35406 65046 35458 65098
rect 35458 65046 35460 65098
rect 35404 65044 35460 65046
rect 35868 65490 35924 65492
rect 35868 65438 35870 65490
rect 35870 65438 35922 65490
rect 35922 65438 35924 65490
rect 35868 65436 35924 65438
rect 35644 64988 35700 65044
rect 34860 64594 34916 64596
rect 34860 64542 34862 64594
rect 34862 64542 34914 64594
rect 34914 64542 34916 64594
rect 34860 64540 34916 64542
rect 33852 61180 33908 61236
rect 33852 60620 33908 60676
rect 33404 59778 33460 59780
rect 33404 59726 33406 59778
rect 33406 59726 33458 59778
rect 33458 59726 33460 59778
rect 33404 59724 33460 59726
rect 33292 59276 33348 59332
rect 33516 58492 33572 58548
rect 34188 60786 34244 60788
rect 34188 60734 34190 60786
rect 34190 60734 34242 60786
rect 34242 60734 34244 60786
rect 34188 60732 34244 60734
rect 33852 58716 33908 58772
rect 33964 58492 34020 58548
rect 34972 63084 35028 63140
rect 34748 60956 34804 61012
rect 34860 61964 34916 62020
rect 35196 63530 35252 63532
rect 35196 63478 35198 63530
rect 35198 63478 35250 63530
rect 35250 63478 35252 63530
rect 35196 63476 35252 63478
rect 35300 63530 35356 63532
rect 35300 63478 35302 63530
rect 35302 63478 35354 63530
rect 35354 63478 35356 63530
rect 35300 63476 35356 63478
rect 35404 63530 35460 63532
rect 35404 63478 35406 63530
rect 35406 63478 35458 63530
rect 35458 63478 35460 63530
rect 35404 63476 35460 63478
rect 35196 63308 35252 63364
rect 35868 64706 35924 64708
rect 35868 64654 35870 64706
rect 35870 64654 35922 64706
rect 35922 64654 35924 64706
rect 35868 64652 35924 64654
rect 35868 63868 35924 63924
rect 36764 65324 36820 65380
rect 36316 64818 36372 64820
rect 36316 64766 36318 64818
rect 36318 64766 36370 64818
rect 36370 64766 36372 64818
rect 36316 64764 36372 64766
rect 36204 64428 36260 64484
rect 36092 64092 36148 64148
rect 36428 63026 36484 63028
rect 36428 62974 36430 63026
rect 36430 62974 36482 63026
rect 36482 62974 36484 63026
rect 36428 62972 36484 62974
rect 36652 63308 36708 63364
rect 35084 62076 35140 62132
rect 37324 65324 37380 65380
rect 36988 64988 37044 65044
rect 36988 64818 37044 64820
rect 36988 64766 36990 64818
rect 36990 64766 37042 64818
rect 37042 64766 37044 64818
rect 36988 64764 37044 64766
rect 37100 64204 37156 64260
rect 35196 61962 35252 61964
rect 35196 61910 35198 61962
rect 35198 61910 35250 61962
rect 35250 61910 35252 61962
rect 35196 61908 35252 61910
rect 35300 61962 35356 61964
rect 35300 61910 35302 61962
rect 35302 61910 35354 61962
rect 35354 61910 35356 61962
rect 35300 61908 35356 61910
rect 35404 61962 35460 61964
rect 35404 61910 35406 61962
rect 35406 61910 35458 61962
rect 35458 61910 35460 61962
rect 35404 61908 35460 61910
rect 35308 61404 35364 61460
rect 34860 60508 34916 60564
rect 34412 59724 34468 59780
rect 35196 60394 35252 60396
rect 35196 60342 35198 60394
rect 35198 60342 35250 60394
rect 35250 60342 35252 60394
rect 35196 60340 35252 60342
rect 35300 60394 35356 60396
rect 35300 60342 35302 60394
rect 35302 60342 35354 60394
rect 35354 60342 35356 60394
rect 35300 60340 35356 60342
rect 35404 60394 35460 60396
rect 35404 60342 35406 60394
rect 35406 60342 35458 60394
rect 35458 60342 35460 60394
rect 35404 60340 35460 60342
rect 34860 59388 34916 59444
rect 35308 59276 35364 59332
rect 35532 59164 35588 59220
rect 34972 58940 35028 58996
rect 31948 56978 32004 56980
rect 31948 56926 31950 56978
rect 31950 56926 32002 56978
rect 32002 56926 32004 56978
rect 31948 56924 32004 56926
rect 34300 57484 34356 57540
rect 35196 58826 35252 58828
rect 35196 58774 35198 58826
rect 35198 58774 35250 58826
rect 35250 58774 35252 58826
rect 35196 58772 35252 58774
rect 35300 58826 35356 58828
rect 35300 58774 35302 58826
rect 35302 58774 35354 58826
rect 35354 58774 35356 58826
rect 35300 58772 35356 58774
rect 35404 58826 35460 58828
rect 35404 58774 35406 58826
rect 35406 58774 35458 58826
rect 35458 58774 35460 58826
rect 35404 58772 35460 58774
rect 35084 57484 35140 57540
rect 35196 57258 35252 57260
rect 35196 57206 35198 57258
rect 35198 57206 35250 57258
rect 35250 57206 35252 57258
rect 35196 57204 35252 57206
rect 35300 57258 35356 57260
rect 35300 57206 35302 57258
rect 35302 57206 35354 57258
rect 35354 57206 35356 57258
rect 35300 57204 35356 57206
rect 35404 57258 35460 57260
rect 35404 57206 35406 57258
rect 35406 57206 35458 57258
rect 35458 57206 35460 57258
rect 35404 57204 35460 57206
rect 35868 59724 35924 59780
rect 36316 59330 36372 59332
rect 36316 59278 36318 59330
rect 36318 59278 36370 59330
rect 36370 59278 36372 59330
rect 36316 59276 36372 59278
rect 36428 59218 36484 59220
rect 36428 59166 36430 59218
rect 36430 59166 36482 59218
rect 36482 59166 36484 59218
rect 36428 59164 36484 59166
rect 36204 58940 36260 58996
rect 35868 58604 35924 58660
rect 37324 64316 37380 64372
rect 37436 64540 37492 64596
rect 37548 65660 37604 65716
rect 37884 65212 37940 65268
rect 37548 63362 37604 63364
rect 37548 63310 37550 63362
rect 37550 63310 37602 63362
rect 37602 63310 37604 63362
rect 37548 63308 37604 63310
rect 37996 63868 38052 63924
rect 38220 64092 38276 64148
rect 37548 63138 37604 63140
rect 37548 63086 37550 63138
rect 37550 63086 37602 63138
rect 37602 63086 37604 63138
rect 37548 63084 37604 63086
rect 36988 61740 37044 61796
rect 37212 61292 37268 61348
rect 37100 60508 37156 60564
rect 36988 59724 37044 59780
rect 37212 59612 37268 59668
rect 37212 58604 37268 58660
rect 37660 62076 37716 62132
rect 37548 60956 37604 61012
rect 38220 62972 38276 63028
rect 38108 62076 38164 62132
rect 37884 61964 37940 62020
rect 37884 61740 37940 61796
rect 37772 61682 37828 61684
rect 37772 61630 37774 61682
rect 37774 61630 37826 61682
rect 37826 61630 37828 61682
rect 37772 61628 37828 61630
rect 37660 60508 37716 60564
rect 38108 61628 38164 61684
rect 37660 59612 37716 59668
rect 37884 59442 37940 59444
rect 37884 59390 37886 59442
rect 37886 59390 37938 59442
rect 37938 59390 37940 59442
rect 37884 59388 37940 59390
rect 37996 59330 38052 59332
rect 37996 59278 37998 59330
rect 37998 59278 38050 59330
rect 38050 59278 38052 59330
rect 37996 59276 38052 59278
rect 37772 58604 37828 58660
rect 38220 58268 38276 58324
rect 31836 56252 31892 56308
rect 35196 55690 35252 55692
rect 35196 55638 35198 55690
rect 35198 55638 35250 55690
rect 35250 55638 35252 55690
rect 35196 55636 35252 55638
rect 35300 55690 35356 55692
rect 35300 55638 35302 55690
rect 35302 55638 35354 55690
rect 35354 55638 35356 55690
rect 35300 55636 35356 55638
rect 35404 55690 35460 55692
rect 35404 55638 35406 55690
rect 35406 55638 35458 55690
rect 35458 55638 35460 55690
rect 35404 55636 35460 55638
rect 32284 55410 32340 55412
rect 32284 55358 32286 55410
rect 32286 55358 32338 55410
rect 32338 55358 32340 55410
rect 32284 55356 32340 55358
rect 32060 54348 32116 54404
rect 31836 53676 31892 53732
rect 31500 52780 31556 52836
rect 31388 52668 31444 52724
rect 31164 51324 31220 51380
rect 30716 49308 30772 49364
rect 30380 49196 30436 49252
rect 30604 48914 30660 48916
rect 30604 48862 30606 48914
rect 30606 48862 30658 48914
rect 30658 48862 30660 48914
rect 30604 48860 30660 48862
rect 30492 48076 30548 48132
rect 29932 46450 29988 46452
rect 29932 46398 29934 46450
rect 29934 46398 29986 46450
rect 29986 46398 29988 46450
rect 29932 46396 29988 46398
rect 31164 49196 31220 49252
rect 30828 47458 30884 47460
rect 30828 47406 30830 47458
rect 30830 47406 30882 47458
rect 30882 47406 30884 47458
rect 30828 47404 30884 47406
rect 31052 47404 31108 47460
rect 30940 47180 30996 47236
rect 30604 46396 30660 46452
rect 30492 46172 30548 46228
rect 30268 46060 30324 46116
rect 30604 46002 30660 46004
rect 30604 45950 30606 46002
rect 30606 45950 30658 46002
rect 30658 45950 30660 46002
rect 30604 45948 30660 45950
rect 30156 44380 30212 44436
rect 30828 44604 30884 44660
rect 30492 44492 30548 44548
rect 31724 48300 31780 48356
rect 31388 48130 31444 48132
rect 31388 48078 31390 48130
rect 31390 48078 31442 48130
rect 31442 48078 31444 48130
rect 31388 48076 31444 48078
rect 31836 47458 31892 47460
rect 31836 47406 31838 47458
rect 31838 47406 31890 47458
rect 31890 47406 31892 47458
rect 31836 47404 31892 47406
rect 31500 47346 31556 47348
rect 31500 47294 31502 47346
rect 31502 47294 31554 47346
rect 31554 47294 31556 47346
rect 31500 47292 31556 47294
rect 31164 46396 31220 46452
rect 31164 46060 31220 46116
rect 30940 44380 30996 44436
rect 30604 44210 30660 44212
rect 30604 44158 30606 44210
rect 30606 44158 30658 44210
rect 30658 44158 30660 44210
rect 30604 44156 30660 44158
rect 30828 44156 30884 44212
rect 30044 43260 30100 43316
rect 29932 42812 29988 42868
rect 30380 44098 30436 44100
rect 30380 44046 30382 44098
rect 30382 44046 30434 44098
rect 30434 44046 30436 44098
rect 30380 44044 30436 44046
rect 30716 43260 30772 43316
rect 30828 43372 30884 43428
rect 30604 42812 30660 42868
rect 29932 42140 29988 42196
rect 30380 42140 30436 42196
rect 30492 41970 30548 41972
rect 30492 41918 30494 41970
rect 30494 41918 30546 41970
rect 30546 41918 30548 41970
rect 30492 41916 30548 41918
rect 30940 43260 30996 43316
rect 30940 42978 30996 42980
rect 30940 42926 30942 42978
rect 30942 42926 30994 42978
rect 30994 42926 30996 42978
rect 30940 42924 30996 42926
rect 30828 42028 30884 42084
rect 30940 41692 30996 41748
rect 30940 41468 30996 41524
rect 30492 41356 30548 41412
rect 30044 40236 30100 40292
rect 28924 37490 28980 37492
rect 28924 37438 28926 37490
rect 28926 37438 28978 37490
rect 28978 37438 28980 37490
rect 28924 37436 28980 37438
rect 29148 37548 29204 37604
rect 28924 35810 28980 35812
rect 28924 35758 28926 35810
rect 28926 35758 28978 35810
rect 28978 35758 28980 35810
rect 28924 35756 28980 35758
rect 29148 35698 29204 35700
rect 29148 35646 29150 35698
rect 29150 35646 29202 35698
rect 29202 35646 29204 35698
rect 29148 35644 29204 35646
rect 30492 39788 30548 39844
rect 30268 36652 30324 36708
rect 30492 39228 30548 39284
rect 30604 38946 30660 38948
rect 30604 38894 30606 38946
rect 30606 38894 30658 38946
rect 30658 38894 30660 38946
rect 30604 38892 30660 38894
rect 30492 38780 30548 38836
rect 30716 38556 30772 38612
rect 30044 34524 30100 34580
rect 29484 33516 29540 33572
rect 29260 33292 29316 33348
rect 28812 32956 28868 33012
rect 31164 42924 31220 42980
rect 31388 43148 31444 43204
rect 31500 43036 31556 43092
rect 32060 46956 32116 47012
rect 31948 44604 32004 44660
rect 31948 42476 32004 42532
rect 31276 42082 31332 42084
rect 31276 42030 31278 42082
rect 31278 42030 31330 42082
rect 31330 42030 31332 42082
rect 31276 42028 31332 42030
rect 31500 41804 31556 41860
rect 31052 37436 31108 37492
rect 30604 35810 30660 35812
rect 30604 35758 30606 35810
rect 30606 35758 30658 35810
rect 30658 35758 30660 35810
rect 30604 35756 30660 35758
rect 31052 35922 31108 35924
rect 31052 35870 31054 35922
rect 31054 35870 31106 35922
rect 31106 35870 31108 35922
rect 31052 35868 31108 35870
rect 30268 34914 30324 34916
rect 30268 34862 30270 34914
rect 30270 34862 30322 34914
rect 30322 34862 30324 34914
rect 30268 34860 30324 34862
rect 30828 34860 30884 34916
rect 30156 34300 30212 34356
rect 31388 41580 31444 41636
rect 31500 41356 31556 41412
rect 31724 39676 31780 39732
rect 34860 55186 34916 55188
rect 34860 55134 34862 55186
rect 34862 55134 34914 55186
rect 34914 55134 34916 55186
rect 34860 55132 34916 55134
rect 35420 55132 35476 55188
rect 36428 55132 36484 55188
rect 32396 53730 32452 53732
rect 32396 53678 32398 53730
rect 32398 53678 32450 53730
rect 32450 53678 32452 53730
rect 32396 53676 32452 53678
rect 33852 53676 33908 53732
rect 33852 53116 33908 53172
rect 32284 52946 32340 52948
rect 32284 52894 32286 52946
rect 32286 52894 32338 52946
rect 32338 52894 32340 52946
rect 32284 52892 32340 52894
rect 33404 52722 33460 52724
rect 33404 52670 33406 52722
rect 33406 52670 33458 52722
rect 33458 52670 33460 52722
rect 33404 52668 33460 52670
rect 35196 54122 35252 54124
rect 35196 54070 35198 54122
rect 35198 54070 35250 54122
rect 35250 54070 35252 54122
rect 35196 54068 35252 54070
rect 35300 54122 35356 54124
rect 35300 54070 35302 54122
rect 35302 54070 35354 54122
rect 35354 54070 35356 54122
rect 35300 54068 35356 54070
rect 35404 54122 35460 54124
rect 35404 54070 35406 54122
rect 35406 54070 35458 54122
rect 35458 54070 35460 54122
rect 35404 54068 35460 54070
rect 34972 53170 35028 53172
rect 34972 53118 34974 53170
rect 34974 53118 35026 53170
rect 35026 53118 35028 53170
rect 34972 53116 35028 53118
rect 34076 52668 34132 52724
rect 35308 52834 35364 52836
rect 35308 52782 35310 52834
rect 35310 52782 35362 52834
rect 35362 52782 35364 52834
rect 35308 52780 35364 52782
rect 35196 52554 35252 52556
rect 35196 52502 35198 52554
rect 35198 52502 35250 52554
rect 35250 52502 35252 52554
rect 35196 52500 35252 52502
rect 35300 52554 35356 52556
rect 35300 52502 35302 52554
rect 35302 52502 35354 52554
rect 35354 52502 35356 52554
rect 35300 52500 35356 52502
rect 35404 52554 35460 52556
rect 35404 52502 35406 52554
rect 35406 52502 35458 52554
rect 35458 52502 35460 52554
rect 35404 52500 35460 52502
rect 35644 52668 35700 52724
rect 35644 52108 35700 52164
rect 35196 50986 35252 50988
rect 35196 50934 35198 50986
rect 35198 50934 35250 50986
rect 35250 50934 35252 50986
rect 35196 50932 35252 50934
rect 35300 50986 35356 50988
rect 35300 50934 35302 50986
rect 35302 50934 35354 50986
rect 35354 50934 35356 50986
rect 35300 50932 35356 50934
rect 35404 50986 35460 50988
rect 35404 50934 35406 50986
rect 35406 50934 35458 50986
rect 35458 50934 35460 50986
rect 35404 50932 35460 50934
rect 34748 50316 34804 50372
rect 33740 49196 33796 49252
rect 34188 48860 34244 48916
rect 33852 48466 33908 48468
rect 33852 48414 33854 48466
rect 33854 48414 33906 48466
rect 33906 48414 33908 48466
rect 33852 48412 33908 48414
rect 34972 49810 35028 49812
rect 34972 49758 34974 49810
rect 34974 49758 35026 49810
rect 35026 49758 35028 49810
rect 34972 49756 35028 49758
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 36316 52162 36372 52164
rect 36316 52110 36318 52162
rect 36318 52110 36370 52162
rect 36370 52110 36372 52162
rect 36316 52108 36372 52110
rect 35644 49756 35700 49812
rect 35756 51996 35812 52052
rect 34860 48748 34916 48804
rect 35196 48802 35252 48804
rect 35196 48750 35198 48802
rect 35198 48750 35250 48802
rect 35250 48750 35252 48802
rect 35196 48748 35252 48750
rect 34748 48466 34804 48468
rect 34748 48414 34750 48466
rect 34750 48414 34802 48466
rect 34802 48414 34804 48466
rect 34748 48412 34804 48414
rect 32284 48130 32340 48132
rect 32284 48078 32286 48130
rect 32286 48078 32338 48130
rect 32338 48078 32340 48130
rect 32284 48076 32340 48078
rect 32620 47346 32676 47348
rect 32620 47294 32622 47346
rect 32622 47294 32674 47346
rect 32674 47294 32676 47346
rect 32620 47292 32676 47294
rect 33180 46956 33236 47012
rect 33404 46898 33460 46900
rect 33404 46846 33406 46898
rect 33406 46846 33458 46898
rect 33458 46846 33460 46898
rect 33404 46844 33460 46846
rect 32396 44322 32452 44324
rect 32396 44270 32398 44322
rect 32398 44270 32450 44322
rect 32450 44270 32452 44322
rect 32396 44268 32452 44270
rect 32844 44098 32900 44100
rect 32844 44046 32846 44098
rect 32846 44046 32898 44098
rect 32898 44046 32900 44098
rect 32844 44044 32900 44046
rect 33180 43596 33236 43652
rect 32284 43036 32340 43092
rect 33068 43372 33124 43428
rect 32396 42476 32452 42532
rect 33180 42476 33236 42532
rect 32284 41858 32340 41860
rect 32284 41806 32286 41858
rect 32286 41806 32338 41858
rect 32338 41806 32340 41858
rect 32284 41804 32340 41806
rect 32172 41356 32228 41412
rect 32732 41244 32788 41300
rect 32508 39730 32564 39732
rect 32508 39678 32510 39730
rect 32510 39678 32562 39730
rect 32562 39678 32564 39730
rect 32508 39676 32564 39678
rect 31948 39564 32004 39620
rect 33180 39618 33236 39620
rect 33180 39566 33182 39618
rect 33182 39566 33234 39618
rect 33234 39566 33236 39618
rect 33180 39564 33236 39566
rect 31388 38668 31444 38724
rect 33740 39618 33796 39620
rect 33740 39566 33742 39618
rect 33742 39566 33794 39618
rect 33794 39566 33796 39618
rect 33740 39564 33796 39566
rect 33180 38892 33236 38948
rect 32172 38834 32228 38836
rect 32172 38782 32174 38834
rect 32174 38782 32226 38834
rect 32226 38782 32228 38834
rect 32172 38780 32228 38782
rect 31836 38668 31892 38724
rect 34076 47516 34132 47572
rect 34748 47570 34804 47572
rect 34748 47518 34750 47570
rect 34750 47518 34802 47570
rect 34802 47518 34804 47570
rect 34748 47516 34804 47518
rect 35532 48636 35588 48692
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 35532 47628 35588 47684
rect 35084 46898 35140 46900
rect 35084 46846 35086 46898
rect 35086 46846 35138 46898
rect 35138 46846 35140 46898
rect 35084 46844 35140 46846
rect 35308 46396 35364 46452
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 34972 45666 35028 45668
rect 34972 45614 34974 45666
rect 34974 45614 35026 45666
rect 35026 45614 35028 45666
rect 34972 45612 35028 45614
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 34972 43596 35028 43652
rect 34636 43426 34692 43428
rect 34636 43374 34638 43426
rect 34638 43374 34690 43426
rect 34690 43374 34692 43426
rect 34636 43372 34692 43374
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 36204 48636 36260 48692
rect 36204 47628 36260 47684
rect 36204 47292 36260 47348
rect 35532 42924 35588 42980
rect 35644 44044 35700 44100
rect 34524 42700 34580 42756
rect 35308 42140 35364 42196
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 35868 43596 35924 43652
rect 35868 42812 35924 42868
rect 35308 41298 35364 41300
rect 35308 41246 35310 41298
rect 35310 41246 35362 41298
rect 35362 41246 35364 41298
rect 35308 41244 35364 41246
rect 35420 40572 35476 40628
rect 34972 40236 35028 40292
rect 34300 39842 34356 39844
rect 34300 39790 34302 39842
rect 34302 39790 34354 39842
rect 34354 39790 34356 39842
rect 34300 39788 34356 39790
rect 35756 41244 35812 41300
rect 36092 41298 36148 41300
rect 36092 41246 36094 41298
rect 36094 41246 36146 41298
rect 36146 41246 36148 41298
rect 36092 41244 36148 41246
rect 37548 51996 37604 52052
rect 38108 51996 38164 52052
rect 37884 50316 37940 50372
rect 36988 47346 37044 47348
rect 36988 47294 36990 47346
rect 36990 47294 37042 47346
rect 37042 47294 37044 47346
rect 36988 47292 37044 47294
rect 37548 47570 37604 47572
rect 37548 47518 37550 47570
rect 37550 47518 37602 47570
rect 37602 47518 37604 47570
rect 37548 47516 37604 47518
rect 36428 46732 36484 46788
rect 37212 46956 37268 47012
rect 36988 46396 37044 46452
rect 37436 46786 37492 46788
rect 37436 46734 37438 46786
rect 37438 46734 37490 46786
rect 37490 46734 37492 46786
rect 37436 46732 37492 46734
rect 36428 42866 36484 42868
rect 36428 42814 36430 42866
rect 36430 42814 36482 42866
rect 36482 42814 36484 42866
rect 36428 42812 36484 42814
rect 36428 42588 36484 42644
rect 35644 40236 35700 40292
rect 35532 40124 35588 40180
rect 31612 38556 31668 38612
rect 31164 35196 31220 35252
rect 29260 31948 29316 32004
rect 30044 31948 30100 32004
rect 30492 30882 30548 30884
rect 30492 30830 30494 30882
rect 30494 30830 30546 30882
rect 30546 30830 30548 30882
rect 30492 30828 30548 30830
rect 29820 30098 29876 30100
rect 29820 30046 29822 30098
rect 29822 30046 29874 30098
rect 29874 30046 29876 30098
rect 29820 30044 29876 30046
rect 29820 29372 29876 29428
rect 27804 29202 27860 29204
rect 27804 29150 27806 29202
rect 27806 29150 27858 29202
rect 27858 29150 27860 29202
rect 27804 29148 27860 29150
rect 29260 28028 29316 28084
rect 27468 27468 27524 27524
rect 28028 27468 28084 27524
rect 26908 26908 26964 26964
rect 26572 26684 26628 26740
rect 26460 26236 26516 26292
rect 26572 26460 26628 26516
rect 26348 25618 26404 25620
rect 26348 25566 26350 25618
rect 26350 25566 26402 25618
rect 26402 25566 26404 25618
rect 26348 25564 26404 25566
rect 26124 25394 26180 25396
rect 26124 25342 26126 25394
rect 26126 25342 26178 25394
rect 26178 25342 26180 25394
rect 26124 25340 26180 25342
rect 25564 23938 25620 23940
rect 25564 23886 25566 23938
rect 25566 23886 25618 23938
rect 25618 23886 25620 23938
rect 25564 23884 25620 23886
rect 25676 23772 25732 23828
rect 25564 23492 25620 23548
rect 25228 23042 25284 23044
rect 25228 22990 25230 23042
rect 25230 22990 25282 23042
rect 25282 22990 25284 23042
rect 25228 22988 25284 22990
rect 26012 22988 26068 23044
rect 25564 17778 25620 17780
rect 25564 17726 25566 17778
rect 25566 17726 25618 17778
rect 25618 17726 25620 17778
rect 25564 17724 25620 17726
rect 24220 15426 24276 15428
rect 24220 15374 24222 15426
rect 24222 15374 24274 15426
rect 24274 15374 24276 15426
rect 24220 15372 24276 15374
rect 24108 15314 24164 15316
rect 24108 15262 24110 15314
rect 24110 15262 24162 15314
rect 24162 15262 24164 15314
rect 24108 15260 24164 15262
rect 24556 13186 24612 13188
rect 24556 13134 24558 13186
rect 24558 13134 24610 13186
rect 24610 13134 24612 13186
rect 24556 13132 24612 13134
rect 26236 17052 26292 17108
rect 25676 16716 25732 16772
rect 25340 15372 25396 15428
rect 26012 15484 26068 15540
rect 23772 12236 23828 12292
rect 24220 12290 24276 12292
rect 24220 12238 24222 12290
rect 24222 12238 24274 12290
rect 24274 12238 24276 12290
rect 24220 12236 24276 12238
rect 21868 10108 21924 10164
rect 21756 9548 21812 9604
rect 20412 7308 20468 7364
rect 20188 5292 20244 5348
rect 20412 6636 20468 6692
rect 19740 5234 19796 5236
rect 19740 5182 19742 5234
rect 19742 5182 19794 5234
rect 19794 5182 19796 5234
rect 19740 5180 19796 5182
rect 20412 5180 20468 5236
rect 21308 6636 21364 6692
rect 24220 10834 24276 10836
rect 24220 10782 24222 10834
rect 24222 10782 24274 10834
rect 24274 10782 24276 10834
rect 24220 10780 24276 10782
rect 22204 5516 22260 5572
rect 22316 5852 22372 5908
rect 21532 5346 21588 5348
rect 21532 5294 21534 5346
rect 21534 5294 21586 5346
rect 21586 5294 21588 5346
rect 21532 5292 21588 5294
rect 23212 5852 23268 5908
rect 24220 5906 24276 5908
rect 24220 5854 24222 5906
rect 24222 5854 24274 5906
rect 24274 5854 24276 5906
rect 24220 5852 24276 5854
rect 25228 13132 25284 13188
rect 25116 12236 25172 12292
rect 25228 12124 25284 12180
rect 24668 10610 24724 10612
rect 24668 10558 24670 10610
rect 24670 10558 24722 10610
rect 24722 10558 24724 10610
rect 24668 10556 24724 10558
rect 26460 15426 26516 15428
rect 26460 15374 26462 15426
rect 26462 15374 26514 15426
rect 26514 15374 26516 15426
rect 26460 15372 26516 15374
rect 27132 26348 27188 26404
rect 26684 25282 26740 25284
rect 26684 25230 26686 25282
rect 26686 25230 26738 25282
rect 26738 25230 26740 25282
rect 26684 25228 26740 25230
rect 27020 25228 27076 25284
rect 26796 25116 26852 25172
rect 26684 20578 26740 20580
rect 26684 20526 26686 20578
rect 26686 20526 26738 20578
rect 26738 20526 26740 20578
rect 26684 20524 26740 20526
rect 26684 19964 26740 20020
rect 26684 19234 26740 19236
rect 26684 19182 26686 19234
rect 26686 19182 26738 19234
rect 26738 19182 26740 19234
rect 26684 19180 26740 19182
rect 26684 16940 26740 16996
rect 27020 24722 27076 24724
rect 27020 24670 27022 24722
rect 27022 24670 27074 24722
rect 27074 24670 27076 24722
rect 27020 24668 27076 24670
rect 27804 25676 27860 25732
rect 27804 25282 27860 25284
rect 27804 25230 27806 25282
rect 27806 25230 27858 25282
rect 27858 25230 27860 25282
rect 27804 25228 27860 25230
rect 27916 23324 27972 23380
rect 28028 23212 28084 23268
rect 29260 27468 29316 27524
rect 30044 28812 30100 28868
rect 30156 28028 30212 28084
rect 30380 26962 30436 26964
rect 30380 26910 30382 26962
rect 30382 26910 30434 26962
rect 30434 26910 30436 26962
rect 30380 26908 30436 26910
rect 30492 25228 30548 25284
rect 30268 25116 30324 25172
rect 29708 24668 29764 24724
rect 29708 23938 29764 23940
rect 29708 23886 29710 23938
rect 29710 23886 29762 23938
rect 29762 23886 29764 23938
rect 29708 23884 29764 23886
rect 29820 23996 29876 24052
rect 29148 23436 29204 23492
rect 28588 23266 28644 23268
rect 28588 23214 28590 23266
rect 28590 23214 28642 23266
rect 28642 23214 28644 23266
rect 28588 23212 28644 23214
rect 27244 20524 27300 20580
rect 27132 19180 27188 19236
rect 27692 17724 27748 17780
rect 26908 17106 26964 17108
rect 26908 17054 26910 17106
rect 26910 17054 26962 17106
rect 26962 17054 26964 17106
rect 26908 17052 26964 17054
rect 27692 16940 27748 16996
rect 26796 16716 26852 16772
rect 29260 23378 29316 23380
rect 29260 23326 29262 23378
rect 29262 23326 29314 23378
rect 29314 23326 29316 23378
rect 29260 23324 29316 23326
rect 29596 21474 29652 21476
rect 29596 21422 29598 21474
rect 29598 21422 29650 21474
rect 29650 21422 29652 21474
rect 29596 21420 29652 21422
rect 29260 20524 29316 20580
rect 29708 19404 29764 19460
rect 29260 19346 29316 19348
rect 29260 19294 29262 19346
rect 29262 19294 29314 19346
rect 29314 19294 29316 19346
rect 29260 19292 29316 19294
rect 28028 15820 28084 15876
rect 28588 17724 28644 17780
rect 29260 17724 29316 17780
rect 30044 17778 30100 17780
rect 30044 17726 30046 17778
rect 30046 17726 30098 17778
rect 30098 17726 30100 17778
rect 30044 17724 30100 17726
rect 30492 23826 30548 23828
rect 30492 23774 30494 23826
rect 30494 23774 30546 23826
rect 30546 23774 30548 23826
rect 30492 23772 30548 23774
rect 31836 36204 31892 36260
rect 31612 34802 31668 34804
rect 31612 34750 31614 34802
rect 31614 34750 31666 34802
rect 31666 34750 31668 34802
rect 31612 34748 31668 34750
rect 31500 34130 31556 34132
rect 31500 34078 31502 34130
rect 31502 34078 31554 34130
rect 31554 34078 31556 34130
rect 31500 34076 31556 34078
rect 31500 33516 31556 33572
rect 31500 33346 31556 33348
rect 31500 33294 31502 33346
rect 31502 33294 31554 33346
rect 31554 33294 31556 33346
rect 31500 33292 31556 33294
rect 30940 32284 30996 32340
rect 30716 30828 30772 30884
rect 31948 34524 32004 34580
rect 31948 34354 32004 34356
rect 31948 34302 31950 34354
rect 31950 34302 32002 34354
rect 32002 34302 32004 34354
rect 31948 34300 32004 34302
rect 31836 32620 31892 32676
rect 32172 35532 32228 35588
rect 32172 33516 32228 33572
rect 31612 30828 31668 30884
rect 30828 30098 30884 30100
rect 30828 30046 30830 30098
rect 30830 30046 30882 30098
rect 30882 30046 30884 30098
rect 30828 30044 30884 30046
rect 30716 29596 30772 29652
rect 30716 28866 30772 28868
rect 30716 28814 30718 28866
rect 30718 28814 30770 28866
rect 30770 28814 30772 28866
rect 30716 28812 30772 28814
rect 31612 30210 31668 30212
rect 31612 30158 31614 30210
rect 31614 30158 31666 30210
rect 31666 30158 31668 30210
rect 31612 30156 31668 30158
rect 32060 30044 32116 30100
rect 31276 29596 31332 29652
rect 31164 28812 31220 28868
rect 30716 28082 30772 28084
rect 30716 28030 30718 28082
rect 30718 28030 30770 28082
rect 30770 28030 30772 28082
rect 30716 28028 30772 28030
rect 31500 27746 31556 27748
rect 31500 27694 31502 27746
rect 31502 27694 31554 27746
rect 31554 27694 31556 27746
rect 31500 27692 31556 27694
rect 32396 35756 32452 35812
rect 33404 37772 33460 37828
rect 32844 36258 32900 36260
rect 32844 36206 32846 36258
rect 32846 36206 32898 36258
rect 32898 36206 32900 36258
rect 32844 36204 32900 36206
rect 32956 35532 33012 35588
rect 32844 35420 32900 35476
rect 32732 34802 32788 34804
rect 32732 34750 32734 34802
rect 32734 34750 32786 34802
rect 32786 34750 32788 34802
rect 32732 34748 32788 34750
rect 33404 34354 33460 34356
rect 33404 34302 33406 34354
rect 33406 34302 33458 34354
rect 33458 34302 33460 34354
rect 33404 34300 33460 34302
rect 33068 33570 33124 33572
rect 33068 33518 33070 33570
rect 33070 33518 33122 33570
rect 33122 33518 33124 33570
rect 33068 33516 33124 33518
rect 33852 37826 33908 37828
rect 33852 37774 33854 37826
rect 33854 37774 33906 37826
rect 33906 37774 33908 37826
rect 33852 37772 33908 37774
rect 33852 36988 33908 37044
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 35196 39676 35252 39732
rect 35308 39618 35364 39620
rect 35308 39566 35310 39618
rect 35310 39566 35362 39618
rect 35362 39566 35364 39618
rect 35308 39564 35364 39566
rect 35756 39730 35812 39732
rect 35756 39678 35758 39730
rect 35758 39678 35810 39730
rect 35810 39678 35812 39730
rect 35756 39676 35812 39678
rect 36092 40572 36148 40628
rect 36204 40124 36260 40180
rect 35532 39116 35588 39172
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 35308 37154 35364 37156
rect 35308 37102 35310 37154
rect 35310 37102 35362 37154
rect 35362 37102 35364 37154
rect 35308 37100 35364 37102
rect 36428 39564 36484 39620
rect 36428 38050 36484 38052
rect 36428 37998 36430 38050
rect 36430 37998 36482 38050
rect 36482 37998 36484 38050
rect 36428 37996 36484 37998
rect 35868 37100 35924 37156
rect 36428 37100 36484 37156
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 33740 35196 33796 35252
rect 33740 34748 33796 34804
rect 34076 34860 34132 34916
rect 34076 34354 34132 34356
rect 34076 34302 34078 34354
rect 34078 34302 34130 34354
rect 34130 34302 34132 34354
rect 34076 34300 34132 34302
rect 34524 34636 34580 34692
rect 32396 30882 32452 30884
rect 32396 30830 32398 30882
rect 32398 30830 32450 30882
rect 32450 30830 32452 30882
rect 32396 30828 32452 30830
rect 33068 32674 33124 32676
rect 33068 32622 33070 32674
rect 33070 32622 33122 32674
rect 33122 32622 33124 32674
rect 33068 32620 33124 32622
rect 34300 33404 34356 33460
rect 33852 31948 33908 32004
rect 32956 30828 33012 30884
rect 33516 30828 33572 30884
rect 32732 30210 32788 30212
rect 32732 30158 32734 30210
rect 32734 30158 32786 30210
rect 32786 30158 32788 30210
rect 32732 30156 32788 30158
rect 32508 30098 32564 30100
rect 32508 30046 32510 30098
rect 32510 30046 32562 30098
rect 32562 30046 32564 30098
rect 32508 30044 32564 30046
rect 31388 26962 31444 26964
rect 31388 26910 31390 26962
rect 31390 26910 31442 26962
rect 31442 26910 31444 26962
rect 31388 26908 31444 26910
rect 31052 25282 31108 25284
rect 31052 25230 31054 25282
rect 31054 25230 31106 25282
rect 31106 25230 31108 25282
rect 31052 25228 31108 25230
rect 33852 29596 33908 29652
rect 32844 28028 32900 28084
rect 32508 27692 32564 27748
rect 35532 36652 35588 36708
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35644 35196 35700 35252
rect 35756 35756 35812 35812
rect 35084 34860 35140 34916
rect 35420 34972 35476 35028
rect 35196 34242 35252 34244
rect 35196 34190 35198 34242
rect 35198 34190 35250 34242
rect 35250 34190 35252 34242
rect 35196 34188 35252 34190
rect 35644 35026 35700 35028
rect 35644 34974 35646 35026
rect 35646 34974 35698 35026
rect 35698 34974 35700 35026
rect 35644 34972 35700 34974
rect 35532 34802 35588 34804
rect 35532 34750 35534 34802
rect 35534 34750 35586 34802
rect 35586 34750 35588 34802
rect 35532 34748 35588 34750
rect 36092 35586 36148 35588
rect 36092 35534 36094 35586
rect 36094 35534 36146 35586
rect 36146 35534 36148 35586
rect 36092 35532 36148 35534
rect 35980 35308 36036 35364
rect 35868 34914 35924 34916
rect 35868 34862 35870 34914
rect 35870 34862 35922 34914
rect 35922 34862 35924 34914
rect 35868 34860 35924 34862
rect 35644 34300 35700 34356
rect 35532 34018 35588 34020
rect 35532 33966 35534 34018
rect 35534 33966 35586 34018
rect 35586 33966 35588 34018
rect 35532 33964 35588 33966
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 34860 33404 34916 33460
rect 35308 33458 35364 33460
rect 35308 33406 35310 33458
rect 35310 33406 35362 33458
rect 35362 33406 35364 33458
rect 35308 33404 35364 33406
rect 34972 33346 35028 33348
rect 34972 33294 34974 33346
rect 34974 33294 35026 33346
rect 35026 33294 35028 33346
rect 34972 33292 35028 33294
rect 35532 33346 35588 33348
rect 35532 33294 35534 33346
rect 35534 33294 35586 33346
rect 35586 33294 35588 33346
rect 35532 33292 35588 33294
rect 36204 34300 36260 34356
rect 36428 35420 36484 35476
rect 36204 33964 36260 34020
rect 36092 33292 36148 33348
rect 35868 33234 35924 33236
rect 35868 33182 35870 33234
rect 35870 33182 35922 33234
rect 35922 33182 35924 33234
rect 35868 33180 35924 33182
rect 35084 32284 35140 32340
rect 35868 32284 35924 32340
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35644 31948 35700 32004
rect 36204 31666 36260 31668
rect 36204 31614 36206 31666
rect 36206 31614 36258 31666
rect 36258 31614 36260 31666
rect 36204 31612 36260 31614
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 34748 29596 34804 29652
rect 35308 29314 35364 29316
rect 35308 29262 35310 29314
rect 35310 29262 35362 29314
rect 35362 29262 35364 29314
rect 35308 29260 35364 29262
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 35308 27244 35364 27300
rect 31164 25116 31220 25172
rect 31500 25282 31556 25284
rect 31500 25230 31502 25282
rect 31502 25230 31554 25282
rect 31554 25230 31556 25282
rect 31500 25228 31556 25230
rect 30828 24610 30884 24612
rect 30828 24558 30830 24610
rect 30830 24558 30882 24610
rect 30882 24558 30884 24610
rect 30828 24556 30884 24558
rect 31500 24668 31556 24724
rect 31388 24556 31444 24612
rect 33404 24834 33460 24836
rect 33404 24782 33406 24834
rect 33406 24782 33458 24834
rect 33458 24782 33460 24834
rect 33404 24780 33460 24782
rect 32060 24722 32116 24724
rect 32060 24670 32062 24722
rect 32062 24670 32114 24722
rect 32114 24670 32116 24722
rect 32060 24668 32116 24670
rect 31836 24332 31892 24388
rect 32172 23996 32228 24052
rect 32620 24332 32676 24388
rect 32956 24050 33012 24052
rect 32956 23998 32958 24050
rect 32958 23998 33010 24050
rect 33010 23998 33012 24050
rect 32956 23996 33012 23998
rect 31164 23772 31220 23828
rect 33180 23884 33236 23940
rect 30492 19404 30548 19460
rect 32508 21586 32564 21588
rect 32508 21534 32510 21586
rect 32510 21534 32562 21586
rect 32562 21534 32564 21586
rect 32508 21532 32564 21534
rect 31836 21308 31892 21364
rect 33068 21362 33124 21364
rect 33068 21310 33070 21362
rect 33070 21310 33122 21362
rect 33122 21310 33124 21362
rect 33068 21308 33124 21310
rect 32732 20578 32788 20580
rect 32732 20526 32734 20578
rect 32734 20526 32786 20578
rect 32786 20526 32788 20578
rect 32732 20524 32788 20526
rect 33404 20524 33460 20580
rect 32844 19404 32900 19460
rect 30828 19292 30884 19348
rect 32396 19346 32452 19348
rect 32396 19294 32398 19346
rect 32398 19294 32450 19346
rect 32450 19294 32452 19346
rect 32396 19292 32452 19294
rect 33628 19852 33684 19908
rect 33740 19964 33796 20020
rect 33292 19292 33348 19348
rect 33628 19404 33684 19460
rect 36204 27186 36260 27188
rect 36204 27134 36206 27186
rect 36206 27134 36258 27186
rect 36258 27134 36260 27186
rect 36204 27132 36260 27134
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 35420 25394 35476 25396
rect 35420 25342 35422 25394
rect 35422 25342 35474 25394
rect 35474 25342 35476 25394
rect 35420 25340 35476 25342
rect 35868 25340 35924 25396
rect 35084 24780 35140 24836
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 34636 23884 34692 23940
rect 35756 23938 35812 23940
rect 35756 23886 35758 23938
rect 35758 23886 35810 23938
rect 35810 23886 35812 23938
rect 35756 23884 35812 23886
rect 34972 23436 35028 23492
rect 34076 19964 34132 20020
rect 34188 22876 34244 22932
rect 34972 23154 35028 23156
rect 34972 23102 34974 23154
rect 34974 23102 35026 23154
rect 35026 23102 35028 23154
rect 34972 23100 35028 23102
rect 34524 21586 34580 21588
rect 34524 21534 34526 21586
rect 34526 21534 34578 21586
rect 34578 21534 34580 21586
rect 34524 21532 34580 21534
rect 35532 23154 35588 23156
rect 35532 23102 35534 23154
rect 35534 23102 35586 23154
rect 35586 23102 35588 23154
rect 35532 23100 35588 23102
rect 35196 22876 35252 22932
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 34188 20188 34244 20244
rect 34860 20524 34916 20580
rect 34636 20130 34692 20132
rect 34636 20078 34638 20130
rect 34638 20078 34690 20130
rect 34690 20078 34692 20130
rect 34636 20076 34692 20078
rect 34076 19292 34132 19348
rect 34524 20018 34580 20020
rect 34524 19966 34526 20018
rect 34526 19966 34578 20018
rect 34578 19966 34580 20018
rect 34524 19964 34580 19966
rect 34748 20018 34804 20020
rect 34748 19966 34750 20018
rect 34750 19966 34802 20018
rect 34802 19966 34804 20018
rect 34748 19964 34804 19966
rect 34972 20188 35028 20244
rect 35532 19964 35588 20020
rect 35308 19906 35364 19908
rect 35308 19854 35310 19906
rect 35310 19854 35362 19906
rect 35362 19854 35364 19906
rect 35308 19852 35364 19854
rect 30492 18338 30548 18340
rect 30492 18286 30494 18338
rect 30494 18286 30546 18338
rect 30546 18286 30548 18338
rect 30492 18284 30548 18286
rect 30828 18338 30884 18340
rect 30828 18286 30830 18338
rect 30830 18286 30882 18338
rect 30882 18286 30884 18338
rect 30828 18284 30884 18286
rect 30492 17724 30548 17780
rect 30268 17052 30324 17108
rect 26460 14924 26516 14980
rect 25340 10834 25396 10836
rect 25340 10782 25342 10834
rect 25342 10782 25394 10834
rect 25394 10782 25396 10834
rect 25340 10780 25396 10782
rect 25676 10610 25732 10612
rect 25676 10558 25678 10610
rect 25678 10558 25730 10610
rect 25730 10558 25732 10610
rect 25676 10556 25732 10558
rect 26236 11452 26292 11508
rect 27020 14924 27076 14980
rect 26012 10556 26068 10612
rect 28700 16716 28756 16772
rect 28700 16044 28756 16100
rect 29708 16098 29764 16100
rect 29708 16046 29710 16098
rect 29710 16046 29762 16098
rect 29762 16046 29764 16098
rect 29708 16044 29764 16046
rect 29484 14924 29540 14980
rect 29036 13580 29092 13636
rect 30044 13580 30100 13636
rect 28588 12124 28644 12180
rect 29708 12178 29764 12180
rect 29708 12126 29710 12178
rect 29710 12126 29762 12178
rect 29762 12126 29764 12178
rect 29708 12124 29764 12126
rect 28028 12012 28084 12068
rect 26348 10780 26404 10836
rect 26796 11228 26852 11284
rect 26348 9996 26404 10052
rect 26460 9938 26516 9940
rect 26460 9886 26462 9938
rect 26462 9886 26514 9938
rect 26514 9886 26516 9938
rect 26460 9884 26516 9886
rect 26684 9884 26740 9940
rect 26908 10610 26964 10612
rect 26908 10558 26910 10610
rect 26910 10558 26962 10610
rect 26962 10558 26964 10610
rect 26908 10556 26964 10558
rect 27468 10556 27524 10612
rect 28924 12066 28980 12068
rect 28924 12014 28926 12066
rect 28926 12014 28978 12066
rect 28978 12014 28980 12066
rect 28924 12012 28980 12014
rect 25452 8428 25508 8484
rect 25564 8258 25620 8260
rect 25564 8206 25566 8258
rect 25566 8206 25618 8258
rect 25618 8206 25620 8258
rect 25564 8204 25620 8206
rect 25116 8034 25172 8036
rect 25116 7982 25118 8034
rect 25118 7982 25170 8034
rect 25170 7982 25172 8034
rect 25116 7980 25172 7982
rect 24892 5852 24948 5908
rect 22316 5292 22372 5348
rect 23100 5404 23156 5460
rect 23324 5180 23380 5236
rect 20076 4898 20132 4900
rect 20076 4846 20078 4898
rect 20078 4846 20130 4898
rect 20130 4846 20132 4898
rect 20076 4844 20132 4846
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 25564 6636 25620 6692
rect 25564 5906 25620 5908
rect 25564 5854 25566 5906
rect 25566 5854 25618 5906
rect 25618 5854 25620 5906
rect 25564 5852 25620 5854
rect 26348 7980 26404 8036
rect 27020 8258 27076 8260
rect 27020 8206 27022 8258
rect 27022 8206 27074 8258
rect 27074 8206 27076 8258
rect 27020 8204 27076 8206
rect 27244 8204 27300 8260
rect 26908 7586 26964 7588
rect 26908 7534 26910 7586
rect 26910 7534 26962 7586
rect 26962 7534 26964 7586
rect 26908 7532 26964 7534
rect 26572 7308 26628 7364
rect 25116 5404 25172 5460
rect 24220 5180 24276 5236
rect 24444 5068 24500 5124
rect 14476 2492 14532 2548
rect 15148 3276 15204 3332
rect 15260 2882 15316 2884
rect 15260 2830 15262 2882
rect 15262 2830 15314 2882
rect 15314 2830 15316 2882
rect 15260 2828 15316 2830
rect 16156 3330 16212 3332
rect 16156 3278 16158 3330
rect 16158 3278 16210 3330
rect 16210 3278 16212 3330
rect 16156 3276 16212 3278
rect 16380 2940 16436 2996
rect 16380 2716 16436 2772
rect 17612 2770 17668 2772
rect 17612 2718 17614 2770
rect 17614 2718 17666 2770
rect 17666 2718 17668 2770
rect 17612 2716 17668 2718
rect 17836 3388 17892 3444
rect 17276 1762 17332 1764
rect 17276 1710 17278 1762
rect 17278 1710 17330 1762
rect 17330 1710 17332 1762
rect 17276 1708 17332 1710
rect 18172 2770 18228 2772
rect 18172 2718 18174 2770
rect 18174 2718 18226 2770
rect 18226 2718 18228 2770
rect 18172 2716 18228 2718
rect 25228 5068 25284 5124
rect 25228 4450 25284 4452
rect 25228 4398 25230 4450
rect 25230 4398 25282 4450
rect 25282 4398 25284 4450
rect 25228 4396 25284 4398
rect 18620 3442 18676 3444
rect 18620 3390 18622 3442
rect 18622 3390 18674 3442
rect 18674 3390 18676 3442
rect 18620 3388 18676 3390
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 19852 2994 19908 2996
rect 19852 2942 19854 2994
rect 19854 2942 19906 2994
rect 19906 2942 19908 2994
rect 19852 2940 19908 2942
rect 18172 1708 18228 1764
rect 19836 1594 19892 1596
rect 19836 1542 19838 1594
rect 19838 1542 19890 1594
rect 19890 1542 19892 1594
rect 19836 1540 19892 1542
rect 19940 1594 19996 1596
rect 19940 1542 19942 1594
rect 19942 1542 19994 1594
rect 19994 1542 19996 1594
rect 19940 1540 19996 1542
rect 20044 1594 20100 1596
rect 20044 1542 20046 1594
rect 20046 1542 20098 1594
rect 20098 1542 20100 1594
rect 20044 1540 20100 1542
rect 21420 2828 21476 2884
rect 22316 2882 22372 2884
rect 22316 2830 22318 2882
rect 22318 2830 22370 2882
rect 22370 2830 22372 2882
rect 22316 2828 22372 2830
rect 21980 1986 22036 1988
rect 21980 1934 21982 1986
rect 21982 1934 22034 1986
rect 22034 1934 22036 1986
rect 21980 1932 22036 1934
rect 25564 3276 25620 3332
rect 26572 5180 26628 5236
rect 27916 9996 27972 10052
rect 29148 9884 29204 9940
rect 29708 9660 29764 9716
rect 28700 8428 28756 8484
rect 29932 8482 29988 8484
rect 29932 8430 29934 8482
rect 29934 8430 29986 8482
rect 29986 8430 29988 8482
rect 29932 8428 29988 8430
rect 30716 16156 30772 16212
rect 30604 14924 30660 14980
rect 30604 14642 30660 14644
rect 30604 14590 30606 14642
rect 30606 14590 30658 14642
rect 30658 14590 30660 14642
rect 30604 14588 30660 14590
rect 30156 13132 30212 13188
rect 31052 18732 31108 18788
rect 31388 18338 31444 18340
rect 31388 18286 31390 18338
rect 31390 18286 31442 18338
rect 31442 18286 31444 18338
rect 31388 18284 31444 18286
rect 32060 18284 32116 18340
rect 32508 17724 32564 17780
rect 33292 17778 33348 17780
rect 33292 17726 33294 17778
rect 33294 17726 33346 17778
rect 33346 17726 33348 17778
rect 33292 17724 33348 17726
rect 33180 17612 33236 17668
rect 31052 16156 31108 16212
rect 32508 17106 32564 17108
rect 32508 17054 32510 17106
rect 32510 17054 32562 17106
rect 32562 17054 32564 17106
rect 32508 17052 32564 17054
rect 33180 17052 33236 17108
rect 34300 18732 34356 18788
rect 34636 18396 34692 18452
rect 34188 17778 34244 17780
rect 34188 17726 34190 17778
rect 34190 17726 34242 17778
rect 34242 17726 34244 17778
rect 34188 17724 34244 17726
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 34860 19404 34916 19460
rect 35196 19010 35252 19012
rect 35196 18958 35198 19010
rect 35198 18958 35250 19010
rect 35250 18958 35252 19010
rect 35196 18956 35252 18958
rect 34860 18732 34916 18788
rect 34972 18508 35028 18564
rect 36092 21420 36148 21476
rect 35756 19404 35812 19460
rect 36428 33292 36484 33348
rect 36428 30882 36484 30884
rect 36428 30830 36430 30882
rect 36430 30830 36482 30882
rect 36482 30830 36484 30882
rect 36428 30828 36484 30830
rect 36764 35586 36820 35588
rect 36764 35534 36766 35586
rect 36766 35534 36818 35586
rect 36818 35534 36820 35586
rect 36764 35532 36820 35534
rect 36876 42924 36932 42980
rect 36988 42642 37044 42644
rect 36988 42590 36990 42642
rect 36990 42590 37042 42642
rect 37042 42590 37044 42642
rect 36988 42588 37044 42590
rect 37436 41410 37492 41412
rect 37436 41358 37438 41410
rect 37438 41358 37490 41410
rect 37490 41358 37492 41410
rect 37436 41356 37492 41358
rect 37100 41298 37156 41300
rect 37100 41246 37102 41298
rect 37102 41246 37154 41298
rect 37154 41246 37156 41298
rect 37100 41244 37156 41246
rect 37996 46956 38052 47012
rect 38108 45612 38164 45668
rect 38220 42866 38276 42868
rect 38220 42814 38222 42866
rect 38222 42814 38274 42866
rect 38274 42814 38276 42866
rect 38220 42812 38276 42814
rect 36988 37938 37044 37940
rect 36988 37886 36990 37938
rect 36990 37886 37042 37938
rect 37042 37886 37044 37938
rect 36988 37884 37044 37886
rect 38220 41692 38276 41748
rect 37772 38050 37828 38052
rect 37772 37998 37774 38050
rect 37774 37998 37826 38050
rect 37826 37998 37828 38050
rect 37772 37996 37828 37998
rect 37548 37884 37604 37940
rect 36988 35756 37044 35812
rect 37212 35532 37268 35588
rect 36988 35308 37044 35364
rect 36876 34188 36932 34244
rect 37436 37154 37492 37156
rect 37436 37102 37438 37154
rect 37438 37102 37490 37154
rect 37490 37102 37492 37154
rect 37436 37100 37492 37102
rect 36876 33292 36932 33348
rect 38220 34300 38276 34356
rect 36988 33234 37044 33236
rect 36988 33182 36990 33234
rect 36990 33182 37042 33234
rect 37042 33182 37044 33234
rect 36988 33180 37044 33182
rect 36988 31666 37044 31668
rect 36988 31614 36990 31666
rect 36990 31614 37042 31666
rect 37042 31614 37044 31666
rect 36988 31612 37044 31614
rect 36988 27244 37044 27300
rect 36764 25340 36820 25396
rect 36540 23436 36596 23492
rect 36988 21474 37044 21476
rect 36988 21422 36990 21474
rect 36990 21422 37042 21474
rect 37042 21422 37044 21474
rect 36988 21420 37044 21422
rect 36316 20076 36372 20132
rect 36988 18956 37044 19012
rect 35756 18508 35812 18564
rect 35980 18396 36036 18452
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 35084 17666 35140 17668
rect 35084 17614 35086 17666
rect 35086 17614 35138 17666
rect 35138 17614 35140 17666
rect 35084 17612 35140 17614
rect 30940 15260 30996 15316
rect 31836 15260 31892 15316
rect 31164 14642 31220 14644
rect 31164 14590 31166 14642
rect 31166 14590 31218 14642
rect 31218 14590 31220 14642
rect 31164 14588 31220 14590
rect 34636 16044 34692 16100
rect 34636 15148 34692 15204
rect 36652 18284 36708 18340
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 35196 16098 35252 16100
rect 35196 16046 35198 16098
rect 35198 16046 35250 16098
rect 35250 16046 35252 16098
rect 35196 16044 35252 16046
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 31500 14306 31556 14308
rect 31500 14254 31502 14306
rect 31502 14254 31554 14306
rect 31554 14254 31556 14306
rect 31500 14252 31556 14254
rect 31500 13634 31556 13636
rect 31500 13582 31502 13634
rect 31502 13582 31554 13634
rect 31554 13582 31556 13634
rect 31500 13580 31556 13582
rect 33292 14252 33348 14308
rect 31948 13580 32004 13636
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 31164 13186 31220 13188
rect 31164 13134 31166 13186
rect 31166 13134 31218 13186
rect 31218 13134 31220 13186
rect 31164 13132 31220 13134
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 30268 11506 30324 11508
rect 30268 11454 30270 11506
rect 30270 11454 30322 11506
rect 30322 11454 30324 11506
rect 30268 11452 30324 11454
rect 31388 11228 31444 11284
rect 32396 11282 32452 11284
rect 32396 11230 32398 11282
rect 32398 11230 32450 11282
rect 32450 11230 32452 11282
rect 32396 11228 32452 11230
rect 31724 9938 31780 9940
rect 31724 9886 31726 9938
rect 31726 9886 31778 9938
rect 31778 9886 31780 9938
rect 31724 9884 31780 9886
rect 31500 9826 31556 9828
rect 31500 9774 31502 9826
rect 31502 9774 31554 9826
rect 31554 9774 31556 9826
rect 31500 9772 31556 9774
rect 30828 9714 30884 9716
rect 30828 9662 30830 9714
rect 30830 9662 30882 9714
rect 30882 9662 30884 9714
rect 30828 9660 30884 9662
rect 30156 8428 30212 8484
rect 30044 7644 30100 7700
rect 27692 7532 27748 7588
rect 30156 7362 30212 7364
rect 30156 7310 30158 7362
rect 30158 7310 30210 7362
rect 30210 7310 30212 7362
rect 30156 7308 30212 7310
rect 27356 6636 27412 6692
rect 32172 9826 32228 9828
rect 32172 9774 32174 9826
rect 32174 9774 32226 9826
rect 32226 9774 32228 9826
rect 32172 9772 32228 9774
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 38220 30828 38276 30884
rect 38220 27132 38276 27188
rect 37548 25394 37604 25396
rect 37548 25342 37550 25394
rect 37550 25342 37602 25394
rect 37602 25342 37604 25394
rect 37548 25340 37604 25342
rect 38220 25116 38276 25172
rect 37884 24892 37940 24948
rect 37772 21586 37828 21588
rect 37772 21534 37774 21586
rect 37774 21534 37826 21586
rect 37826 21534 37828 21586
rect 37772 21532 37828 21534
rect 37436 18338 37492 18340
rect 37436 18286 37438 18338
rect 37438 18286 37490 18338
rect 37490 18286 37492 18338
rect 37436 18284 37492 18286
rect 38108 17612 38164 17668
rect 37212 9660 37268 9716
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 38332 8540 38388 8596
rect 31948 8428 32004 8484
rect 31276 7980 31332 8036
rect 31388 7698 31444 7700
rect 31388 7646 31390 7698
rect 31390 7646 31442 7698
rect 31442 7646 31444 7698
rect 31388 7644 31444 7646
rect 31948 8034 32004 8036
rect 31948 7982 31950 8034
rect 31950 7982 32002 8034
rect 32002 7982 32004 8034
rect 31948 7980 32004 7982
rect 31500 7308 31556 7364
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35196 5514 35252 5516
rect 27356 5404 27412 5460
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 27692 5180 27748 5236
rect 23212 2716 23268 2772
rect 25228 2770 25284 2772
rect 25228 2718 25230 2770
rect 25230 2718 25282 2770
rect 25282 2718 25284 2770
rect 25228 2716 25284 2718
rect 23660 1986 23716 1988
rect 23660 1934 23662 1986
rect 23662 1934 23714 1986
rect 23714 1934 23716 1986
rect 23660 1932 23716 1934
rect 25788 2828 25844 2884
rect 26796 2882 26852 2884
rect 26796 2830 26798 2882
rect 26798 2830 26850 2882
rect 26850 2830 26852 2882
rect 26796 2828 26852 2830
rect 26572 2604 26628 2660
rect 27020 3330 27076 3332
rect 27020 3278 27022 3330
rect 27022 3278 27074 3330
rect 27074 3278 27076 3330
rect 27020 3276 27076 3278
rect 27356 2658 27412 2660
rect 27356 2606 27358 2658
rect 27358 2606 27410 2658
rect 27410 2606 27412 2658
rect 27356 2604 27412 2606
rect 27916 1708 27972 1764
rect 29148 1762 29204 1764
rect 29148 1710 29150 1762
rect 29150 1710 29202 1762
rect 29202 1710 29204 1762
rect 29148 1708 29204 1710
rect 32508 3388 32564 3444
rect 33628 3442 33684 3444
rect 33628 3390 33630 3442
rect 33630 3390 33682 3442
rect 33682 3390 33684 3442
rect 33628 3388 33684 3390
rect 33180 2546 33236 2548
rect 33180 2494 33182 2546
rect 33182 2494 33234 2546
rect 33234 2494 33236 2546
rect 33180 2492 33236 2494
rect 34412 2940 34468 2996
rect 33740 1986 33796 1988
rect 33740 1934 33742 1986
rect 33742 1934 33794 1986
rect 33794 1934 33796 1986
rect 33740 1932 33796 1934
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 34748 3052 34804 3108
rect 36652 3052 36708 3108
rect 35980 2940 36036 2996
rect 34860 2604 34916 2660
rect 35196 2378 35252 2380
rect 35196 2326 35198 2378
rect 35198 2326 35250 2378
rect 35250 2326 35252 2378
rect 35196 2324 35252 2326
rect 35300 2378 35356 2380
rect 35300 2326 35302 2378
rect 35302 2326 35354 2378
rect 35354 2326 35356 2378
rect 35300 2324 35356 2326
rect 35404 2378 35460 2380
rect 35404 2326 35406 2378
rect 35406 2326 35458 2378
rect 35458 2326 35460 2378
rect 35404 2324 35460 2326
rect 35308 1986 35364 1988
rect 35308 1934 35310 1986
rect 35310 1934 35362 1986
rect 35362 1934 35364 1986
rect 35308 1932 35364 1934
rect 35196 1820 35252 1876
rect 36092 2658 36148 2660
rect 36092 2606 36094 2658
rect 36094 2606 36146 2658
rect 36146 2606 36148 2658
rect 36092 2604 36148 2606
rect 36204 1820 36260 1876
rect 36092 1708 36148 1764
rect 36876 1708 36932 1764
rect 37436 1762 37492 1764
rect 37436 1710 37438 1762
rect 37438 1710 37490 1762
rect 37490 1710 37492 1762
rect 37436 1708 37492 1710
<< metal3 >>
rect 4466 97972 4476 98028
rect 4532 97972 4580 98028
rect 4636 97972 4684 98028
rect 4740 97972 4750 98028
rect 35186 97972 35196 98028
rect 35252 97972 35300 98028
rect 35356 97972 35404 98028
rect 35460 97972 35470 98028
rect 13010 97468 13020 97524
rect 13076 97468 14476 97524
rect 14532 97468 14542 97524
rect 13682 97356 13692 97412
rect 13748 97356 15708 97412
rect 15764 97356 15774 97412
rect 16146 97356 16156 97412
rect 16212 97356 16940 97412
rect 16996 97356 17006 97412
rect 26786 97356 26796 97412
rect 26852 97356 28476 97412
rect 28532 97356 28542 97412
rect 19826 97188 19836 97244
rect 19892 97188 19940 97244
rect 19996 97188 20044 97244
rect 20100 97188 20110 97244
rect 32274 96796 32284 96852
rect 32340 96796 32956 96852
rect 33012 96796 35196 96852
rect 35252 96796 35262 96852
rect 6178 96572 6188 96628
rect 6244 96572 6860 96628
rect 6916 96572 7644 96628
rect 7700 96572 7710 96628
rect 4466 96404 4476 96460
rect 4532 96404 4580 96460
rect 4636 96404 4684 96460
rect 4740 96404 4750 96460
rect 35186 96404 35196 96460
rect 35252 96404 35300 96460
rect 35356 96404 35404 96460
rect 35460 96404 35470 96460
rect 25330 96124 25340 96180
rect 25396 96124 35868 96180
rect 35924 96124 35934 96180
rect 6738 96012 6748 96068
rect 6804 96012 8876 96068
rect 8932 96012 9324 96068
rect 9380 96012 9390 96068
rect 30146 96012 30156 96068
rect 30212 96012 31276 96068
rect 31332 96012 31342 96068
rect 24210 95900 24220 95956
rect 24276 95900 33404 95956
rect 33460 95900 33470 95956
rect 8642 95788 8652 95844
rect 8708 95788 9660 95844
rect 9716 95788 10332 95844
rect 10388 95788 11676 95844
rect 11732 95788 11742 95844
rect 21410 95788 21420 95844
rect 21476 95788 22092 95844
rect 22148 95788 22158 95844
rect 26450 95788 26460 95844
rect 26516 95788 27356 95844
rect 27412 95788 27422 95844
rect 33170 95788 33180 95844
rect 33236 95788 35196 95844
rect 35252 95788 35262 95844
rect 13570 95676 13580 95732
rect 13636 95676 14700 95732
rect 14756 95676 14766 95732
rect 16258 95676 16268 95732
rect 16324 95676 19516 95732
rect 19572 95676 19582 95732
rect 26002 95676 26012 95732
rect 26068 95676 30940 95732
rect 30996 95676 31006 95732
rect 19826 95620 19836 95676
rect 19892 95620 19940 95676
rect 19996 95620 20044 95676
rect 20100 95620 20110 95676
rect 12338 95452 12348 95508
rect 12404 95452 13916 95508
rect 13972 95452 14476 95508
rect 14532 95452 15148 95508
rect 15204 95452 15214 95508
rect 23538 95452 23548 95508
rect 23604 95452 25116 95508
rect 25172 95452 25182 95508
rect 16818 95340 16828 95396
rect 16884 95340 17500 95396
rect 17556 95340 17566 95396
rect 20626 95228 20636 95284
rect 20692 95228 21196 95284
rect 21252 95228 22316 95284
rect 22372 95228 23324 95284
rect 23380 95228 24668 95284
rect 24724 95228 26012 95284
rect 26068 95228 26078 95284
rect 27794 95228 27804 95284
rect 27860 95228 29148 95284
rect 29204 95228 29596 95284
rect 29652 95228 30156 95284
rect 30212 95228 30222 95284
rect 33058 95228 33068 95284
rect 33124 95228 35644 95284
rect 35700 95228 35710 95284
rect 34066 95116 34076 95172
rect 34132 95116 36428 95172
rect 36484 95116 36494 95172
rect 35186 95004 35196 95060
rect 35252 95004 37772 95060
rect 37828 95004 37838 95060
rect 4466 94836 4476 94892
rect 4532 94836 4580 94892
rect 4636 94836 4684 94892
rect 4740 94836 4750 94892
rect 35186 94836 35196 94892
rect 35252 94836 35300 94892
rect 35356 94836 35404 94892
rect 35460 94836 35470 94892
rect 14690 94668 14700 94724
rect 14756 94668 15596 94724
rect 15652 94668 15662 94724
rect 26226 94556 26236 94612
rect 26292 94556 27356 94612
rect 27412 94556 27422 94612
rect 17490 94444 17500 94500
rect 17556 94444 18508 94500
rect 18564 94444 18574 94500
rect 0 94388 400 94416
rect 0 94332 1708 94388
rect 1764 94332 1774 94388
rect 20290 94332 20300 94388
rect 20356 94332 21980 94388
rect 22036 94332 22046 94388
rect 0 94304 400 94332
rect 19826 94052 19836 94108
rect 19892 94052 19940 94108
rect 19996 94052 20044 94108
rect 20100 94052 20110 94108
rect 17266 93996 17276 94052
rect 17332 93996 17724 94052
rect 17780 93996 17790 94052
rect 31826 93996 31836 94052
rect 31892 93996 32844 94052
rect 32900 93996 32910 94052
rect 20626 93884 20636 93940
rect 20692 93884 21532 93940
rect 21588 93884 21598 93940
rect 27458 93884 27468 93940
rect 27524 93884 30492 93940
rect 30548 93884 30558 93940
rect 2930 93660 2940 93716
rect 2996 93660 4172 93716
rect 4228 93660 6748 93716
rect 6804 93660 6814 93716
rect 10322 93660 10332 93716
rect 10388 93660 12012 93716
rect 12068 93660 12078 93716
rect 13346 93660 13356 93716
rect 13412 93660 14140 93716
rect 14196 93660 14206 93716
rect 15922 93660 15932 93716
rect 15988 93660 16604 93716
rect 16660 93660 17052 93716
rect 17108 93660 17118 93716
rect 18386 93660 18396 93716
rect 18452 93660 19292 93716
rect 19348 93660 19358 93716
rect 12674 93548 12684 93604
rect 12740 93548 14588 93604
rect 14644 93548 14654 93604
rect 2034 93436 2044 93492
rect 2100 93436 3388 93492
rect 3444 93436 3454 93492
rect 24406 93436 24444 93492
rect 24500 93436 24510 93492
rect 17714 93324 17724 93380
rect 17780 93324 20076 93380
rect 20132 93324 20748 93380
rect 20804 93324 23212 93380
rect 23268 93324 24668 93380
rect 24724 93324 24734 93380
rect 4466 93268 4476 93324
rect 4532 93268 4580 93324
rect 4636 93268 4684 93324
rect 4740 93268 4750 93324
rect 35186 93268 35196 93324
rect 35252 93268 35300 93324
rect 35356 93268 35404 93324
rect 35460 93268 35470 93324
rect 30930 93100 30940 93156
rect 30996 93100 31500 93156
rect 31556 93100 31948 93156
rect 31892 93044 31948 93100
rect 14242 92988 14252 93044
rect 14308 92988 17276 93044
rect 17332 92988 18620 93044
rect 18676 92988 20972 93044
rect 21028 92988 21038 93044
rect 31892 92988 32508 93044
rect 32564 92988 32574 93044
rect 30146 92876 30156 92932
rect 30212 92876 32732 92932
rect 32788 92876 33852 92932
rect 33908 92876 33918 92932
rect 9650 92764 9660 92820
rect 9716 92764 10780 92820
rect 10836 92764 10846 92820
rect 12562 92764 12572 92820
rect 12628 92764 13804 92820
rect 13860 92764 13870 92820
rect 26226 92764 26236 92820
rect 26292 92764 26684 92820
rect 26740 92764 26750 92820
rect 27458 92764 27468 92820
rect 27524 92764 29260 92820
rect 29316 92764 31836 92820
rect 31892 92764 33180 92820
rect 33236 92764 33246 92820
rect 17938 92652 17948 92708
rect 18004 92652 19404 92708
rect 19460 92652 22204 92708
rect 22260 92652 22270 92708
rect 25218 92652 25228 92708
rect 25284 92652 26124 92708
rect 26180 92652 26190 92708
rect 32498 92652 32508 92708
rect 32564 92652 34076 92708
rect 34132 92652 35084 92708
rect 35140 92652 35150 92708
rect 6514 92540 6524 92596
rect 6580 92540 6972 92596
rect 7028 92540 10780 92596
rect 10836 92540 10846 92596
rect 19826 92484 19836 92540
rect 19892 92484 19940 92540
rect 19996 92484 20044 92540
rect 20100 92484 20110 92540
rect 7298 92428 7308 92484
rect 7364 92428 7756 92484
rect 7812 92428 9660 92484
rect 9716 92428 9726 92484
rect 23874 92428 23884 92484
rect 23940 92428 25564 92484
rect 25620 92428 26460 92484
rect 26516 92428 26526 92484
rect 13570 92316 13580 92372
rect 13636 92316 14364 92372
rect 14420 92316 14430 92372
rect 10210 92204 10220 92260
rect 10276 92204 12908 92260
rect 12964 92204 14700 92260
rect 14756 92204 15148 92260
rect 15204 92204 16828 92260
rect 16884 92204 16894 92260
rect 26114 92204 26124 92260
rect 26180 92204 26908 92260
rect 26852 92148 26908 92204
rect 3826 92092 3836 92148
rect 3892 92092 4956 92148
rect 5012 92092 5022 92148
rect 12338 92092 12348 92148
rect 12404 92092 25340 92148
rect 25396 92092 25676 92148
rect 25732 92092 25742 92148
rect 26852 92092 27356 92148
rect 27412 92092 27422 92148
rect 21634 91980 21644 92036
rect 21700 91980 23324 92036
rect 23380 91980 23390 92036
rect 26852 91980 28364 92036
rect 28420 91980 28430 92036
rect 37650 91980 37660 92036
rect 37716 91980 38220 92036
rect 38276 91980 38286 92036
rect 26852 91924 26908 91980
rect 20962 91868 20972 91924
rect 21028 91868 22428 91924
rect 22484 91868 23996 91924
rect 24052 91868 24668 91924
rect 24724 91868 26124 91924
rect 26180 91868 26908 91924
rect 4466 91700 4476 91756
rect 4532 91700 4580 91756
rect 4636 91700 4684 91756
rect 4740 91700 4750 91756
rect 35186 91700 35196 91756
rect 35252 91700 35300 91756
rect 35356 91700 35404 91756
rect 35460 91700 35470 91756
rect 39600 91476 40000 91504
rect 38210 91420 38220 91476
rect 38276 91420 40000 91476
rect 39600 91392 40000 91420
rect 11554 91308 11564 91364
rect 11620 91308 12012 91364
rect 12068 91308 13580 91364
rect 13636 91308 13646 91364
rect 33170 91308 33180 91364
rect 33236 91308 34524 91364
rect 34580 91308 34590 91364
rect 19826 90916 19836 90972
rect 19892 90916 19940 90972
rect 19996 90916 20044 90972
rect 20100 90916 20110 90972
rect 11666 90636 11676 90692
rect 11732 90636 12348 90692
rect 12404 90636 12414 90692
rect 24098 90636 24108 90692
rect 24164 90636 24556 90692
rect 24612 90636 29708 90692
rect 29764 90636 30156 90692
rect 30212 90636 35084 90692
rect 35140 90636 35150 90692
rect 22978 90524 22988 90580
rect 23044 90524 25116 90580
rect 25172 90524 25508 90580
rect 25452 90468 25508 90524
rect 21858 90412 21868 90468
rect 21924 90412 23548 90468
rect 23604 90412 23614 90468
rect 25442 90412 25452 90468
rect 25508 90412 28252 90468
rect 28308 90412 28318 90468
rect 4466 90132 4476 90188
rect 4532 90132 4580 90188
rect 4636 90132 4684 90188
rect 4740 90132 4750 90188
rect 35186 90132 35196 90188
rect 35252 90132 35300 90188
rect 35356 90132 35404 90188
rect 35460 90132 35470 90188
rect 21634 89852 21644 89908
rect 21700 89852 21980 89908
rect 22036 89852 23436 89908
rect 23492 89852 23502 89908
rect 3154 89740 3164 89796
rect 3220 89740 4284 89796
rect 4340 89740 4350 89796
rect 19954 89740 19964 89796
rect 20020 89740 24556 89796
rect 24612 89740 24622 89796
rect 22082 89628 22092 89684
rect 22148 89628 22876 89684
rect 22932 89628 22942 89684
rect 17490 89516 17500 89572
rect 17556 89516 19516 89572
rect 19572 89516 19582 89572
rect 21746 89516 21756 89572
rect 21812 89516 23324 89572
rect 23380 89516 23390 89572
rect 26114 89516 26124 89572
rect 26180 89516 27468 89572
rect 27524 89516 27534 89572
rect 21858 89404 21868 89460
rect 21924 89404 22540 89460
rect 22596 89404 23212 89460
rect 23268 89404 24444 89460
rect 24500 89404 26236 89460
rect 26292 89404 26908 89460
rect 19826 89348 19836 89404
rect 19892 89348 19940 89404
rect 19996 89348 20044 89404
rect 20100 89348 20110 89404
rect 23538 89292 23548 89348
rect 23604 89292 24108 89348
rect 24164 89292 24174 89348
rect 22866 89180 22876 89236
rect 22932 89180 23660 89236
rect 23716 89180 24892 89236
rect 24948 89180 24958 89236
rect 14242 89068 14252 89124
rect 14308 89068 15932 89124
rect 15988 89068 16716 89124
rect 16772 89068 19628 89124
rect 19684 89068 19694 89124
rect 22082 89068 22092 89124
rect 22148 89068 24220 89124
rect 24276 89068 24286 89124
rect 24770 89068 24780 89124
rect 24836 89068 25228 89124
rect 25284 89068 25294 89124
rect 26852 89068 26908 89404
rect 26964 89068 28028 89124
rect 28084 89068 29260 89124
rect 29316 89068 29326 89124
rect 6850 88956 6860 89012
rect 6916 88956 7980 89012
rect 8036 88956 8046 89012
rect 13346 88956 13356 89012
rect 13412 88956 16044 89012
rect 16100 88956 16110 89012
rect 21186 88956 21196 89012
rect 21252 88956 22204 89012
rect 22260 88956 23436 89012
rect 23492 88956 23502 89012
rect 24434 88956 24444 89012
rect 24500 88956 27468 89012
rect 27524 88956 27534 89012
rect 18274 88844 18284 88900
rect 18340 88844 19516 88900
rect 19572 88844 19582 88900
rect 22978 88844 22988 88900
rect 23044 88844 23996 88900
rect 24052 88844 25788 88900
rect 25844 88844 25854 88900
rect 27682 88844 27692 88900
rect 27748 88844 30156 88900
rect 30212 88844 30222 88900
rect 19170 88732 19180 88788
rect 19236 88732 25116 88788
rect 25172 88732 25900 88788
rect 25956 88732 25966 88788
rect 19058 88620 19068 88676
rect 19124 88620 27356 88676
rect 27412 88620 27422 88676
rect 4466 88564 4476 88620
rect 4532 88564 4580 88620
rect 4636 88564 4684 88620
rect 4740 88564 4750 88620
rect 35186 88564 35196 88620
rect 35252 88564 35300 88620
rect 35356 88564 35404 88620
rect 35460 88564 35470 88620
rect 23874 88508 23884 88564
rect 23940 88508 23950 88564
rect 20626 88396 20636 88452
rect 20692 88396 22764 88452
rect 22820 88396 22830 88452
rect 23884 88340 23940 88508
rect 16706 88284 16716 88340
rect 16772 88284 16940 88340
rect 16996 88284 17006 88340
rect 23874 88284 23884 88340
rect 23940 88284 23950 88340
rect 7970 88172 7980 88228
rect 8036 88172 9660 88228
rect 9716 88172 9726 88228
rect 21522 88172 21532 88228
rect 21588 88172 22204 88228
rect 22260 88172 22428 88228
rect 22484 88172 22494 88228
rect 28578 88172 28588 88228
rect 28644 88172 29260 88228
rect 29316 88172 31052 88228
rect 31108 88172 32508 88228
rect 32564 88172 32574 88228
rect 8372 88060 9324 88116
rect 9380 88060 10556 88116
rect 10612 88060 10622 88116
rect 24098 88060 24108 88116
rect 24164 88060 27804 88116
rect 27860 88060 27870 88116
rect 8372 88004 8428 88060
rect 7746 87948 7756 88004
rect 7812 87948 8428 88004
rect 8484 87948 8494 88004
rect 10658 87948 10668 88004
rect 10724 87948 12236 88004
rect 12292 87948 12302 88004
rect 13794 87948 13804 88004
rect 13860 87948 14252 88004
rect 14308 87948 14318 88004
rect 19730 87948 19740 88004
rect 19796 87948 20188 88004
rect 20244 87948 21196 88004
rect 21252 87948 21262 88004
rect 24770 87948 24780 88004
rect 24836 87948 25564 88004
rect 25620 87948 27020 88004
rect 27076 87948 29148 88004
rect 29204 87948 29214 88004
rect 35074 87948 35084 88004
rect 35140 87948 35532 88004
rect 35588 87948 36204 88004
rect 36260 87948 36270 88004
rect 9538 87836 9548 87892
rect 9604 87836 12012 87892
rect 12068 87836 12078 87892
rect 24546 87836 24556 87892
rect 24612 87836 25004 87892
rect 25060 87836 25070 87892
rect 27346 87836 27356 87892
rect 27412 87836 29484 87892
rect 29540 87836 29550 87892
rect 19826 87780 19836 87836
rect 19892 87780 19940 87836
rect 19996 87780 20044 87836
rect 20100 87780 20110 87836
rect 12450 87724 12460 87780
rect 12516 87724 14140 87780
rect 14196 87724 14206 87780
rect 20402 87724 20412 87780
rect 20468 87724 22764 87780
rect 22820 87724 22830 87780
rect 15250 87612 15260 87668
rect 15316 87612 15708 87668
rect 15764 87612 16044 87668
rect 16100 87612 16716 87668
rect 16772 87612 17500 87668
rect 17556 87612 18732 87668
rect 18788 87612 20076 87668
rect 20132 87612 21196 87668
rect 21252 87612 21262 87668
rect 23762 87612 23772 87668
rect 23828 87612 25452 87668
rect 25508 87612 26236 87668
rect 26292 87612 26302 87668
rect 31892 87612 32060 87668
rect 32116 87612 32126 87668
rect 10546 87500 10556 87556
rect 10612 87500 13580 87556
rect 13636 87500 13646 87556
rect 15092 87500 21084 87556
rect 21140 87500 21252 87556
rect 24518 87500 24556 87556
rect 24612 87500 24622 87556
rect 25330 87500 25340 87556
rect 25396 87500 27244 87556
rect 27300 87500 27310 87556
rect 15092 87444 15148 87500
rect 13010 87388 13020 87444
rect 13076 87388 13916 87444
rect 13972 87388 15148 87444
rect 15586 87388 15596 87444
rect 15652 87388 17836 87444
rect 17892 87388 17902 87444
rect 19618 87388 19628 87444
rect 19684 87388 20972 87444
rect 21028 87388 21038 87444
rect 21196 87220 21252 87500
rect 31892 87444 31948 87612
rect 24658 87388 24668 87444
rect 24724 87388 26572 87444
rect 26628 87388 26638 87444
rect 30370 87388 30380 87444
rect 30436 87388 31052 87444
rect 31108 87388 31948 87444
rect 32050 87388 32060 87444
rect 32116 87388 32956 87444
rect 33012 87388 33022 87444
rect 33506 87276 33516 87332
rect 33572 87276 34972 87332
rect 35028 87276 35038 87332
rect 6962 87164 6972 87220
rect 7028 87164 9100 87220
rect 9156 87164 9166 87220
rect 21196 87164 27132 87220
rect 27188 87164 27198 87220
rect 4466 86996 4476 87052
rect 4532 86996 4580 87052
rect 4636 86996 4684 87052
rect 4740 86996 4750 87052
rect 35186 86996 35196 87052
rect 35252 86996 35300 87052
rect 35356 86996 35404 87052
rect 35460 86996 35470 87052
rect 25106 86940 25116 86996
rect 25172 86940 28028 86996
rect 28084 86940 28094 86996
rect 20738 86828 20748 86884
rect 20804 86828 22652 86884
rect 22708 86828 22718 86884
rect 24434 86828 24444 86884
rect 24500 86828 24668 86884
rect 24724 86828 24734 86884
rect 15092 86716 20636 86772
rect 20692 86716 21980 86772
rect 22036 86716 22046 86772
rect 22194 86716 22204 86772
rect 22260 86716 22876 86772
rect 22932 86716 25116 86772
rect 25172 86716 25182 86772
rect 29586 86716 29596 86772
rect 29652 86716 30828 86772
rect 30884 86716 30894 86772
rect 9314 86604 9324 86660
rect 9380 86604 10108 86660
rect 10164 86604 10174 86660
rect 15092 86548 15148 86716
rect 15810 86604 15820 86660
rect 15876 86604 16940 86660
rect 16996 86604 17006 86660
rect 20738 86604 20748 86660
rect 20804 86604 23660 86660
rect 23716 86604 23726 86660
rect 24882 86604 24892 86660
rect 24948 86604 26012 86660
rect 26068 86604 26124 86660
rect 26180 86604 26190 86660
rect 4274 86492 4284 86548
rect 4340 86492 10892 86548
rect 10948 86492 10958 86548
rect 14130 86492 14140 86548
rect 14196 86492 15148 86548
rect 26898 86492 26908 86548
rect 26964 86492 27692 86548
rect 27748 86492 27758 86548
rect 21074 86380 21084 86436
rect 21140 86380 23660 86436
rect 23716 86380 24108 86436
rect 24164 86380 24174 86436
rect 24658 86380 24668 86436
rect 24724 86380 27916 86436
rect 27972 86380 27982 86436
rect 19826 86212 19836 86268
rect 19892 86212 19940 86268
rect 19996 86212 20044 86268
rect 20100 86212 20110 86268
rect 21746 86156 21756 86212
rect 21812 86156 24332 86212
rect 24388 86156 24398 86212
rect 11554 86044 11564 86100
rect 11620 86044 12124 86100
rect 12180 86044 12796 86100
rect 12852 86044 12862 86100
rect 23538 86044 23548 86100
rect 23604 86044 24892 86100
rect 24948 86044 24958 86100
rect 32834 86044 32844 86100
rect 32900 86044 33628 86100
rect 33684 86044 33694 86100
rect 5394 85820 5404 85876
rect 5460 85820 6972 85876
rect 7028 85820 7038 85876
rect 20738 85820 20748 85876
rect 20804 85820 25228 85876
rect 25284 85820 25294 85876
rect 29922 85820 29932 85876
rect 29988 85820 31164 85876
rect 31220 85820 31230 85876
rect 21970 85708 21980 85764
rect 22036 85708 28924 85764
rect 28980 85708 28990 85764
rect 30706 85708 30716 85764
rect 30772 85708 31836 85764
rect 31892 85708 31902 85764
rect 32498 85708 32508 85764
rect 32564 85708 33684 85764
rect 25890 85596 25900 85652
rect 25956 85596 27356 85652
rect 27412 85596 28476 85652
rect 28532 85596 28542 85652
rect 33628 85540 33684 85708
rect 33628 85484 33852 85540
rect 33908 85484 34524 85540
rect 34580 85484 34590 85540
rect 4466 85428 4476 85484
rect 4532 85428 4580 85484
rect 4636 85428 4684 85484
rect 4740 85428 4750 85484
rect 35186 85428 35196 85484
rect 35252 85428 35300 85484
rect 35356 85428 35404 85484
rect 35460 85428 35470 85484
rect 14018 85260 14028 85316
rect 14084 85260 15148 85316
rect 15204 85260 15214 85316
rect 31938 85260 31948 85316
rect 32004 85260 32508 85316
rect 32564 85260 33292 85316
rect 33348 85260 33358 85316
rect 18834 85148 18844 85204
rect 18900 85148 26908 85204
rect 29138 85148 29148 85204
rect 29204 85148 30828 85204
rect 30884 85148 30894 85204
rect 34738 85148 34748 85204
rect 34804 85148 35980 85204
rect 36036 85148 36876 85204
rect 36932 85148 36942 85204
rect 26852 85092 26908 85148
rect 13682 85036 13692 85092
rect 13748 85036 14588 85092
rect 14644 85036 15596 85092
rect 15652 85036 15662 85092
rect 19170 85036 19180 85092
rect 19236 85036 20188 85092
rect 20244 85036 21420 85092
rect 21476 85036 21486 85092
rect 26852 85036 31276 85092
rect 31332 85036 32060 85092
rect 32116 85036 32126 85092
rect 33618 85036 33628 85092
rect 33684 85036 34412 85092
rect 34468 85036 35084 85092
rect 35140 85036 35868 85092
rect 35924 85036 35934 85092
rect 27458 84924 27468 84980
rect 27524 84924 38332 84980
rect 38388 84924 38398 84980
rect 12898 84812 12908 84868
rect 12964 84812 13804 84868
rect 13860 84812 13870 84868
rect 18722 84812 18732 84868
rect 18788 84812 20076 84868
rect 20132 84812 20142 84868
rect 31490 84812 31500 84868
rect 31556 84812 32732 84868
rect 32788 84812 32798 84868
rect 34962 84812 34972 84868
rect 35028 84812 37660 84868
rect 37716 84812 37726 84868
rect 26226 84700 26236 84756
rect 26292 84700 30156 84756
rect 30212 84700 33964 84756
rect 34020 84700 35420 84756
rect 35476 84700 35486 84756
rect 19826 84644 19836 84700
rect 19892 84644 19940 84700
rect 19996 84644 20044 84700
rect 20100 84644 20110 84700
rect 20402 84588 20412 84644
rect 20468 84588 24220 84644
rect 24276 84588 29372 84644
rect 29428 84588 29438 84644
rect 30594 84588 30604 84644
rect 30660 84588 31052 84644
rect 31108 84588 36540 84644
rect 36596 84588 36606 84644
rect 0 84532 400 84560
rect 30604 84532 30660 84588
rect 0 84476 4956 84532
rect 5012 84476 5022 84532
rect 13906 84476 13916 84532
rect 13972 84476 17612 84532
rect 17668 84476 18844 84532
rect 18900 84476 18910 84532
rect 22306 84476 22316 84532
rect 22372 84476 23884 84532
rect 23940 84476 23950 84532
rect 25666 84476 25676 84532
rect 25732 84476 26236 84532
rect 26292 84476 26302 84532
rect 27346 84476 27356 84532
rect 27412 84476 28028 84532
rect 28084 84476 30660 84532
rect 34738 84476 34748 84532
rect 34804 84476 35308 84532
rect 35364 84476 35374 84532
rect 36418 84476 36428 84532
rect 36484 84476 37100 84532
rect 37156 84476 37166 84532
rect 0 84448 400 84476
rect 19954 84364 19964 84420
rect 20020 84364 23324 84420
rect 23380 84364 23390 84420
rect 28466 84364 28476 84420
rect 28532 84364 29708 84420
rect 29764 84364 29774 84420
rect 18834 84252 18844 84308
rect 18900 84252 20636 84308
rect 20692 84252 20702 84308
rect 24434 84252 24444 84308
rect 24500 84252 26908 84308
rect 26964 84252 27356 84308
rect 27412 84252 27422 84308
rect 12562 84140 12572 84196
rect 12628 84140 13692 84196
rect 13748 84140 13758 84196
rect 24210 84140 24220 84196
rect 24276 84140 25116 84196
rect 25172 84140 25788 84196
rect 25844 84140 25854 84196
rect 26012 84140 26908 84196
rect 27346 84140 27356 84196
rect 27412 84140 27468 84196
rect 27524 84140 27534 84196
rect 26012 84084 26068 84140
rect 16146 84028 16156 84084
rect 16212 84028 19740 84084
rect 19796 84028 22316 84084
rect 22372 84028 26068 84084
rect 26852 84084 26908 84140
rect 26852 84028 28476 84084
rect 28532 84028 28542 84084
rect 31938 84028 31948 84084
rect 32004 84028 34524 84084
rect 34580 84028 35700 84084
rect 37202 84028 37212 84084
rect 37268 84028 38108 84084
rect 38164 84028 38174 84084
rect 35644 83972 35700 84028
rect 35634 83916 35644 83972
rect 35700 83916 37660 83972
rect 37716 83916 38220 83972
rect 38276 83916 38286 83972
rect 4466 83860 4476 83916
rect 4532 83860 4580 83916
rect 4636 83860 4684 83916
rect 4740 83860 4750 83916
rect 35186 83860 35196 83916
rect 35252 83860 35300 83916
rect 35356 83860 35404 83916
rect 35460 83860 35470 83916
rect 17714 83692 17724 83748
rect 17780 83692 19180 83748
rect 19236 83692 19246 83748
rect 20066 83692 20076 83748
rect 20132 83692 20412 83748
rect 20468 83692 20478 83748
rect 27794 83692 27804 83748
rect 27860 83692 29260 83748
rect 29316 83692 29326 83748
rect 36082 83692 36092 83748
rect 36148 83692 37100 83748
rect 37156 83692 37166 83748
rect 19282 83580 19292 83636
rect 19348 83580 19964 83636
rect 20020 83580 20030 83636
rect 28354 83580 28364 83636
rect 28420 83580 30492 83636
rect 30548 83580 30558 83636
rect 18498 83468 18508 83524
rect 18564 83468 19516 83524
rect 19572 83468 21868 83524
rect 21924 83468 21934 83524
rect 34850 83468 34860 83524
rect 34916 83468 35980 83524
rect 36036 83468 36046 83524
rect 3266 83356 3276 83412
rect 3332 83356 4396 83412
rect 4452 83356 4462 83412
rect 13794 83356 13804 83412
rect 13860 83356 15596 83412
rect 15652 83356 17836 83412
rect 17892 83356 17902 83412
rect 18050 83356 18060 83412
rect 18116 83356 19292 83412
rect 19348 83356 20300 83412
rect 20356 83356 29596 83412
rect 29652 83356 31388 83412
rect 31444 83356 31454 83412
rect 36194 83356 36204 83412
rect 36260 83356 36988 83412
rect 37044 83356 37054 83412
rect 18284 83300 18340 83356
rect 12674 83244 12684 83300
rect 12740 83244 15260 83300
rect 15316 83244 15326 83300
rect 16594 83244 16604 83300
rect 16660 83244 17164 83300
rect 17220 83244 18284 83300
rect 18340 83244 18350 83300
rect 20402 83244 20412 83300
rect 20468 83244 22092 83300
rect 22148 83244 26012 83300
rect 26068 83244 26236 83300
rect 26292 83244 28364 83300
rect 28420 83244 30044 83300
rect 30100 83244 30940 83300
rect 30996 83244 31006 83300
rect 34626 83244 34636 83300
rect 34692 83244 37548 83300
rect 37604 83244 37614 83300
rect 16604 83188 16660 83244
rect 15362 83132 15372 83188
rect 15428 83132 16660 83188
rect 25890 83132 25900 83188
rect 25956 83132 30604 83188
rect 30660 83132 30670 83188
rect 19826 83076 19836 83132
rect 19892 83076 19940 83132
rect 19996 83076 20044 83132
rect 20100 83076 20110 83132
rect 14802 83020 14812 83076
rect 14868 83020 16156 83076
rect 16212 83020 16222 83076
rect 21410 83020 21420 83076
rect 21476 83020 22876 83076
rect 22932 83020 30156 83076
rect 30212 83020 30222 83076
rect 8418 82908 8428 82964
rect 8484 82908 9660 82964
rect 9716 82908 9726 82964
rect 14130 82908 14140 82964
rect 14196 82908 25900 82964
rect 25956 82908 25966 82964
rect 27122 82908 27132 82964
rect 27188 82908 29036 82964
rect 29092 82908 29102 82964
rect 10210 82796 10220 82852
rect 10276 82796 20524 82852
rect 20580 82796 20590 82852
rect 26450 82796 26460 82852
rect 26516 82796 29148 82852
rect 29204 82796 29214 82852
rect 22306 82684 22316 82740
rect 22372 82684 22988 82740
rect 23044 82684 25228 82740
rect 25284 82684 25294 82740
rect 26562 82684 26572 82740
rect 26628 82684 29372 82740
rect 29428 82684 29438 82740
rect 4946 82572 4956 82628
rect 5012 82572 6076 82628
rect 6132 82572 9772 82628
rect 9828 82572 9838 82628
rect 19394 82572 19404 82628
rect 19460 82572 20972 82628
rect 21028 82572 21038 82628
rect 27010 82572 27020 82628
rect 27076 82572 27356 82628
rect 27412 82572 28924 82628
rect 28980 82572 28990 82628
rect 31602 82572 31612 82628
rect 31668 82572 33180 82628
rect 33236 82572 34524 82628
rect 34580 82572 34590 82628
rect 7186 82460 7196 82516
rect 7252 82460 7980 82516
rect 8036 82460 8764 82516
rect 8820 82460 10668 82516
rect 10724 82460 11004 82516
rect 11060 82460 11070 82516
rect 14018 82460 14028 82516
rect 14084 82460 15148 82516
rect 15204 82460 15214 82516
rect 16930 82460 16940 82516
rect 16996 82460 18172 82516
rect 18228 82460 18396 82516
rect 18452 82460 20412 82516
rect 20468 82460 21084 82516
rect 21140 82460 21150 82516
rect 25442 82460 25452 82516
rect 25508 82460 26908 82516
rect 26964 82460 26974 82516
rect 27122 82460 27132 82516
rect 27188 82460 28028 82516
rect 28084 82460 28094 82516
rect 10434 82348 10444 82404
rect 10500 82348 11564 82404
rect 11620 82348 11630 82404
rect 12002 82348 12012 82404
rect 12068 82348 15148 82404
rect 24098 82348 24108 82404
rect 24164 82348 25788 82404
rect 25844 82348 25854 82404
rect 27206 82348 27244 82404
rect 27300 82348 27310 82404
rect 29810 82348 29820 82404
rect 29876 82348 33852 82404
rect 33908 82348 34636 82404
rect 34692 82348 34702 82404
rect 4466 82292 4476 82348
rect 4532 82292 4580 82348
rect 4636 82292 4684 82348
rect 4740 82292 4750 82348
rect 15092 82292 15148 82348
rect 35186 82292 35196 82348
rect 35252 82292 35300 82348
rect 35356 82292 35404 82348
rect 35460 82292 35470 82348
rect 15092 82236 15484 82292
rect 15540 82236 16380 82292
rect 16436 82236 16446 82292
rect 25890 82236 25900 82292
rect 25956 82236 27692 82292
rect 27748 82236 30380 82292
rect 30436 82236 30446 82292
rect 23650 82124 23660 82180
rect 23716 82124 24108 82180
rect 24164 82124 24174 82180
rect 26674 82124 26684 82180
rect 26740 82124 27356 82180
rect 27412 82124 28812 82180
rect 28868 82124 28878 82180
rect 24882 82012 24892 82068
rect 24948 82012 27804 82068
rect 27860 82012 27870 82068
rect 6626 81900 6636 81956
rect 6692 81900 21196 81956
rect 21252 81900 21262 81956
rect 24994 81900 25004 81956
rect 25060 81900 26348 81956
rect 26404 81900 26414 81956
rect 32946 81900 32956 81956
rect 33012 81900 34188 81956
rect 34244 81900 35196 81956
rect 35252 81900 36204 81956
rect 36260 81900 37884 81956
rect 37940 81900 37950 81956
rect 9650 81788 9660 81844
rect 9716 81788 10892 81844
rect 10948 81788 10958 81844
rect 25442 81788 25452 81844
rect 25508 81788 26908 81844
rect 26964 81788 28588 81844
rect 28644 81788 28654 81844
rect 5842 81676 5852 81732
rect 5908 81676 7196 81732
rect 7252 81676 7262 81732
rect 23090 81676 23100 81732
rect 23156 81676 24892 81732
rect 24948 81676 27132 81732
rect 27188 81676 28364 81732
rect 28420 81676 28430 81732
rect 29698 81676 29708 81732
rect 29764 81676 31276 81732
rect 31332 81676 31342 81732
rect 34402 81676 34412 81732
rect 34468 81676 35308 81732
rect 35364 81676 35644 81732
rect 35700 81676 35710 81732
rect 19826 81508 19836 81564
rect 19892 81508 19940 81564
rect 19996 81508 20044 81564
rect 20100 81508 20110 81564
rect 27458 81452 27468 81508
rect 27524 81452 28140 81508
rect 28196 81452 28206 81508
rect 6514 81340 6524 81396
rect 6580 81340 7084 81396
rect 7140 81340 8988 81396
rect 9044 81340 9054 81396
rect 9874 81340 9884 81396
rect 9940 81340 10780 81396
rect 10836 81340 10846 81396
rect 13682 81340 13692 81396
rect 13748 81340 14476 81396
rect 14532 81340 14924 81396
rect 14980 81340 14990 81396
rect 15092 81340 27356 81396
rect 27412 81340 27422 81396
rect 30370 81340 30380 81396
rect 30436 81340 31612 81396
rect 31668 81340 31678 81396
rect 15092 81284 15148 81340
rect 4834 81228 4844 81284
rect 4900 81228 5628 81284
rect 5684 81228 5694 81284
rect 10210 81228 10220 81284
rect 10276 81228 15148 81284
rect 16482 81228 16492 81284
rect 16548 81228 18508 81284
rect 18564 81228 18574 81284
rect 20178 81228 20188 81284
rect 20244 81228 21980 81284
rect 22036 81228 22652 81284
rect 22708 81228 22718 81284
rect 23986 81228 23996 81284
rect 24052 81228 25004 81284
rect 25060 81228 25070 81284
rect 25442 81228 25452 81284
rect 25508 81228 25518 81284
rect 27682 81228 27692 81284
rect 27748 81228 29596 81284
rect 29652 81228 29662 81284
rect 7410 81116 7420 81172
rect 7476 81116 9772 81172
rect 9828 81116 9838 81172
rect 21858 81116 21868 81172
rect 21924 81116 23100 81172
rect 23156 81116 23166 81172
rect 25452 81060 25508 81228
rect 27122 81116 27132 81172
rect 27188 81116 28476 81172
rect 28532 81116 28542 81172
rect 9986 81004 9996 81060
rect 10052 81004 10668 81060
rect 10724 81004 10734 81060
rect 16370 81004 16380 81060
rect 16436 81004 17052 81060
rect 17108 81004 17388 81060
rect 17444 81004 17454 81060
rect 18610 81004 18620 81060
rect 18676 81004 20300 81060
rect 20356 81004 20366 81060
rect 22082 81004 22092 81060
rect 22148 81004 23324 81060
rect 23380 81004 26684 81060
rect 26740 81004 26750 81060
rect 26852 81004 29260 81060
rect 29316 81004 29326 81060
rect 13458 80892 13468 80948
rect 13524 80892 14028 80948
rect 14084 80892 14094 80948
rect 21970 80892 21980 80948
rect 22036 80892 25676 80948
rect 25732 80892 25742 80948
rect 26852 80836 26908 81004
rect 28466 80892 28476 80948
rect 28532 80892 29932 80948
rect 29988 80892 29998 80948
rect 22754 80780 22764 80836
rect 22820 80780 26572 80836
rect 26628 80780 26908 80836
rect 4466 80724 4476 80780
rect 4532 80724 4580 80780
rect 4636 80724 4684 80780
rect 4740 80724 4750 80780
rect 35186 80724 35196 80780
rect 35252 80724 35300 80780
rect 35356 80724 35404 80780
rect 35460 80724 35470 80780
rect 18834 80668 18844 80724
rect 18900 80668 20076 80724
rect 20132 80668 20142 80724
rect 24770 80668 24780 80724
rect 24836 80668 25452 80724
rect 25508 80668 25518 80724
rect 25890 80668 25900 80724
rect 25956 80668 26404 80724
rect 34150 80668 34188 80724
rect 34244 80668 34254 80724
rect 26348 80612 26404 80668
rect 17378 80556 17388 80612
rect 17444 80556 26012 80612
rect 26068 80556 26078 80612
rect 26338 80556 26348 80612
rect 26404 80556 26414 80612
rect 17042 80444 17052 80500
rect 17108 80444 23772 80500
rect 23828 80444 23838 80500
rect 24098 80444 24108 80500
rect 24164 80444 25788 80500
rect 25844 80444 25854 80500
rect 17826 80332 17836 80388
rect 17892 80332 20524 80388
rect 20580 80332 23660 80388
rect 23716 80332 23726 80388
rect 20850 80220 20860 80276
rect 20916 80220 22428 80276
rect 22484 80220 22494 80276
rect 19394 80108 19404 80164
rect 19460 80108 20076 80164
rect 20132 80108 20244 80164
rect 20626 80108 20636 80164
rect 20692 80108 22092 80164
rect 22148 80108 22158 80164
rect 20188 80052 20244 80108
rect 20188 79996 20972 80052
rect 21028 79996 21532 80052
rect 21588 79996 22316 80052
rect 22372 79996 22382 80052
rect 19826 79940 19836 79996
rect 19892 79940 19940 79996
rect 19996 79940 20044 79996
rect 20100 79940 20110 79996
rect 14140 79772 16268 79828
rect 16324 79772 16334 79828
rect 18050 79772 18060 79828
rect 18116 79772 22204 79828
rect 22260 79772 22270 79828
rect 14140 79604 14196 79772
rect 18284 79660 27692 79716
rect 27748 79660 27758 79716
rect 18284 79604 18340 79660
rect 10546 79548 10556 79604
rect 10612 79548 11564 79604
rect 11620 79548 13580 79604
rect 13636 79548 14140 79604
rect 14196 79548 14206 79604
rect 18274 79548 18284 79604
rect 18340 79548 18350 79604
rect 18610 79548 18620 79604
rect 18676 79548 23436 79604
rect 23492 79548 23502 79604
rect 23874 79548 23884 79604
rect 23940 79548 26124 79604
rect 26180 79548 26908 79604
rect 26964 79548 26974 79604
rect 5954 79436 5964 79492
rect 6020 79436 8988 79492
rect 9044 79436 9660 79492
rect 9716 79436 9726 79492
rect 16818 79436 16828 79492
rect 16884 79436 18060 79492
rect 18116 79436 23660 79492
rect 23716 79436 23726 79492
rect 24994 79436 25004 79492
rect 25060 79436 27244 79492
rect 27300 79436 27310 79492
rect 29362 79436 29372 79492
rect 29428 79436 30268 79492
rect 30324 79436 30334 79492
rect 27682 79324 27692 79380
rect 27748 79324 30940 79380
rect 30996 79324 31006 79380
rect 30454 79212 30492 79268
rect 30548 79212 30558 79268
rect 4466 79156 4476 79212
rect 4532 79156 4580 79212
rect 4636 79156 4684 79212
rect 4740 79156 4750 79212
rect 35186 79156 35196 79212
rect 35252 79156 35300 79212
rect 35356 79156 35404 79212
rect 35460 79156 35470 79212
rect 27010 79100 27020 79156
rect 27076 79100 27132 79156
rect 27188 79100 27198 79156
rect 17276 78988 17780 79044
rect 24322 78988 24332 79044
rect 24388 78988 25564 79044
rect 25620 78988 25630 79044
rect 27542 78988 27580 79044
rect 27636 78988 27646 79044
rect 17276 78932 17332 78988
rect 17724 78932 17780 78988
rect 5954 78876 5964 78932
rect 6020 78876 7084 78932
rect 7140 78876 7150 78932
rect 10658 78876 10668 78932
rect 10724 78876 17332 78932
rect 17490 78876 17500 78932
rect 17556 78876 17566 78932
rect 17724 78876 23884 78932
rect 23940 78876 23950 78932
rect 26898 78876 26908 78932
rect 26964 78876 27132 78932
rect 27188 78876 27916 78932
rect 27972 78876 27982 78932
rect 28130 78876 28140 78932
rect 28196 78876 29148 78932
rect 29204 78876 29214 78932
rect 29698 78876 29708 78932
rect 29764 78876 30604 78932
rect 30660 78876 32396 78932
rect 32452 78876 33292 78932
rect 33348 78876 33358 78932
rect 17500 78820 17556 78876
rect 6850 78764 6860 78820
rect 6916 78764 7532 78820
rect 7588 78764 11564 78820
rect 11620 78764 12460 78820
rect 12516 78764 12526 78820
rect 17500 78764 18396 78820
rect 18452 78764 20524 78820
rect 20580 78764 20590 78820
rect 23986 78764 23996 78820
rect 24052 78764 27020 78820
rect 27076 78764 27086 78820
rect 27234 78764 27244 78820
rect 27300 78764 28028 78820
rect 28084 78764 28094 78820
rect 28354 78764 28364 78820
rect 28420 78764 28700 78820
rect 28756 78764 29484 78820
rect 29540 78764 29550 78820
rect 30034 78764 30044 78820
rect 30100 78764 30492 78820
rect 30548 78764 30558 78820
rect 6514 78652 6524 78708
rect 6580 78652 20636 78708
rect 20692 78652 20702 78708
rect 22540 78652 23436 78708
rect 23492 78652 23502 78708
rect 25974 78652 26012 78708
rect 26068 78652 26078 78708
rect 31490 78652 31500 78708
rect 31556 78652 32060 78708
rect 32116 78652 32126 78708
rect 22540 78596 22596 78652
rect 7298 78540 7308 78596
rect 7364 78540 10220 78596
rect 10276 78540 10286 78596
rect 13458 78540 13468 78596
rect 13524 78540 15820 78596
rect 15876 78540 15886 78596
rect 20066 78540 20076 78596
rect 20132 78540 21644 78596
rect 21700 78540 22540 78596
rect 22596 78540 22606 78596
rect 22754 78540 22764 78596
rect 22820 78540 24332 78596
rect 24388 78540 24780 78596
rect 24836 78540 24846 78596
rect 25778 78540 25788 78596
rect 25844 78540 26684 78596
rect 26740 78540 26750 78596
rect 27458 78540 27468 78596
rect 27524 78540 28252 78596
rect 28308 78540 28318 78596
rect 29138 78540 29148 78596
rect 29204 78540 30156 78596
rect 30212 78540 30492 78596
rect 30548 78540 31836 78596
rect 31892 78540 31902 78596
rect 32722 78540 32732 78596
rect 32788 78540 34860 78596
rect 34916 78540 34926 78596
rect 35858 78540 35868 78596
rect 35924 78540 37996 78596
rect 38052 78540 38062 78596
rect 3602 78428 3612 78484
rect 3668 78428 6076 78484
rect 6132 78428 6142 78484
rect 19826 78372 19836 78428
rect 19892 78372 19940 78428
rect 19996 78372 20044 78428
rect 20100 78372 20110 78428
rect 16706 78316 16716 78372
rect 16772 78316 18732 78372
rect 18788 78316 18798 78372
rect 31714 78316 31724 78372
rect 31780 78316 32396 78372
rect 32452 78316 32462 78372
rect 11106 78204 11116 78260
rect 11172 78204 18620 78260
rect 18676 78204 19628 78260
rect 19684 78204 19694 78260
rect 28802 78204 28812 78260
rect 28868 78204 29260 78260
rect 29316 78204 32172 78260
rect 32228 78204 32238 78260
rect 35298 78204 35308 78260
rect 35364 78204 37324 78260
rect 37380 78204 37390 78260
rect 15810 78092 15820 78148
rect 15876 78092 17612 78148
rect 17668 78092 17678 78148
rect 25750 78092 25788 78148
rect 25844 78092 25854 78148
rect 26086 78092 26124 78148
rect 26180 78092 26190 78148
rect 30380 78092 31556 78148
rect 34626 78092 34636 78148
rect 34692 78092 35756 78148
rect 35812 78092 37100 78148
rect 37156 78092 37166 78148
rect 30380 78036 30436 78092
rect 31500 78036 31556 78092
rect 16706 77980 16716 78036
rect 16772 77980 17388 78036
rect 17444 77980 17454 78036
rect 22530 77980 22540 78036
rect 22596 77980 26348 78036
rect 26404 77980 28476 78036
rect 28532 77980 28542 78036
rect 30370 77980 30380 78036
rect 30436 77980 30446 78036
rect 31266 77980 31276 78036
rect 31332 77980 31342 78036
rect 31490 77980 31500 78036
rect 31556 77980 32844 78036
rect 32900 77980 32910 78036
rect 34402 77980 34412 78036
rect 34468 77980 35084 78036
rect 35140 77980 35150 78036
rect 35522 77980 35532 78036
rect 35588 77980 35598 78036
rect 35858 77980 35868 78036
rect 35924 77980 37212 78036
rect 37268 77980 37278 78036
rect 31276 77924 31332 77980
rect 35532 77924 35588 77980
rect 11330 77868 11340 77924
rect 11396 77868 12908 77924
rect 12964 77868 14140 77924
rect 14196 77868 14206 77924
rect 15250 77868 15260 77924
rect 15316 77868 16268 77924
rect 16324 77868 16828 77924
rect 16884 77868 16894 77924
rect 23762 77868 23772 77924
rect 23828 77868 25788 77924
rect 25844 77868 28028 77924
rect 28084 77868 28094 77924
rect 31276 77868 34076 77924
rect 34132 77868 34142 77924
rect 35532 77868 36092 77924
rect 36148 77868 36316 77924
rect 36372 77868 36382 77924
rect 31276 77812 31332 77868
rect 22082 77756 22092 77812
rect 22148 77756 27244 77812
rect 27300 77756 27310 77812
rect 30818 77756 30828 77812
rect 30884 77756 31332 77812
rect 35074 77756 35084 77812
rect 35140 77756 36540 77812
rect 36596 77756 36606 77812
rect 21858 77644 21868 77700
rect 21924 77644 25564 77700
rect 25620 77644 27020 77700
rect 27076 77644 27086 77700
rect 30258 77644 30268 77700
rect 30324 77644 33180 77700
rect 33236 77644 33246 77700
rect 4466 77588 4476 77644
rect 4532 77588 4580 77644
rect 4636 77588 4684 77644
rect 4740 77588 4750 77644
rect 35186 77588 35196 77644
rect 35252 77588 35300 77644
rect 35356 77588 35404 77644
rect 35460 77588 35470 77644
rect 25218 77532 25228 77588
rect 25284 77532 26684 77588
rect 26740 77532 26750 77588
rect 31014 77532 31052 77588
rect 31108 77532 31118 77588
rect 31602 77532 31612 77588
rect 31668 77532 34524 77588
rect 34580 77532 34590 77588
rect 35718 77532 35756 77588
rect 35812 77532 35822 77588
rect 6850 77420 6860 77476
rect 6916 77420 7308 77476
rect 7364 77420 7374 77476
rect 27010 77420 27020 77476
rect 27076 77420 27114 77476
rect 30930 77420 30940 77476
rect 30996 77420 31006 77476
rect 32050 77420 32060 77476
rect 32116 77420 33068 77476
rect 33124 77420 33134 77476
rect 34738 77420 34748 77476
rect 34804 77420 36204 77476
rect 36260 77420 36270 77476
rect 36642 77420 36652 77476
rect 36708 77420 37212 77476
rect 37268 77420 37884 77476
rect 37940 77420 37950 77476
rect 30940 77364 30996 77420
rect 6962 77308 6972 77364
rect 7028 77308 8372 77364
rect 12898 77308 12908 77364
rect 12964 77308 13804 77364
rect 13860 77308 13870 77364
rect 30940 77308 31164 77364
rect 31220 77308 31230 77364
rect 32386 77308 32396 77364
rect 32452 77308 35644 77364
rect 35700 77308 35710 77364
rect 8316 77252 8372 77308
rect 8316 77196 10108 77252
rect 10164 77196 10174 77252
rect 19506 77196 19516 77252
rect 19572 77196 26012 77252
rect 26068 77196 26908 77252
rect 29250 77196 29260 77252
rect 29316 77196 29326 77252
rect 29698 77196 29708 77252
rect 29764 77196 32172 77252
rect 32228 77196 32238 77252
rect 34402 77196 34412 77252
rect 34468 77196 36428 77252
rect 36484 77196 36876 77252
rect 36932 77196 36942 77252
rect 37426 77196 37436 77252
rect 37492 77196 38108 77252
rect 38164 77196 38174 77252
rect 26852 77140 26908 77196
rect 29260 77140 29316 77196
rect 12338 77084 12348 77140
rect 12404 77084 13692 77140
rect 13748 77084 14812 77140
rect 14868 77084 15148 77140
rect 15204 77084 16828 77140
rect 16884 77084 17948 77140
rect 18004 77084 18014 77140
rect 26852 77084 29316 77140
rect 31490 77084 31500 77140
rect 31556 77084 33292 77140
rect 33348 77084 33358 77140
rect 34178 77084 34188 77140
rect 34244 77084 36988 77140
rect 37044 77084 37054 77140
rect 15474 76972 15484 77028
rect 15540 76972 16044 77028
rect 16100 76972 17724 77028
rect 17780 76972 20244 77028
rect 27346 76972 27356 77028
rect 27412 76972 27468 77028
rect 27524 76972 27534 77028
rect 28578 76972 28588 77028
rect 28644 76972 29708 77028
rect 29764 76972 30380 77028
rect 30436 76972 30446 77028
rect 31266 76972 31276 77028
rect 31332 76972 34300 77028
rect 34356 76972 34366 77028
rect 35410 76972 35420 77028
rect 35476 76972 37100 77028
rect 37156 76972 37166 77028
rect 19826 76804 19836 76860
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 20100 76804 20110 76860
rect 20188 76804 20244 76972
rect 28588 76916 28644 76972
rect 26338 76860 26348 76916
rect 26404 76860 28644 76916
rect 31154 76860 31164 76916
rect 31220 76860 32060 76916
rect 32116 76860 32126 76916
rect 32386 76860 32396 76916
rect 32452 76860 33180 76916
rect 33236 76860 33246 76916
rect 33618 76860 33628 76916
rect 33684 76860 37660 76916
rect 37716 76860 37726 76916
rect 20188 76748 27804 76804
rect 27860 76748 27870 76804
rect 28354 76748 28364 76804
rect 28420 76748 30156 76804
rect 30212 76748 30222 76804
rect 31714 76748 31724 76804
rect 31780 76748 32508 76804
rect 32564 76748 32574 76804
rect 35410 76748 35420 76804
rect 35476 76748 36428 76804
rect 36484 76748 37212 76804
rect 37268 76748 37278 76804
rect 15922 76636 15932 76692
rect 15988 76636 16604 76692
rect 16660 76636 21644 76692
rect 21700 76636 21710 76692
rect 24546 76636 24556 76692
rect 24612 76636 25340 76692
rect 25396 76636 25406 76692
rect 26786 76636 26796 76692
rect 26852 76636 26908 76692
rect 26964 76636 26974 76692
rect 36092 76580 36148 76748
rect 8306 76524 8316 76580
rect 8372 76524 9548 76580
rect 9604 76524 9614 76580
rect 19618 76524 19628 76580
rect 19684 76524 20636 76580
rect 20692 76524 20702 76580
rect 24098 76524 24108 76580
rect 24164 76524 27244 76580
rect 27300 76524 27310 76580
rect 27458 76524 27468 76580
rect 27524 76524 27580 76580
rect 27636 76524 27646 76580
rect 30482 76524 30492 76580
rect 30548 76524 32956 76580
rect 33012 76524 33022 76580
rect 33516 76524 34412 76580
rect 34468 76524 34478 76580
rect 36082 76524 36092 76580
rect 36148 76524 36158 76580
rect 36306 76524 36316 76580
rect 36372 76524 37884 76580
rect 37940 76524 37950 76580
rect 33516 76468 33572 76524
rect 7634 76412 7644 76468
rect 7700 76412 9772 76468
rect 9828 76412 9838 76468
rect 10210 76412 10220 76468
rect 10276 76412 24220 76468
rect 24276 76412 24286 76468
rect 24658 76412 24668 76468
rect 24724 76412 25564 76468
rect 25620 76412 25630 76468
rect 27346 76412 27356 76468
rect 27412 76412 29596 76468
rect 29652 76412 29662 76468
rect 33506 76412 33516 76468
rect 33572 76412 33582 76468
rect 33954 76412 33964 76468
rect 34020 76412 35308 76468
rect 35364 76412 35374 76468
rect 36418 76412 36428 76468
rect 36484 76412 37100 76468
rect 37156 76412 37166 76468
rect 10322 76300 10332 76356
rect 10388 76300 10668 76356
rect 10724 76300 10734 76356
rect 11106 76300 11116 76356
rect 11172 76300 13468 76356
rect 13524 76300 13534 76356
rect 26002 76300 26012 76356
rect 26068 76300 26124 76356
rect 26180 76300 26190 76356
rect 27122 76300 27132 76356
rect 27188 76300 27916 76356
rect 27972 76300 27982 76356
rect 35746 76300 35756 76356
rect 35812 76300 37436 76356
rect 37492 76300 37502 76356
rect 11116 76244 11172 76300
rect 8754 76188 8764 76244
rect 8820 76188 11172 76244
rect 26786 76188 26796 76244
rect 26852 76188 28252 76244
rect 28308 76188 28318 76244
rect 29698 76188 29708 76244
rect 29764 76188 30380 76244
rect 30436 76188 30716 76244
rect 30772 76188 30782 76244
rect 33394 76188 33404 76244
rect 33460 76188 34188 76244
rect 34244 76188 34254 76244
rect 34514 76188 34524 76244
rect 34580 76188 35532 76244
rect 35588 76188 35598 76244
rect 4466 76020 4476 76076
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4740 76020 4750 76076
rect 35186 76020 35196 76076
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35460 76020 35470 76076
rect 5954 75964 5964 76020
rect 6020 75964 7308 76020
rect 7364 75964 7374 76020
rect 15026 75964 15036 76020
rect 15092 75964 19292 76020
rect 19348 75964 19358 76020
rect 29138 75964 29148 76020
rect 29204 75964 31052 76020
rect 31108 75964 31118 76020
rect 6850 75852 6860 75908
rect 6916 75852 21980 75908
rect 22036 75852 22046 75908
rect 24546 75852 24556 75908
rect 24612 75852 26348 75908
rect 26404 75852 26684 75908
rect 26740 75852 28700 75908
rect 28756 75852 28766 75908
rect 34066 75852 34076 75908
rect 34132 75852 37996 75908
rect 38052 75852 38062 75908
rect 4834 75740 4844 75796
rect 4900 75740 7644 75796
rect 7700 75740 7710 75796
rect 27794 75740 27804 75796
rect 27860 75740 29260 75796
rect 29316 75740 30156 75796
rect 30212 75740 30380 75796
rect 30436 75740 30446 75796
rect 32274 75740 32284 75796
rect 32340 75740 37100 75796
rect 37156 75740 37166 75796
rect 4274 75628 4284 75684
rect 4340 75628 6300 75684
rect 6356 75628 6366 75684
rect 14466 75628 14476 75684
rect 14532 75628 15932 75684
rect 15988 75628 15998 75684
rect 24434 75628 24444 75684
rect 24500 75628 27580 75684
rect 27636 75628 27646 75684
rect 30594 75628 30604 75684
rect 30660 75628 31948 75684
rect 32004 75628 32014 75684
rect 34402 75628 34412 75684
rect 34468 75628 36092 75684
rect 36148 75628 37212 75684
rect 37268 75628 37278 75684
rect 13906 75516 13916 75572
rect 13972 75516 18060 75572
rect 18116 75516 18126 75572
rect 19058 75516 19068 75572
rect 19124 75516 20412 75572
rect 20468 75516 20478 75572
rect 27234 75516 27244 75572
rect 27300 75516 28364 75572
rect 28420 75516 29820 75572
rect 29876 75516 29886 75572
rect 30930 75516 30940 75572
rect 30996 75516 31836 75572
rect 31892 75516 31902 75572
rect 32386 75516 32396 75572
rect 32452 75516 32462 75572
rect 33506 75516 33516 75572
rect 33572 75516 34972 75572
rect 35028 75516 36988 75572
rect 37044 75516 37054 75572
rect 15036 75460 15092 75516
rect 32396 75460 32452 75516
rect 15026 75404 15036 75460
rect 15092 75404 15102 75460
rect 30034 75404 30044 75460
rect 30100 75404 31612 75460
rect 31668 75404 32452 75460
rect 33730 75404 33740 75460
rect 33796 75404 34636 75460
rect 34692 75404 34702 75460
rect 35298 75404 35308 75460
rect 35364 75404 35756 75460
rect 35812 75404 36092 75460
rect 36148 75404 36158 75460
rect 35308 75348 35364 75404
rect 25778 75292 25788 75348
rect 25844 75292 26236 75348
rect 26292 75292 27804 75348
rect 27860 75292 27870 75348
rect 33282 75292 33292 75348
rect 33348 75292 33964 75348
rect 34020 75292 35364 75348
rect 35970 75292 35980 75348
rect 36036 75292 36046 75348
rect 19826 75236 19836 75292
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 20100 75236 20110 75292
rect 30454 75180 30492 75236
rect 30548 75180 30558 75236
rect 31042 75180 31052 75236
rect 31108 75180 31836 75236
rect 31892 75180 31902 75236
rect 35980 75124 36036 75292
rect 16034 75068 16044 75124
rect 16100 75068 17500 75124
rect 17556 75068 17566 75124
rect 17714 75068 17724 75124
rect 17780 75068 18172 75124
rect 18228 75068 18238 75124
rect 22866 75068 22876 75124
rect 22932 75068 22942 75124
rect 25218 75068 25228 75124
rect 25284 75068 25676 75124
rect 25732 75068 25742 75124
rect 31714 75068 31724 75124
rect 31780 75068 32508 75124
rect 32564 75068 32574 75124
rect 34066 75068 34076 75124
rect 34132 75068 35196 75124
rect 35252 75068 35262 75124
rect 35970 75068 35980 75124
rect 36036 75068 36046 75124
rect 36306 75068 36316 75124
rect 36372 75068 37436 75124
rect 37492 75068 37502 75124
rect 22876 75012 22932 75068
rect 36316 75012 36372 75068
rect 8306 74956 8316 75012
rect 8372 74956 8764 75012
rect 8820 74956 22932 75012
rect 23762 74956 23772 75012
rect 23828 74956 24332 75012
rect 24388 74956 24398 75012
rect 25330 74956 25340 75012
rect 25396 74956 27132 75012
rect 27188 74956 27198 75012
rect 34626 74956 34636 75012
rect 34692 74956 34972 75012
rect 35028 74956 36372 75012
rect 39600 74900 40000 74928
rect 7298 74844 7308 74900
rect 7364 74844 7756 74900
rect 7812 74844 8428 74900
rect 8484 74844 8494 74900
rect 22978 74844 22988 74900
rect 23044 74844 23884 74900
rect 23940 74844 23950 74900
rect 25218 74844 25228 74900
rect 25284 74844 26460 74900
rect 26516 74844 27020 74900
rect 27076 74844 27086 74900
rect 29586 74844 29596 74900
rect 29652 74844 30604 74900
rect 30660 74844 30670 74900
rect 38210 74844 38220 74900
rect 38276 74844 40000 74900
rect 39600 74816 40000 74844
rect 4162 74732 4172 74788
rect 4228 74732 4396 74788
rect 4452 74732 4462 74788
rect 6514 74732 6524 74788
rect 6580 74732 8092 74788
rect 8148 74732 8158 74788
rect 13682 74732 13692 74788
rect 13748 74732 15260 74788
rect 15316 74732 15326 74788
rect 18050 74732 18060 74788
rect 18116 74732 19740 74788
rect 19796 74732 19806 74788
rect 28466 74732 28476 74788
rect 28532 74732 29260 74788
rect 29316 74732 29326 74788
rect 32722 74732 32732 74788
rect 32788 74732 37660 74788
rect 37716 74732 37726 74788
rect 0 74676 400 74704
rect 0 74620 4844 74676
rect 4900 74620 4910 74676
rect 10882 74620 10892 74676
rect 10948 74620 11452 74676
rect 11508 74620 11518 74676
rect 35718 74620 35756 74676
rect 35812 74620 36428 74676
rect 36484 74620 36876 74676
rect 36932 74620 36942 74676
rect 0 74592 400 74620
rect 4466 74452 4476 74508
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4740 74452 4750 74508
rect 35186 74452 35196 74508
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35460 74452 35470 74508
rect 7074 74396 7084 74452
rect 7140 74396 7868 74452
rect 7924 74396 7934 74452
rect 5282 74284 5292 74340
rect 5348 74284 7196 74340
rect 7252 74284 7262 74340
rect 20066 74284 20076 74340
rect 20132 74284 21420 74340
rect 21476 74284 22540 74340
rect 22596 74284 22606 74340
rect 35298 74284 35308 74340
rect 35364 74284 35756 74340
rect 35812 74284 35822 74340
rect 2146 74172 2156 74228
rect 2212 74172 3388 74228
rect 19058 74172 19068 74228
rect 19124 74172 21644 74228
rect 21700 74172 21710 74228
rect 29810 74172 29820 74228
rect 29876 74172 30268 74228
rect 30324 74172 30716 74228
rect 30772 74172 31500 74228
rect 31556 74172 31566 74228
rect 34402 74172 34412 74228
rect 34468 74172 35644 74228
rect 35700 74172 35710 74228
rect 3332 74004 3388 74172
rect 4162 74060 4172 74116
rect 4228 74060 6748 74116
rect 6804 74060 6814 74116
rect 17938 74060 17948 74116
rect 18004 74060 19852 74116
rect 19908 74060 23100 74116
rect 23156 74060 23166 74116
rect 27794 74060 27804 74116
rect 27860 74060 28364 74116
rect 28420 74060 28430 74116
rect 29250 74060 29260 74116
rect 29316 74060 32732 74116
rect 32788 74060 32798 74116
rect 35410 74060 35420 74116
rect 35476 74060 36092 74116
rect 36148 74060 36158 74116
rect 3332 73948 3724 74004
rect 3780 73948 5852 74004
rect 5908 73948 5918 74004
rect 6972 73948 7196 74004
rect 7252 73948 7980 74004
rect 8036 73948 8046 74004
rect 15026 73948 15036 74004
rect 15092 73948 15372 74004
rect 15428 73948 15438 74004
rect 15922 73948 15932 74004
rect 15988 73948 17220 74004
rect 19730 73948 19740 74004
rect 19796 73948 20524 74004
rect 20580 73948 22204 74004
rect 22260 73948 22270 74004
rect 31490 73948 31500 74004
rect 31556 73948 31948 74004
rect 6972 73892 7028 73948
rect 5730 73836 5740 73892
rect 5796 73836 6188 73892
rect 6244 73836 6636 73892
rect 6692 73836 7028 73892
rect 17164 73892 17220 73948
rect 17164 73836 17500 73892
rect 17556 73836 18844 73892
rect 18900 73836 19516 73892
rect 19572 73836 19582 73892
rect 31892 73836 31948 73948
rect 32004 73836 32014 73892
rect 35718 73836 35756 73892
rect 35812 73836 35822 73892
rect 19826 73668 19836 73724
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 20100 73668 20110 73724
rect 28130 73612 28140 73668
rect 28196 73612 29260 73668
rect 29316 73612 29326 73668
rect 27570 73500 27580 73556
rect 27636 73500 30492 73556
rect 30548 73500 30558 73556
rect 34066 73500 34076 73556
rect 34132 73500 34412 73556
rect 34468 73500 34478 73556
rect 24322 73388 24332 73444
rect 24388 73388 29820 73444
rect 29876 73388 31052 73444
rect 31108 73388 31118 73444
rect 28354 73276 28364 73332
rect 28420 73276 29036 73332
rect 29092 73276 29102 73332
rect 17714 73164 17724 73220
rect 17780 73164 18396 73220
rect 18452 73164 21084 73220
rect 21140 73164 24668 73220
rect 24724 73164 24734 73220
rect 26226 73164 26236 73220
rect 26292 73164 28252 73220
rect 28308 73164 28318 73220
rect 26114 73052 26124 73108
rect 26180 73052 26908 73108
rect 26964 73052 27804 73108
rect 27860 73052 28028 73108
rect 28084 73052 29260 73108
rect 29316 73052 29326 73108
rect 4466 72884 4476 72940
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4740 72884 4750 72940
rect 35186 72884 35196 72940
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35460 72884 35470 72940
rect 22530 72716 22540 72772
rect 22596 72716 23548 72772
rect 23604 72716 23614 72772
rect 24770 72716 24780 72772
rect 24836 72716 25564 72772
rect 25620 72716 25630 72772
rect 25218 72604 25228 72660
rect 25284 72604 29820 72660
rect 29876 72604 29886 72660
rect 19954 72492 19964 72548
rect 20020 72492 20412 72548
rect 20468 72492 27804 72548
rect 27860 72492 31276 72548
rect 31332 72492 31342 72548
rect 26786 72380 26796 72436
rect 26852 72380 28140 72436
rect 28196 72380 28206 72436
rect 7410 72268 7420 72324
rect 7476 72268 8092 72324
rect 8148 72268 8158 72324
rect 10994 72268 11004 72324
rect 11060 72268 11564 72324
rect 11620 72268 11630 72324
rect 33730 72268 33740 72324
rect 33796 72268 35644 72324
rect 35700 72268 35710 72324
rect 36054 72268 36092 72324
rect 36148 72268 36764 72324
rect 36820 72268 36830 72324
rect 13906 72156 13916 72212
rect 13972 72156 18844 72212
rect 18900 72156 18910 72212
rect 23986 72156 23996 72212
rect 24052 72156 25004 72212
rect 25060 72156 25070 72212
rect 33618 72156 33628 72212
rect 33684 72156 34076 72212
rect 34132 72156 34142 72212
rect 19826 72100 19836 72156
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 20100 72100 20110 72156
rect 32162 72044 32172 72100
rect 32228 72044 33852 72100
rect 33908 72044 33918 72100
rect 32386 71932 32396 71988
rect 32452 71932 33740 71988
rect 33796 71932 33806 71988
rect 7522 71820 7532 71876
rect 7588 71820 8540 71876
rect 8596 71820 8606 71876
rect 34402 71820 34412 71876
rect 34468 71820 34748 71876
rect 34804 71820 34814 71876
rect 11106 71708 11116 71764
rect 11172 71708 14476 71764
rect 14532 71708 15036 71764
rect 15092 71708 15102 71764
rect 16818 71708 16828 71764
rect 16884 71708 17500 71764
rect 17556 71708 19180 71764
rect 19236 71708 21868 71764
rect 21924 71708 21934 71764
rect 22866 71596 22876 71652
rect 22932 71596 24668 71652
rect 24724 71596 26012 71652
rect 26068 71596 28140 71652
rect 28196 71596 28206 71652
rect 36306 71596 36316 71652
rect 36372 71596 37212 71652
rect 37268 71596 37660 71652
rect 37716 71596 37726 71652
rect 29362 71484 29372 71540
rect 29428 71484 30268 71540
rect 30324 71484 30334 71540
rect 33282 71484 33292 71540
rect 33348 71484 35532 71540
rect 35588 71484 35598 71540
rect 12674 71372 12684 71428
rect 12740 71372 13468 71428
rect 13524 71372 13534 71428
rect 4466 71316 4476 71372
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4740 71316 4750 71372
rect 35186 71316 35196 71372
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35460 71316 35470 71372
rect 28914 71148 28924 71204
rect 28980 71148 29596 71204
rect 29652 71148 32508 71204
rect 32564 71148 32574 71204
rect 33618 71148 33628 71204
rect 33684 71148 34636 71204
rect 34692 71148 34702 71204
rect 29922 71036 29932 71092
rect 29988 71036 34188 71092
rect 34244 71036 35308 71092
rect 35364 71036 36316 71092
rect 36372 71036 36382 71092
rect 24322 70924 24332 70980
rect 24388 70924 25564 70980
rect 25620 70924 25630 70980
rect 28018 70924 28028 70980
rect 28084 70924 28252 70980
rect 28308 70924 29372 70980
rect 29428 70924 29438 70980
rect 30594 70924 30604 70980
rect 30660 70924 32732 70980
rect 32788 70924 32798 70980
rect 32956 70924 37212 70980
rect 37268 70924 37278 70980
rect 32956 70868 33012 70924
rect 9538 70812 9548 70868
rect 9604 70812 9996 70868
rect 10052 70812 11900 70868
rect 11956 70812 11966 70868
rect 30258 70812 30268 70868
rect 30324 70812 30716 70868
rect 30772 70812 31052 70868
rect 31108 70812 32284 70868
rect 32340 70812 33012 70868
rect 33394 70812 33404 70868
rect 33460 70812 35420 70868
rect 35476 70812 35486 70868
rect 26852 70700 27692 70756
rect 27748 70700 31724 70756
rect 31780 70700 31790 70756
rect 26852 70644 26908 70700
rect 12898 70588 12908 70644
rect 12964 70588 14028 70644
rect 14084 70588 15484 70644
rect 15540 70588 15550 70644
rect 26450 70588 26460 70644
rect 26516 70588 26908 70644
rect 27122 70588 27132 70644
rect 27188 70588 29820 70644
rect 29876 70588 29886 70644
rect 30370 70588 30380 70644
rect 30436 70588 31052 70644
rect 31108 70588 31118 70644
rect 34738 70588 34748 70644
rect 34804 70588 36092 70644
rect 36148 70588 38220 70644
rect 38276 70588 38286 70644
rect 19826 70532 19836 70588
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 20100 70532 20110 70588
rect 25890 70476 25900 70532
rect 25956 70476 27468 70532
rect 27524 70476 27534 70532
rect 25330 70364 25340 70420
rect 25396 70364 27804 70420
rect 27860 70364 27870 70420
rect 28130 70364 28140 70420
rect 28196 70364 28206 70420
rect 29110 70364 29148 70420
rect 29204 70364 29214 70420
rect 31826 70364 31836 70420
rect 31892 70364 34076 70420
rect 34132 70364 34142 70420
rect 28140 70308 28196 70364
rect 14578 70252 14588 70308
rect 14644 70252 15708 70308
rect 15764 70252 16604 70308
rect 16660 70252 16670 70308
rect 25778 70252 25788 70308
rect 25844 70252 28196 70308
rect 15250 70140 15260 70196
rect 15316 70140 15596 70196
rect 15652 70140 15662 70196
rect 18946 70140 18956 70196
rect 19012 70140 22316 70196
rect 22372 70140 22382 70196
rect 28130 70140 28140 70196
rect 28196 70140 29708 70196
rect 29764 70140 29774 70196
rect 30706 70140 30716 70196
rect 30772 70140 31164 70196
rect 31220 70140 31836 70196
rect 31892 70140 34412 70196
rect 34468 70140 34478 70196
rect 36082 70140 36092 70196
rect 36148 70140 37324 70196
rect 37380 70140 37390 70196
rect 6738 70028 6748 70084
rect 6804 70028 8764 70084
rect 8820 70028 9548 70084
rect 9604 70028 9614 70084
rect 9874 70028 9884 70084
rect 9940 70028 10332 70084
rect 10388 70028 10398 70084
rect 18498 70028 18508 70084
rect 18564 70028 19628 70084
rect 19684 70028 19694 70084
rect 10668 69916 11228 69972
rect 11284 69916 13692 69972
rect 13748 69916 13758 69972
rect 26786 69916 26796 69972
rect 26852 69916 27356 69972
rect 27412 69916 28476 69972
rect 28532 69916 28542 69972
rect 33394 69916 33404 69972
rect 33460 69916 36876 69972
rect 36932 69916 36942 69972
rect 4466 69748 4476 69804
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4740 69748 4750 69804
rect 10668 69748 10724 69916
rect 35186 69748 35196 69804
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35460 69748 35470 69804
rect 10658 69692 10668 69748
rect 10724 69692 10734 69748
rect 29250 69692 29260 69748
rect 29316 69692 30940 69748
rect 30996 69692 33068 69748
rect 33124 69692 33134 69748
rect 28354 69580 28364 69636
rect 28420 69580 29596 69636
rect 29652 69580 29662 69636
rect 11890 69468 11900 69524
rect 11956 69468 14028 69524
rect 14084 69468 14476 69524
rect 14532 69468 14812 69524
rect 14868 69468 16268 69524
rect 16324 69468 16334 69524
rect 27906 69468 27916 69524
rect 27972 69468 29372 69524
rect 29428 69468 30492 69524
rect 30548 69468 30558 69524
rect 26114 69356 26124 69412
rect 26180 69356 26684 69412
rect 26740 69356 29148 69412
rect 29204 69356 32284 69412
rect 32340 69356 32350 69412
rect 35074 69356 35084 69412
rect 35140 69356 35868 69412
rect 35924 69356 35934 69412
rect 27458 69244 27468 69300
rect 27524 69244 27916 69300
rect 27972 69244 28252 69300
rect 28308 69244 28318 69300
rect 5282 69132 5292 69188
rect 5348 69132 5964 69188
rect 6020 69132 6636 69188
rect 6692 69132 9660 69188
rect 9716 69132 9726 69188
rect 19826 68964 19836 69020
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 20100 68964 20110 69020
rect 5506 68908 5516 68964
rect 5572 68908 6076 68964
rect 6132 68908 7084 68964
rect 7140 68908 7150 68964
rect 30370 68908 30380 68964
rect 30436 68908 31164 68964
rect 31220 68908 31230 68964
rect 34962 68908 34972 68964
rect 35028 68908 37324 68964
rect 37380 68908 37884 68964
rect 37940 68908 37950 68964
rect 35532 68852 35588 68908
rect 5058 68796 5068 68852
rect 5124 68796 6188 68852
rect 6244 68796 6254 68852
rect 14914 68796 14924 68852
rect 14980 68796 15148 68852
rect 15204 68796 15820 68852
rect 15876 68796 16940 68852
rect 16996 68796 17500 68852
rect 17556 68796 18844 68852
rect 18900 68796 18910 68852
rect 32946 68796 32956 68852
rect 33012 68796 33740 68852
rect 33796 68796 33806 68852
rect 35522 68796 35532 68852
rect 35588 68796 35598 68852
rect 10546 68684 10556 68740
rect 10612 68684 10622 68740
rect 14354 68684 14364 68740
rect 14420 68684 15260 68740
rect 15316 68684 20748 68740
rect 20804 68684 20814 68740
rect 21046 68684 21084 68740
rect 21140 68684 21150 68740
rect 30034 68684 30044 68740
rect 30100 68684 32060 68740
rect 32116 68684 32126 68740
rect 33058 68684 33068 68740
rect 33124 68684 34300 68740
rect 34356 68684 34366 68740
rect 10556 68628 10612 68684
rect 33068 68628 33124 68684
rect 4498 68572 4508 68628
rect 4564 68572 5628 68628
rect 5684 68572 10612 68628
rect 30706 68572 30716 68628
rect 30772 68572 33124 68628
rect 3826 68460 3836 68516
rect 3892 68460 9548 68516
rect 9604 68460 9614 68516
rect 10098 68460 10108 68516
rect 10164 68460 10892 68516
rect 10948 68460 10958 68516
rect 28466 68460 28476 68516
rect 28532 68460 29036 68516
rect 29092 68460 29260 68516
rect 29316 68460 29326 68516
rect 29698 68460 29708 68516
rect 29764 68460 30044 68516
rect 30100 68460 30110 68516
rect 31938 68460 31948 68516
rect 32004 68460 32396 68516
rect 32452 68460 33628 68516
rect 33684 68460 33694 68516
rect 10108 68404 10164 68460
rect 8978 68348 8988 68404
rect 9044 68348 10164 68404
rect 13458 68348 13468 68404
rect 13524 68348 15372 68404
rect 15428 68348 16156 68404
rect 16212 68348 16222 68404
rect 31826 68348 31836 68404
rect 31892 68348 33852 68404
rect 33908 68348 33918 68404
rect 6178 68236 6188 68292
rect 6244 68236 9100 68292
rect 9156 68236 9166 68292
rect 9314 68236 9324 68292
rect 9380 68236 9884 68292
rect 9940 68236 10556 68292
rect 10612 68236 10622 68292
rect 29558 68236 29596 68292
rect 29652 68236 29662 68292
rect 4466 68180 4476 68236
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4740 68180 4750 68236
rect 35186 68180 35196 68236
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35460 68180 35470 68236
rect 6850 68124 6860 68180
rect 6916 68124 7644 68180
rect 7700 68124 7710 68180
rect 27682 68124 27692 68180
rect 27748 68124 29708 68180
rect 29764 68124 29774 68180
rect 33394 68124 33404 68180
rect 33460 68124 34188 68180
rect 34244 68124 34254 68180
rect 33058 68012 33068 68068
rect 33124 68012 34412 68068
rect 34468 68012 34478 68068
rect 18610 67900 18620 67956
rect 18676 67900 20188 67956
rect 20244 67900 21420 67956
rect 21476 67900 22428 67956
rect 22484 67900 22494 67956
rect 28578 67900 28588 67956
rect 28644 67900 29820 67956
rect 29876 67900 31724 67956
rect 31780 67900 31790 67956
rect 33730 67900 33740 67956
rect 33796 67900 37324 67956
rect 37380 67900 37390 67956
rect 32946 67788 32956 67844
rect 33012 67788 36092 67844
rect 36148 67788 37212 67844
rect 37268 67788 37278 67844
rect 16146 67676 16156 67732
rect 16212 67676 16828 67732
rect 16884 67676 17612 67732
rect 17668 67676 21644 67732
rect 21700 67676 21710 67732
rect 19394 67564 19404 67620
rect 19460 67564 21532 67620
rect 21588 67564 21598 67620
rect 36082 67564 36092 67620
rect 36148 67564 36764 67620
rect 36820 67564 36830 67620
rect 10546 67452 10556 67508
rect 10612 67452 11676 67508
rect 11732 67452 11742 67508
rect 19826 67396 19836 67452
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 20100 67396 20110 67452
rect 32498 67228 32508 67284
rect 32564 67228 33404 67284
rect 33460 67228 35308 67284
rect 35364 67228 36988 67284
rect 37044 67228 37436 67284
rect 37492 67228 37502 67284
rect 20066 67116 20076 67172
rect 20132 67116 22316 67172
rect 22372 67116 22382 67172
rect 29586 67116 29596 67172
rect 29652 67116 30492 67172
rect 30548 67116 31164 67172
rect 31220 67116 31230 67172
rect 15026 67004 15036 67060
rect 15092 67004 15484 67060
rect 15540 67004 15550 67060
rect 17938 67004 17948 67060
rect 18004 67004 18620 67060
rect 18676 67004 18956 67060
rect 19012 67004 19022 67060
rect 5058 66892 5068 66948
rect 5124 66892 5852 66948
rect 5908 66892 5918 66948
rect 17378 66892 17388 66948
rect 17444 66892 18172 66948
rect 18228 66892 18238 66948
rect 22092 66724 22148 67116
rect 29596 67060 29652 67116
rect 29138 67004 29148 67060
rect 29204 67004 29652 67060
rect 23202 66892 23212 66948
rect 23268 66892 30044 66948
rect 30100 66892 30110 66948
rect 29474 66780 29484 66836
rect 29540 66780 30940 66836
rect 30996 66780 31006 66836
rect 22082 66668 22092 66724
rect 22148 66668 26012 66724
rect 26068 66668 26078 66724
rect 4466 66612 4476 66668
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4740 66612 4750 66668
rect 35186 66612 35196 66668
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35460 66612 35470 66668
rect 15474 66556 15484 66612
rect 15540 66556 24780 66612
rect 24836 66556 24846 66612
rect 8754 66444 8764 66500
rect 8820 66444 9996 66500
rect 10052 66444 10062 66500
rect 18610 66444 18620 66500
rect 18676 66444 19180 66500
rect 19236 66444 19246 66500
rect 19394 66444 19404 66500
rect 19460 66444 19470 66500
rect 19404 66388 19460 66444
rect 3602 66332 3612 66388
rect 3668 66332 4396 66388
rect 4452 66332 5068 66388
rect 5124 66332 10668 66388
rect 10724 66332 10734 66388
rect 18162 66332 18172 66388
rect 18228 66332 18732 66388
rect 18788 66332 19460 66388
rect 21410 66332 21420 66388
rect 21476 66332 22316 66388
rect 22372 66332 22382 66388
rect 26002 66332 26012 66388
rect 26068 66332 27020 66388
rect 27076 66332 27086 66388
rect 33618 66332 33628 66388
rect 33684 66332 34636 66388
rect 34692 66332 34702 66388
rect 8754 66220 8764 66276
rect 8820 66220 9324 66276
rect 9380 66220 10220 66276
rect 10276 66220 11116 66276
rect 11172 66220 11900 66276
rect 11956 66220 11966 66276
rect 16482 66220 16492 66276
rect 16548 66220 19292 66276
rect 19348 66220 20412 66276
rect 20468 66220 20478 66276
rect 33282 66220 33292 66276
rect 33348 66220 35420 66276
rect 35476 66220 35486 66276
rect 36194 66220 36204 66276
rect 36260 66220 36270 66276
rect 36204 66164 36260 66220
rect 16370 66108 16380 66164
rect 16436 66108 17948 66164
rect 18004 66108 26348 66164
rect 26404 66108 26414 66164
rect 30706 66108 30716 66164
rect 30772 66108 30940 66164
rect 30996 66108 31276 66164
rect 31332 66108 31836 66164
rect 31892 66108 31902 66164
rect 33506 66108 33516 66164
rect 33572 66108 34748 66164
rect 34804 66108 34814 66164
rect 34962 66108 34972 66164
rect 35028 66108 36260 66164
rect 3714 65996 3724 66052
rect 3780 65996 4284 66052
rect 4340 65996 4350 66052
rect 9650 65996 9660 66052
rect 9716 65996 9726 66052
rect 10546 65996 10556 66052
rect 10612 65996 20524 66052
rect 20580 65996 20590 66052
rect 28802 65996 28812 66052
rect 28868 65996 29708 66052
rect 29764 65996 29774 66052
rect 30370 65996 30380 66052
rect 30436 65996 31164 66052
rect 31220 65996 31230 66052
rect 9660 65828 9716 65996
rect 19826 65828 19836 65884
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 20100 65828 20110 65884
rect 9660 65772 18844 65828
rect 18900 65772 18910 65828
rect 11442 65660 11452 65716
rect 11508 65660 19516 65716
rect 19572 65660 19582 65716
rect 33282 65660 33292 65716
rect 33348 65660 37548 65716
rect 37604 65660 37614 65716
rect 16258 65548 16268 65604
rect 16324 65548 17500 65604
rect 17556 65548 17566 65604
rect 30930 65548 30940 65604
rect 30996 65548 33628 65604
rect 33684 65548 33694 65604
rect 6514 65436 6524 65492
rect 6580 65436 7084 65492
rect 7140 65436 7150 65492
rect 14018 65436 14028 65492
rect 14084 65436 15596 65492
rect 15652 65436 15662 65492
rect 21186 65436 21196 65492
rect 21252 65436 23212 65492
rect 23268 65436 23278 65492
rect 23986 65436 23996 65492
rect 24052 65436 24892 65492
rect 24948 65436 25228 65492
rect 25284 65436 25294 65492
rect 29586 65436 29596 65492
rect 29652 65436 30604 65492
rect 30660 65436 30670 65492
rect 33394 65436 33404 65492
rect 33460 65436 34188 65492
rect 34244 65436 34254 65492
rect 34626 65436 34636 65492
rect 34692 65436 35868 65492
rect 35924 65436 35934 65492
rect 12450 65324 12460 65380
rect 12516 65324 13580 65380
rect 13636 65324 13646 65380
rect 19394 65324 19404 65380
rect 19460 65324 21308 65380
rect 21364 65324 21374 65380
rect 22306 65324 22316 65380
rect 22372 65324 24220 65380
rect 24276 65324 24668 65380
rect 24724 65324 25116 65380
rect 25172 65324 25182 65380
rect 25554 65324 25564 65380
rect 25620 65324 26236 65380
rect 26292 65324 26684 65380
rect 26740 65324 26750 65380
rect 31378 65324 31388 65380
rect 31444 65324 31612 65380
rect 31668 65324 31678 65380
rect 33506 65324 33516 65380
rect 33572 65324 36764 65380
rect 36820 65324 37324 65380
rect 37380 65324 37390 65380
rect 3826 65212 3836 65268
rect 3892 65212 4508 65268
rect 4564 65212 4574 65268
rect 21970 65212 21980 65268
rect 22036 65212 22876 65268
rect 22932 65212 22942 65268
rect 24098 65212 24108 65268
rect 24164 65212 24892 65268
rect 24948 65212 25340 65268
rect 25396 65212 25406 65268
rect 32386 65212 32396 65268
rect 32452 65212 33852 65268
rect 33908 65212 33918 65268
rect 35186 65212 35196 65268
rect 35252 65212 37884 65268
rect 37940 65212 37950 65268
rect 4466 65044 4476 65100
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4740 65044 4750 65100
rect 35186 65044 35196 65100
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35460 65044 35470 65100
rect 35634 64988 35644 65044
rect 35700 64988 36988 65044
rect 37044 64988 37054 65044
rect 12450 64876 12460 64932
rect 12516 64876 13468 64932
rect 13524 64876 13534 64932
rect 28578 64876 28588 64932
rect 28644 64876 29484 64932
rect 29540 64876 29550 64932
rect 32498 64876 32508 64932
rect 32564 64876 33404 64932
rect 33460 64876 33470 64932
rect 0 64820 400 64848
rect 0 64764 6748 64820
rect 6804 64764 6814 64820
rect 13010 64764 13020 64820
rect 13076 64764 13692 64820
rect 13748 64764 14364 64820
rect 14420 64764 14430 64820
rect 36306 64764 36316 64820
rect 36372 64764 36988 64820
rect 37044 64764 37054 64820
rect 0 64736 400 64764
rect 13794 64652 13804 64708
rect 13860 64652 14028 64708
rect 14084 64652 14094 64708
rect 20738 64652 20748 64708
rect 20804 64652 24108 64708
rect 24164 64652 24174 64708
rect 32610 64652 32620 64708
rect 32676 64652 35868 64708
rect 35924 64652 35934 64708
rect 4162 64540 4172 64596
rect 4228 64540 4844 64596
rect 4900 64540 4910 64596
rect 21634 64540 21644 64596
rect 21700 64540 22540 64596
rect 22596 64540 22606 64596
rect 23874 64540 23884 64596
rect 23940 64540 24668 64596
rect 24724 64540 24734 64596
rect 27794 64540 27804 64596
rect 27860 64540 29260 64596
rect 29316 64540 31388 64596
rect 31444 64540 31454 64596
rect 34290 64540 34300 64596
rect 34356 64540 34860 64596
rect 34916 64540 37436 64596
rect 37492 64540 37502 64596
rect 5282 64428 5292 64484
rect 5348 64428 7532 64484
rect 7588 64428 8204 64484
rect 8260 64428 8270 64484
rect 12114 64428 12124 64484
rect 12180 64428 14028 64484
rect 14084 64428 14094 64484
rect 18610 64428 18620 64484
rect 18676 64428 21532 64484
rect 21588 64428 21598 64484
rect 26852 64372 26908 64484
rect 26964 64428 26974 64484
rect 29474 64428 29484 64484
rect 29540 64428 30044 64484
rect 30100 64428 30828 64484
rect 30884 64428 30894 64484
rect 32274 64428 32284 64484
rect 32340 64428 36204 64484
rect 36260 64428 36270 64484
rect 11890 64316 11900 64372
rect 11956 64316 13692 64372
rect 13748 64316 13758 64372
rect 23202 64316 23212 64372
rect 23268 64316 23772 64372
rect 23828 64316 24332 64372
rect 24388 64316 26236 64372
rect 26292 64316 26908 64372
rect 32722 64316 32732 64372
rect 32788 64316 37324 64372
rect 37380 64316 37390 64372
rect 19826 64260 19836 64316
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 20100 64260 20110 64316
rect 11442 64204 11452 64260
rect 11508 64204 11788 64260
rect 11844 64204 14924 64260
rect 14980 64204 16828 64260
rect 16884 64204 17948 64260
rect 18004 64204 18014 64260
rect 31938 64204 31948 64260
rect 32004 64204 37100 64260
rect 37156 64204 37166 64260
rect 23884 64092 25564 64148
rect 25620 64092 25630 64148
rect 28130 64092 28140 64148
rect 28196 64092 28812 64148
rect 28868 64092 29148 64148
rect 29204 64092 29484 64148
rect 29540 64092 29550 64148
rect 32498 64092 32508 64148
rect 32564 64092 36092 64148
rect 36148 64092 38220 64148
rect 38276 64092 38286 64148
rect 23884 64036 23940 64092
rect 14018 63980 14028 64036
rect 14084 63980 19964 64036
rect 20020 63980 20030 64036
rect 20850 63980 20860 64036
rect 20916 63980 21868 64036
rect 21924 63980 21934 64036
rect 23314 63980 23324 64036
rect 23380 63980 23940 64036
rect 23884 63924 23940 63980
rect 24220 63980 24668 64036
rect 24724 63980 27132 64036
rect 27188 63980 27198 64036
rect 27794 63980 27804 64036
rect 27860 63980 29260 64036
rect 29316 63980 29326 64036
rect 32274 63980 32284 64036
rect 32340 63980 32732 64036
rect 32788 63980 32798 64036
rect 33506 63980 33516 64036
rect 33572 63980 34412 64036
rect 34468 63980 34478 64036
rect 24220 63924 24276 63980
rect 14354 63868 14364 63924
rect 14420 63868 15708 63924
rect 15764 63868 15774 63924
rect 16370 63868 16380 63924
rect 16436 63868 17500 63924
rect 17556 63868 17566 63924
rect 21186 63868 21196 63924
rect 21252 63868 23548 63924
rect 23604 63868 23614 63924
rect 23874 63868 23884 63924
rect 23940 63868 23950 63924
rect 24210 63868 24220 63924
rect 24276 63868 24286 63924
rect 28914 63868 28924 63924
rect 28980 63868 29932 63924
rect 29988 63868 29998 63924
rect 32610 63868 32620 63924
rect 32676 63868 33852 63924
rect 33908 63868 33918 63924
rect 35858 63868 35868 63924
rect 35924 63868 37996 63924
rect 38052 63868 38062 63924
rect 4610 63756 4620 63812
rect 4676 63756 6972 63812
rect 7028 63756 7038 63812
rect 11218 63756 11228 63812
rect 11284 63756 11900 63812
rect 11956 63756 11966 63812
rect 23650 63756 23660 63812
rect 23716 63756 24332 63812
rect 24388 63756 24398 63812
rect 26450 63756 26460 63812
rect 26516 63756 27356 63812
rect 27412 63756 27422 63812
rect 6178 63644 6188 63700
rect 6244 63644 8876 63700
rect 8932 63644 8942 63700
rect 26674 63644 26684 63700
rect 26740 63644 28252 63700
rect 28308 63644 28318 63700
rect 29474 63644 29484 63700
rect 29540 63644 30828 63700
rect 30884 63644 30894 63700
rect 4466 63476 4476 63532
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4740 63476 4750 63532
rect 35186 63476 35196 63532
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35460 63476 35470 63532
rect 8418 63308 8428 63364
rect 8484 63308 9212 63364
rect 9268 63308 13468 63364
rect 13524 63308 13534 63364
rect 32162 63308 32172 63364
rect 32228 63308 35196 63364
rect 35252 63308 35262 63364
rect 36642 63308 36652 63364
rect 36708 63308 37548 63364
rect 37604 63308 37614 63364
rect 11890 63196 11900 63252
rect 11956 63196 15148 63252
rect 8978 63084 8988 63140
rect 9044 63084 9660 63140
rect 9716 63084 9726 63140
rect 15092 63028 15148 63196
rect 15698 63084 15708 63140
rect 15764 63084 16044 63140
rect 16100 63084 16604 63140
rect 16660 63084 16670 63140
rect 18946 63084 18956 63140
rect 19012 63084 21420 63140
rect 21476 63084 22876 63140
rect 22932 63084 22942 63140
rect 24546 63084 24556 63140
rect 24612 63084 27020 63140
rect 27076 63084 27804 63140
rect 27860 63084 27870 63140
rect 34962 63084 34972 63140
rect 35028 63084 37548 63140
rect 37604 63084 37614 63140
rect 14466 62972 14476 63028
rect 14532 62972 14542 63028
rect 15092 62972 16156 63028
rect 16212 62972 16222 63028
rect 22194 62972 22204 63028
rect 22260 62972 23100 63028
rect 23156 62972 24332 63028
rect 24388 62972 25788 63028
rect 25844 62972 25854 63028
rect 28466 62972 28476 63028
rect 28532 62972 29260 63028
rect 29316 62972 29596 63028
rect 29652 62972 29662 63028
rect 36418 62972 36428 63028
rect 36484 62972 38220 63028
rect 38276 62972 38286 63028
rect 14476 62804 14532 62972
rect 14802 62860 14812 62916
rect 14868 62860 15036 62916
rect 15092 62860 17052 62916
rect 17108 62860 17118 62916
rect 17266 62860 17276 62916
rect 17332 62860 21420 62916
rect 21476 62860 21486 62916
rect 13906 62748 13916 62804
rect 13972 62748 13982 62804
rect 14476 62748 15484 62804
rect 15540 62748 16716 62804
rect 16772 62748 18172 62804
rect 18228 62748 18238 62804
rect 13916 62692 13972 62748
rect 19826 62692 19836 62748
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 20100 62692 20110 62748
rect 5730 62636 5740 62692
rect 5796 62636 6748 62692
rect 6804 62636 6814 62692
rect 13916 62636 14476 62692
rect 14532 62636 14542 62692
rect 15250 62636 15260 62692
rect 15316 62636 16828 62692
rect 16884 62636 16894 62692
rect 9650 62524 9660 62580
rect 9716 62524 12012 62580
rect 12068 62524 12078 62580
rect 18610 62524 18620 62580
rect 18676 62524 18956 62580
rect 19012 62524 19404 62580
rect 19460 62524 19470 62580
rect 23090 62524 23100 62580
rect 23156 62524 25676 62580
rect 25732 62524 26684 62580
rect 26740 62524 26750 62580
rect 29810 62524 29820 62580
rect 29876 62524 30492 62580
rect 30548 62524 30558 62580
rect 20066 62412 20076 62468
rect 20132 62412 22372 62468
rect 14578 62300 14588 62356
rect 14644 62300 15372 62356
rect 15428 62300 15438 62356
rect 18162 62300 18172 62356
rect 18228 62300 21084 62356
rect 21140 62300 21150 62356
rect 22316 62244 22372 62412
rect 29446 62300 29484 62356
rect 29540 62300 29550 62356
rect 1698 62188 1708 62244
rect 1764 62188 2940 62244
rect 2996 62188 5068 62244
rect 5124 62188 5740 62244
rect 5796 62188 5806 62244
rect 16594 62188 16604 62244
rect 16660 62188 17724 62244
rect 17780 62188 21196 62244
rect 21252 62188 21924 62244
rect 22306 62188 22316 62244
rect 22372 62188 23212 62244
rect 23268 62188 23278 62244
rect 18722 62076 18732 62132
rect 18788 62076 19516 62132
rect 19572 62076 19582 62132
rect 21868 62020 21924 62188
rect 31490 62076 31500 62132
rect 31556 62076 35084 62132
rect 35140 62076 37660 62132
rect 37716 62076 38108 62132
rect 38164 62076 38174 62132
rect 21868 61964 23100 62020
rect 23156 61964 23166 62020
rect 28578 61964 28588 62020
rect 28644 61964 29932 62020
rect 29988 61964 29998 62020
rect 32946 61964 32956 62020
rect 33012 61964 34860 62020
rect 34916 61964 34926 62020
rect 37874 61964 37884 62020
rect 37940 61964 37950 62020
rect 4466 61908 4476 61964
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4740 61908 4750 61964
rect 35186 61908 35196 61964
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35460 61908 35470 61964
rect 29250 61852 29260 61908
rect 29316 61852 30156 61908
rect 30212 61852 30716 61908
rect 30772 61852 30782 61908
rect 37884 61796 37940 61964
rect 32274 61740 32284 61796
rect 32340 61740 33180 61796
rect 33236 61740 36988 61796
rect 37044 61740 37054 61796
rect 37874 61740 37884 61796
rect 37940 61740 37950 61796
rect 3938 61628 3948 61684
rect 4004 61628 4396 61684
rect 4452 61628 4462 61684
rect 5954 61628 5964 61684
rect 6020 61628 6524 61684
rect 6580 61628 7980 61684
rect 8036 61628 8988 61684
rect 9044 61628 9996 61684
rect 10052 61628 10668 61684
rect 10724 61628 10734 61684
rect 21074 61628 21084 61684
rect 21140 61628 21420 61684
rect 21476 61628 21756 61684
rect 21812 61628 21822 61684
rect 31714 61628 31724 61684
rect 31780 61628 33012 61684
rect 33282 61628 33292 61684
rect 33348 61628 33628 61684
rect 33684 61628 33694 61684
rect 37762 61628 37772 61684
rect 37828 61628 38108 61684
rect 38164 61628 38174 61684
rect 15092 61460 15148 61572
rect 15204 61516 18956 61572
rect 19012 61516 19022 61572
rect 28466 61516 28476 61572
rect 28532 61516 30492 61572
rect 30548 61516 30558 61572
rect 31042 61516 31052 61572
rect 31108 61516 32060 61572
rect 32116 61516 32284 61572
rect 32340 61516 32350 61572
rect 13570 61404 13580 61460
rect 13636 61404 14700 61460
rect 14756 61404 15148 61460
rect 29110 61404 29148 61460
rect 29204 61404 29214 61460
rect 32956 61348 33012 61628
rect 33170 61516 33180 61572
rect 33236 61516 33740 61572
rect 33796 61516 33806 61572
rect 33394 61404 33404 61460
rect 33460 61404 35308 61460
rect 35364 61404 35374 61460
rect 4162 61292 4172 61348
rect 4228 61292 4508 61348
rect 4564 61292 4574 61348
rect 7634 61292 7644 61348
rect 7700 61292 9100 61348
rect 9156 61292 9166 61348
rect 17154 61292 17164 61348
rect 17220 61292 17948 61348
rect 18004 61292 18014 61348
rect 19394 61292 19404 61348
rect 19460 61292 20076 61348
rect 20132 61292 20142 61348
rect 22642 61292 22652 61348
rect 22708 61292 22988 61348
rect 23044 61292 23884 61348
rect 23940 61292 23950 61348
rect 32956 61292 37212 61348
rect 37268 61292 37278 61348
rect 31938 61180 31948 61236
rect 32004 61180 33852 61236
rect 33908 61180 33918 61236
rect 19826 61124 19836 61180
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 20100 61124 20110 61180
rect 18946 60956 18956 61012
rect 19012 60956 19516 61012
rect 19572 60956 19582 61012
rect 22530 60956 22540 61012
rect 22596 60956 23100 61012
rect 23156 60956 23660 61012
rect 23716 60956 27692 61012
rect 27748 60956 27758 61012
rect 32274 60956 32284 61012
rect 32340 60956 33292 61012
rect 33348 60956 33358 61012
rect 34738 60956 34748 61012
rect 34804 60956 37548 61012
rect 37604 60956 37614 61012
rect 4274 60844 4284 60900
rect 4340 60844 5740 60900
rect 5796 60844 5806 60900
rect 6850 60844 6860 60900
rect 6916 60844 7532 60900
rect 7588 60844 7598 60900
rect 28242 60844 28252 60900
rect 28308 60844 29148 60900
rect 29204 60844 29484 60900
rect 29540 60844 29550 60900
rect 32834 60844 32844 60900
rect 32900 60844 33516 60900
rect 33572 60844 33582 60900
rect 6178 60732 6188 60788
rect 6244 60732 8092 60788
rect 8148 60732 8158 60788
rect 18946 60732 18956 60788
rect 19012 60732 21196 60788
rect 21252 60732 22764 60788
rect 22820 60732 24220 60788
rect 24276 60732 24668 60788
rect 24724 60732 24734 60788
rect 26852 60732 27468 60788
rect 27524 60732 27916 60788
rect 27972 60732 28364 60788
rect 28420 60732 30828 60788
rect 30884 60732 30894 60788
rect 33618 60732 33628 60788
rect 33684 60732 34188 60788
rect 34244 60732 34254 60788
rect 26852 60676 26908 60732
rect 18722 60620 18732 60676
rect 18788 60620 20748 60676
rect 20804 60620 20814 60676
rect 22418 60620 22428 60676
rect 22484 60620 26908 60676
rect 33842 60620 33852 60676
rect 33908 60620 37716 60676
rect 37660 60564 37716 60620
rect 3378 60508 3388 60564
rect 3444 60508 3724 60564
rect 3780 60508 4508 60564
rect 4564 60508 5292 60564
rect 5348 60508 5358 60564
rect 34850 60508 34860 60564
rect 34916 60508 37100 60564
rect 37156 60508 37166 60564
rect 37650 60508 37660 60564
rect 37716 60508 37726 60564
rect 21074 60396 21084 60452
rect 21140 60396 21644 60452
rect 21700 60396 21710 60452
rect 4466 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4750 60396
rect 35186 60340 35196 60396
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35460 60340 35470 60396
rect 17826 60284 17836 60340
rect 17892 60284 20636 60340
rect 20692 60284 20702 60340
rect 31826 60172 31836 60228
rect 31892 60172 32172 60228
rect 32228 60172 33068 60228
rect 33124 60172 33134 60228
rect 32050 60060 32060 60116
rect 32116 60060 32956 60116
rect 33012 60060 33022 60116
rect 4834 59948 4844 60004
rect 4900 59948 5852 60004
rect 5908 59948 5918 60004
rect 7746 59948 7756 60004
rect 7812 59948 8652 60004
rect 8708 59948 9548 60004
rect 9604 59948 9614 60004
rect 23874 59948 23884 60004
rect 23940 59948 24668 60004
rect 24724 59948 24734 60004
rect 25666 59948 25676 60004
rect 25732 59948 26012 60004
rect 26068 59948 26348 60004
rect 26404 59948 26414 60004
rect 29138 59948 29148 60004
rect 29204 59948 29932 60004
rect 29988 59948 29998 60004
rect 30258 59948 30268 60004
rect 30324 59948 30492 60004
rect 30548 59948 31836 60004
rect 31892 59948 31902 60004
rect 5730 59836 5740 59892
rect 5796 59836 7308 59892
rect 7364 59836 7374 59892
rect 27682 59836 27692 59892
rect 27748 59836 31276 59892
rect 31332 59836 31342 59892
rect 4610 59724 4620 59780
rect 4676 59724 5628 59780
rect 5684 59724 5694 59780
rect 28690 59724 28700 59780
rect 28756 59724 29260 59780
rect 29316 59724 29326 59780
rect 29586 59724 29596 59780
rect 29652 59724 30156 59780
rect 30212 59724 30222 59780
rect 33394 59724 33404 59780
rect 33460 59724 34412 59780
rect 34468 59724 35868 59780
rect 35924 59724 36988 59780
rect 37044 59724 37054 59780
rect 37202 59612 37212 59668
rect 37268 59612 37660 59668
rect 37716 59612 37726 59668
rect 19826 59556 19836 59612
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 20100 59556 20110 59612
rect 18722 59388 18732 59444
rect 18788 59388 21532 59444
rect 21588 59388 21598 59444
rect 29810 59388 29820 59444
rect 29876 59388 31724 59444
rect 31780 59388 32844 59444
rect 32900 59388 34692 59444
rect 34850 59388 34860 59444
rect 34916 59388 37884 59444
rect 37940 59388 37950 59444
rect 34636 59332 34692 59388
rect 14466 59276 14476 59332
rect 14532 59276 15484 59332
rect 15540 59276 15550 59332
rect 17490 59276 17500 59332
rect 17556 59276 19516 59332
rect 19572 59276 19582 59332
rect 32386 59276 32396 59332
rect 32452 59276 33292 59332
rect 33348 59276 33358 59332
rect 34636 59276 35308 59332
rect 35364 59276 35374 59332
rect 36306 59276 36316 59332
rect 36372 59276 37996 59332
rect 38052 59276 38062 59332
rect 1810 59164 1820 59220
rect 1876 59164 3388 59220
rect 10882 59164 10892 59220
rect 10948 59164 13468 59220
rect 13524 59164 13534 59220
rect 16258 59164 16268 59220
rect 16324 59164 17388 59220
rect 17444 59164 18172 59220
rect 18228 59164 18238 59220
rect 25638 59164 25676 59220
rect 25732 59164 25742 59220
rect 29474 59164 29484 59220
rect 29540 59164 30492 59220
rect 30548 59164 30558 59220
rect 35522 59164 35532 59220
rect 35588 59164 36428 59220
rect 36484 59164 36494 59220
rect 3332 59108 3388 59164
rect 3332 59052 3836 59108
rect 3892 59052 5404 59108
rect 5460 59052 7196 59108
rect 7252 59052 8316 59108
rect 8372 59052 8382 59108
rect 14242 59052 14252 59108
rect 14308 59052 14644 59108
rect 14588 58996 14644 59052
rect 15036 59052 16380 59108
rect 16436 59052 16446 59108
rect 19394 59052 19404 59108
rect 19460 59052 21084 59108
rect 21140 59052 21150 59108
rect 23202 59052 23212 59108
rect 23268 59052 23660 59108
rect 23716 59052 26348 59108
rect 26404 59052 26414 59108
rect 15036 58996 15092 59052
rect 7634 58940 7644 58996
rect 7700 58940 7710 58996
rect 14578 58940 14588 58996
rect 14644 58940 14654 58996
rect 15026 58940 15036 58996
rect 15092 58940 15102 58996
rect 34962 58940 34972 58996
rect 35028 58940 36204 58996
rect 36260 58940 36270 58996
rect 4466 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4750 58828
rect 6738 58380 6748 58436
rect 6804 58380 7196 58436
rect 7252 58380 7262 58436
rect 7644 58324 7700 58940
rect 35186 58772 35196 58828
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35460 58772 35470 58828
rect 16034 58716 16044 58772
rect 16100 58716 17612 58772
rect 17668 58716 17678 58772
rect 32498 58716 32508 58772
rect 32564 58716 33852 58772
rect 33908 58716 33918 58772
rect 13794 58604 13804 58660
rect 13860 58604 15596 58660
rect 15652 58604 16716 58660
rect 16772 58604 17836 58660
rect 17892 58604 17902 58660
rect 18610 58604 18620 58660
rect 18676 58604 19180 58660
rect 19236 58604 19246 58660
rect 32946 58604 32956 58660
rect 33012 58604 35868 58660
rect 35924 58604 37212 58660
rect 37268 58604 37772 58660
rect 37828 58604 37838 58660
rect 13458 58492 13468 58548
rect 13524 58492 20300 58548
rect 20356 58492 20366 58548
rect 30258 58492 30268 58548
rect 30324 58492 30604 58548
rect 30660 58492 30670 58548
rect 32722 58492 32732 58548
rect 32788 58492 33516 58548
rect 33572 58492 33964 58548
rect 34020 58492 34030 58548
rect 14018 58380 14028 58436
rect 14084 58380 15036 58436
rect 15092 58380 15102 58436
rect 21410 58380 21420 58436
rect 21476 58380 24668 58436
rect 24724 58380 24892 58436
rect 24948 58380 24958 58436
rect 5058 58268 5068 58324
rect 5124 58268 6188 58324
rect 6244 58268 7308 58324
rect 7364 58268 7700 58324
rect 14028 58212 14084 58380
rect 39600 58324 40000 58352
rect 27682 58268 27692 58324
rect 27748 58268 28252 58324
rect 28308 58268 29820 58324
rect 29876 58268 31276 58324
rect 31332 58268 31342 58324
rect 38210 58268 38220 58324
rect 38276 58268 40000 58324
rect 39600 58240 40000 58268
rect 4610 58156 4620 58212
rect 4676 58156 5740 58212
rect 5796 58156 6972 58212
rect 7028 58156 7868 58212
rect 7924 58156 7934 58212
rect 8418 58156 8428 58212
rect 8484 58156 9772 58212
rect 9828 58156 11676 58212
rect 11732 58156 14084 58212
rect 16818 58156 16828 58212
rect 16884 58156 17612 58212
rect 17668 58156 17678 58212
rect 28018 58156 28028 58212
rect 28084 58156 29484 58212
rect 29540 58156 31836 58212
rect 31892 58156 31902 58212
rect 16940 57988 16996 58156
rect 17266 58044 17276 58100
rect 17332 58044 17836 58100
rect 17892 58044 17902 58100
rect 19826 57988 19836 58044
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20100 57988 20110 58044
rect 16930 57932 16940 57988
rect 16996 57932 17006 57988
rect 14578 57820 14588 57876
rect 14644 57820 16044 57876
rect 16100 57820 16110 57876
rect 16790 57708 16828 57764
rect 16884 57708 17388 57764
rect 17444 57708 17454 57764
rect 20178 57708 20188 57764
rect 20244 57708 23268 57764
rect 23212 57652 23268 57708
rect 6962 57596 6972 57652
rect 7028 57596 7532 57652
rect 7588 57596 8204 57652
rect 8260 57596 8270 57652
rect 12450 57596 12460 57652
rect 12516 57596 13692 57652
rect 13748 57596 13758 57652
rect 19954 57596 19964 57652
rect 20020 57596 20636 57652
rect 20692 57596 22316 57652
rect 22372 57596 22382 57652
rect 23202 57596 23212 57652
rect 23268 57596 28028 57652
rect 28084 57596 28094 57652
rect 21858 57484 21868 57540
rect 21924 57484 22764 57540
rect 22820 57484 22830 57540
rect 34290 57484 34300 57540
rect 34356 57484 35084 57540
rect 35140 57484 35150 57540
rect 18498 57372 18508 57428
rect 18564 57372 19628 57428
rect 19684 57372 19694 57428
rect 29698 57260 29708 57316
rect 29764 57260 30380 57316
rect 30436 57260 30940 57316
rect 30996 57260 31006 57316
rect 4466 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4750 57260
rect 35186 57204 35196 57260
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35460 57204 35470 57260
rect 5842 57148 5852 57204
rect 5908 57148 6188 57204
rect 6244 57148 6254 57204
rect 18274 57148 18284 57204
rect 18340 57148 19404 57204
rect 19460 57148 19470 57204
rect 18806 57036 18844 57092
rect 18900 57036 18910 57092
rect 19254 57036 19292 57092
rect 19348 57036 19358 57092
rect 22082 57036 22092 57092
rect 22148 57036 23548 57092
rect 23604 57036 23614 57092
rect 24882 57036 24892 57092
rect 24948 57036 26684 57092
rect 26740 57036 28140 57092
rect 28196 57036 28206 57092
rect 17938 56924 17948 56980
rect 18004 56924 18396 56980
rect 18452 56924 18462 56980
rect 24546 56924 24556 56980
rect 24612 56924 27468 56980
rect 27524 56924 27534 56980
rect 30594 56924 30604 56980
rect 30660 56924 31948 56980
rect 32004 56924 32014 56980
rect 18834 56812 18844 56868
rect 18900 56812 19180 56868
rect 19236 56812 19246 56868
rect 24658 56812 24668 56868
rect 24724 56812 29148 56868
rect 29204 56812 29214 56868
rect 13010 56588 13020 56644
rect 13076 56588 14364 56644
rect 14420 56588 14430 56644
rect 8194 56476 8204 56532
rect 8260 56476 16604 56532
rect 16660 56476 17164 56532
rect 17220 56476 17230 56532
rect 18498 56476 18508 56532
rect 18564 56476 18574 56532
rect 18050 56364 18060 56420
rect 18116 56364 18126 56420
rect 18060 56196 18116 56364
rect 18508 56308 18564 56476
rect 19826 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20110 56476
rect 18508 56252 19740 56308
rect 19796 56252 19806 56308
rect 24882 56252 24892 56308
rect 24948 56252 25340 56308
rect 25396 56252 25406 56308
rect 28130 56252 28140 56308
rect 28196 56252 30940 56308
rect 30996 56252 31836 56308
rect 31892 56252 31902 56308
rect 18060 56140 18508 56196
rect 18564 56140 18574 56196
rect 11554 56028 11564 56084
rect 11620 56028 12236 56084
rect 12292 56028 12302 56084
rect 3378 55916 3388 55972
rect 3444 55916 3948 55972
rect 4004 55916 4014 55972
rect 17938 55916 17948 55972
rect 18004 55916 18732 55972
rect 18788 55916 18798 55972
rect 4466 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4750 55692
rect 35186 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35470 55692
rect 3042 55356 3052 55412
rect 3108 55356 3612 55412
rect 3668 55356 3678 55412
rect 8530 55356 8540 55412
rect 8596 55356 10892 55412
rect 10948 55356 10958 55412
rect 11890 55356 11900 55412
rect 11956 55356 14812 55412
rect 14868 55356 14878 55412
rect 19730 55356 19740 55412
rect 19796 55356 20860 55412
rect 20916 55356 22092 55412
rect 22148 55356 22158 55412
rect 22530 55356 22540 55412
rect 22596 55356 23324 55412
rect 23380 55356 23390 55412
rect 31154 55356 31164 55412
rect 31220 55356 32284 55412
rect 32340 55356 32350 55412
rect 14018 55244 14028 55300
rect 14084 55244 27916 55300
rect 27972 55244 28476 55300
rect 28532 55244 28542 55300
rect 22082 55132 22092 55188
rect 22148 55132 24556 55188
rect 24612 55132 24622 55188
rect 34850 55132 34860 55188
rect 34916 55132 35420 55188
rect 35476 55132 36428 55188
rect 36484 55132 36494 55188
rect 6178 55020 6188 55076
rect 6244 55020 9324 55076
rect 9380 55020 9390 55076
rect 16706 55020 16716 55076
rect 16772 55020 21420 55076
rect 21476 55020 21868 55076
rect 21924 55020 21934 55076
rect 24210 55020 24220 55076
rect 24276 55020 25004 55076
rect 25060 55020 25070 55076
rect 0 54964 400 54992
rect 0 54908 3500 54964
rect 3556 54908 3566 54964
rect 0 54880 400 54908
rect 19826 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20110 54908
rect 11414 54796 11452 54852
rect 11508 54796 11518 54852
rect 3154 54684 3164 54740
rect 3220 54684 3612 54740
rect 3668 54684 3678 54740
rect 11666 54684 11676 54740
rect 11732 54684 12684 54740
rect 12740 54684 12750 54740
rect 28354 54684 28364 54740
rect 28420 54684 30044 54740
rect 30100 54684 31276 54740
rect 31332 54684 31342 54740
rect 6850 54572 6860 54628
rect 6916 54572 9548 54628
rect 9604 54572 9614 54628
rect 27906 54572 27916 54628
rect 27972 54572 29372 54628
rect 29428 54572 29438 54628
rect 8418 54460 8428 54516
rect 8484 54460 8988 54516
rect 9044 54460 11228 54516
rect 11284 54460 11294 54516
rect 21522 54460 21532 54516
rect 21588 54460 27076 54516
rect 28466 54460 28476 54516
rect 28532 54460 28812 54516
rect 28868 54460 29148 54516
rect 29204 54460 29214 54516
rect 3938 54348 3948 54404
rect 4004 54348 4620 54404
rect 4676 54348 11900 54404
rect 11956 54348 11966 54404
rect 23426 54348 23436 54404
rect 23492 54348 24444 54404
rect 24500 54348 24510 54404
rect 27020 54292 27076 54460
rect 30146 54348 30156 54404
rect 30212 54348 32060 54404
rect 32116 54348 32126 54404
rect 23090 54236 23100 54292
rect 23156 54236 23548 54292
rect 23604 54236 24220 54292
rect 24276 54236 24286 54292
rect 27010 54236 27020 54292
rect 27076 54236 27692 54292
rect 27748 54236 28364 54292
rect 28420 54236 28430 54292
rect 4466 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4750 54124
rect 35186 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35470 54124
rect 3910 54012 3948 54068
rect 4004 54012 4014 54068
rect 12338 54012 12348 54068
rect 12404 54012 14812 54068
rect 14868 54012 15596 54068
rect 15652 54012 15662 54068
rect 10882 53900 10892 53956
rect 10948 53900 12236 53956
rect 12292 53900 15148 53956
rect 18498 53900 18508 53956
rect 18564 53900 19180 53956
rect 19236 53900 20748 53956
rect 20804 53900 21644 53956
rect 21700 53900 26012 53956
rect 26068 53900 26078 53956
rect 26786 53900 26796 53956
rect 26852 53900 27356 53956
rect 27412 53900 27422 53956
rect 15092 53844 15148 53900
rect 4834 53788 4844 53844
rect 4900 53788 5068 53844
rect 5124 53788 6188 53844
rect 6244 53788 6254 53844
rect 10770 53788 10780 53844
rect 10836 53788 13468 53844
rect 13524 53788 13534 53844
rect 15092 53788 17052 53844
rect 17108 53788 17118 53844
rect 28466 53788 28476 53844
rect 28532 53788 29372 53844
rect 29428 53788 29438 53844
rect 7298 53676 7308 53732
rect 7364 53676 8204 53732
rect 8260 53676 8652 53732
rect 8708 53676 8988 53732
rect 9044 53676 9054 53732
rect 11778 53676 11788 53732
rect 11844 53676 12908 53732
rect 12964 53676 12974 53732
rect 15092 53676 15820 53732
rect 15876 53676 16828 53732
rect 16884 53676 16894 53732
rect 20402 53676 20412 53732
rect 20468 53676 20636 53732
rect 20692 53676 20702 53732
rect 28914 53676 28924 53732
rect 28980 53676 29484 53732
rect 29540 53676 29550 53732
rect 30482 53676 30492 53732
rect 30548 53676 31836 53732
rect 31892 53676 32396 53732
rect 32452 53676 33852 53732
rect 33908 53676 33918 53732
rect 3714 53564 3724 53620
rect 3780 53564 6300 53620
rect 6356 53564 6366 53620
rect 7970 53564 7980 53620
rect 8036 53564 8428 53620
rect 8484 53564 9660 53620
rect 9716 53564 9726 53620
rect 12338 53564 12348 53620
rect 12404 53564 13804 53620
rect 13860 53564 13870 53620
rect 15092 53508 15148 53676
rect 20290 53564 20300 53620
rect 20356 53564 21868 53620
rect 21924 53564 21934 53620
rect 10098 53452 10108 53508
rect 10164 53452 11564 53508
rect 11620 53452 14252 53508
rect 14308 53452 15148 53508
rect 17826 53452 17836 53508
rect 17892 53452 18172 53508
rect 18228 53452 21980 53508
rect 22036 53452 22046 53508
rect 22306 53452 22316 53508
rect 22372 53452 23436 53508
rect 23492 53452 35364 53508
rect 25890 53340 25900 53396
rect 25956 53340 26796 53396
rect 26852 53340 26862 53396
rect 19826 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20110 53340
rect 4918 53228 4956 53284
rect 5012 53228 5022 53284
rect 4610 53116 4620 53172
rect 4676 53116 5404 53172
rect 5460 53116 5470 53172
rect 6626 53116 6636 53172
rect 6692 53116 7308 53172
rect 7364 53116 7980 53172
rect 8036 53116 8046 53172
rect 11442 53116 11452 53172
rect 11508 53116 12012 53172
rect 12068 53116 12078 53172
rect 15250 53116 15260 53172
rect 15316 53116 16268 53172
rect 16324 53116 16334 53172
rect 21410 53116 21420 53172
rect 21476 53116 23660 53172
rect 23716 53116 23726 53172
rect 33842 53116 33852 53172
rect 33908 53116 34972 53172
rect 35028 53116 35038 53172
rect 4050 53004 4060 53060
rect 4116 53004 4844 53060
rect 4900 53004 4910 53060
rect 16594 53004 16604 53060
rect 16660 53004 18844 53060
rect 18900 53004 18910 53060
rect 19394 53004 19404 53060
rect 19460 53004 20524 53060
rect 20580 53004 20590 53060
rect 5170 52892 5180 52948
rect 5236 52892 6076 52948
rect 6132 52892 6142 52948
rect 15092 52892 16044 52948
rect 16100 52892 16110 52948
rect 18050 52892 18060 52948
rect 18116 52892 20636 52948
rect 20692 52892 20702 52948
rect 21298 52892 21308 52948
rect 21364 52892 22764 52948
rect 22820 52892 22830 52948
rect 29148 52892 32284 52948
rect 32340 52892 32350 52948
rect 15092 52836 15148 52892
rect 29148 52836 29204 52892
rect 35308 52836 35364 53452
rect 6850 52780 6860 52836
rect 6916 52780 13020 52836
rect 13076 52780 15148 52836
rect 18274 52780 18284 52836
rect 18340 52780 18956 52836
rect 19012 52780 19022 52836
rect 20738 52780 20748 52836
rect 20804 52780 21644 52836
rect 21700 52780 21710 52836
rect 28018 52780 28028 52836
rect 28084 52780 28588 52836
rect 28644 52780 29148 52836
rect 29204 52780 29214 52836
rect 31462 52780 31500 52836
rect 31556 52780 31566 52836
rect 35298 52780 35308 52836
rect 35364 52780 35374 52836
rect 3490 52668 3500 52724
rect 3556 52668 7644 52724
rect 7700 52668 7710 52724
rect 16258 52668 16268 52724
rect 16324 52668 17388 52724
rect 17444 52668 17454 52724
rect 17714 52668 17724 52724
rect 17780 52668 21532 52724
rect 21588 52668 23884 52724
rect 23940 52668 23950 52724
rect 31378 52668 31388 52724
rect 31444 52668 33404 52724
rect 33460 52668 34076 52724
rect 34132 52668 35644 52724
rect 35700 52668 35710 52724
rect 7522 52556 7532 52612
rect 7588 52556 8204 52612
rect 8260 52556 8270 52612
rect 16370 52556 16380 52612
rect 16436 52556 17500 52612
rect 17556 52556 18844 52612
rect 18900 52556 23772 52612
rect 23828 52556 23838 52612
rect 4466 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4750 52556
rect 35186 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35470 52556
rect 7298 52444 7308 52500
rect 7364 52444 8316 52500
rect 8372 52444 8382 52500
rect 19954 52444 19964 52500
rect 20020 52444 23324 52500
rect 23380 52444 23436 52500
rect 23492 52444 23502 52500
rect 15092 52332 22316 52388
rect 22372 52332 22382 52388
rect 15092 52276 15148 52332
rect 11778 52220 11788 52276
rect 11844 52220 12908 52276
rect 12964 52220 15148 52276
rect 16818 52220 16828 52276
rect 16884 52220 17164 52276
rect 17220 52220 18060 52276
rect 18116 52220 18126 52276
rect 21410 52220 21420 52276
rect 21476 52220 22092 52276
rect 22148 52220 22158 52276
rect 2034 52108 2044 52164
rect 2100 52108 5068 52164
rect 5124 52108 5134 52164
rect 13010 52108 13020 52164
rect 13076 52108 15596 52164
rect 15652 52108 15662 52164
rect 20066 52108 20076 52164
rect 20132 52108 20860 52164
rect 20916 52108 21084 52164
rect 21140 52108 21150 52164
rect 21298 52108 21308 52164
rect 21364 52108 23996 52164
rect 24052 52108 24668 52164
rect 24724 52108 24734 52164
rect 35634 52108 35644 52164
rect 35700 52108 36316 52164
rect 36372 52108 36382 52164
rect 2706 51996 2716 52052
rect 2772 51996 3836 52052
rect 3892 51996 3902 52052
rect 4918 51996 4956 52052
rect 5012 51996 5022 52052
rect 5618 51996 5628 52052
rect 5684 51996 10220 52052
rect 10276 51996 10286 52052
rect 16790 51996 16828 52052
rect 16884 51996 17948 52052
rect 18004 51996 19964 52052
rect 20020 51996 20030 52052
rect 20290 51996 20300 52052
rect 20356 51996 21756 52052
rect 21812 51996 25340 52052
rect 25396 51996 25406 52052
rect 35746 51996 35756 52052
rect 35812 51996 37548 52052
rect 37604 51996 38108 52052
rect 38164 51996 38174 52052
rect 18834 51884 18844 51940
rect 18900 51884 19292 51940
rect 19348 51884 19358 51940
rect 22194 51884 22204 51940
rect 22260 51884 23436 51940
rect 23492 51884 25116 51940
rect 25172 51884 25182 51940
rect 19826 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20110 51772
rect 15810 51660 15820 51716
rect 15876 51660 15886 51716
rect 17826 51660 17836 51716
rect 17892 51660 19180 51716
rect 19236 51660 19246 51716
rect 19590 51660 19628 51716
rect 19684 51660 19694 51716
rect 15820 51492 15876 51660
rect 16594 51548 16604 51604
rect 16660 51548 18172 51604
rect 18228 51548 19516 51604
rect 19572 51548 19582 51604
rect 15820 51436 18620 51492
rect 18676 51436 18686 51492
rect 20514 51436 20524 51492
rect 20580 51436 23548 51492
rect 23604 51436 23614 51492
rect 4162 51324 4172 51380
rect 4228 51324 6300 51380
rect 6356 51324 6366 51380
rect 16370 51324 16380 51380
rect 16436 51324 18396 51380
rect 18452 51324 19404 51380
rect 19460 51324 19470 51380
rect 22418 51324 22428 51380
rect 22484 51324 22988 51380
rect 23044 51324 23054 51380
rect 27682 51324 27692 51380
rect 27748 51324 30380 51380
rect 30436 51324 31164 51380
rect 31220 51324 31230 51380
rect 9314 51212 9324 51268
rect 9380 51212 10780 51268
rect 10836 51212 10846 51268
rect 12002 51212 12012 51268
rect 12068 51212 26124 51268
rect 26180 51212 26190 51268
rect 19170 51100 19180 51156
rect 19236 51100 28476 51156
rect 28532 51100 28542 51156
rect 16706 50988 16716 51044
rect 16772 50988 18284 51044
rect 18340 50988 18350 51044
rect 18610 50988 18620 51044
rect 18676 50988 22596 51044
rect 4466 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4750 50988
rect 22540 50932 22596 50988
rect 35186 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35470 50988
rect 16258 50876 16268 50932
rect 16324 50876 21532 50932
rect 21588 50876 21598 50932
rect 22530 50876 22540 50932
rect 22596 50876 30380 50932
rect 30436 50876 30446 50932
rect 18610 50764 18620 50820
rect 18676 50764 22204 50820
rect 22260 50764 22270 50820
rect 9426 50652 9436 50708
rect 9492 50652 21980 50708
rect 22036 50652 22046 50708
rect 26114 50652 26124 50708
rect 26180 50652 27692 50708
rect 27748 50652 27758 50708
rect 17714 50540 17724 50596
rect 17780 50540 20636 50596
rect 20692 50540 21756 50596
rect 21812 50540 21822 50596
rect 23986 50540 23996 50596
rect 24052 50540 27244 50596
rect 27300 50540 28028 50596
rect 28084 50540 28094 50596
rect 15362 50428 15372 50484
rect 15428 50428 17612 50484
rect 17668 50428 17678 50484
rect 19506 50428 19516 50484
rect 19572 50428 20076 50484
rect 20132 50428 20142 50484
rect 23426 50428 23436 50484
rect 23492 50428 24612 50484
rect 24546 50372 24556 50428
rect 24612 50372 24622 50428
rect 15922 50316 15932 50372
rect 15988 50316 18508 50372
rect 18564 50316 18574 50372
rect 34738 50316 34748 50372
rect 34804 50316 37884 50372
rect 37940 50316 37950 50372
rect 19826 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20110 50204
rect 20402 50092 20412 50148
rect 20468 50092 23100 50148
rect 23156 50092 23166 50148
rect 5058 49980 5068 50036
rect 5124 49980 5964 50036
rect 6020 49980 6030 50036
rect 10098 49980 10108 50036
rect 10164 49980 11116 50036
rect 11172 49980 11676 50036
rect 11732 49980 17052 50036
rect 17108 49980 17118 50036
rect 19394 49980 19404 50036
rect 19460 49980 20860 50036
rect 20916 49980 23380 50036
rect 23324 49924 23380 49980
rect 17602 49868 17612 49924
rect 17668 49868 18620 49924
rect 18676 49868 20748 49924
rect 20804 49868 20814 49924
rect 23314 49868 23324 49924
rect 23380 49868 23548 49924
rect 23604 49868 23614 49924
rect 26908 49868 27244 49924
rect 27300 49868 27310 49924
rect 26908 49812 26964 49868
rect 10434 49756 10444 49812
rect 10500 49756 11004 49812
rect 11060 49756 11070 49812
rect 11666 49756 11676 49812
rect 11732 49756 14364 49812
rect 14420 49756 14924 49812
rect 14980 49756 14990 49812
rect 17826 49756 17836 49812
rect 17892 49756 20188 49812
rect 20244 49756 20254 49812
rect 24210 49756 24220 49812
rect 24276 49756 25228 49812
rect 25284 49756 25294 49812
rect 26898 49756 26908 49812
rect 26964 49756 26974 49812
rect 34962 49756 34972 49812
rect 35028 49756 35644 49812
rect 35700 49756 35710 49812
rect 12338 49644 12348 49700
rect 12404 49644 13580 49700
rect 13636 49644 13646 49700
rect 21074 49644 21084 49700
rect 21140 49644 22988 49700
rect 23044 49644 23054 49700
rect 4722 49532 4732 49588
rect 4788 49532 4900 49588
rect 15250 49532 15260 49588
rect 15316 49532 16828 49588
rect 16884 49532 17500 49588
rect 17556 49532 20524 49588
rect 20580 49532 20590 49588
rect 4844 49476 4900 49532
rect 26908 49476 26964 49756
rect 27346 49644 27356 49700
rect 27412 49644 27692 49700
rect 27748 49644 27758 49700
rect 4844 49420 4956 49476
rect 5012 49420 5022 49476
rect 7634 49420 7644 49476
rect 7700 49420 17836 49476
rect 17892 49420 17902 49476
rect 26908 49420 27692 49476
rect 27748 49420 28476 49476
rect 28532 49420 29708 49476
rect 29764 49420 30268 49476
rect 30324 49420 30334 49476
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 10322 49308 10332 49364
rect 10388 49308 15596 49364
rect 15652 49308 15662 49364
rect 16482 49308 16492 49364
rect 16548 49308 21420 49364
rect 21476 49308 21486 49364
rect 24658 49308 24668 49364
rect 24724 49308 25340 49364
rect 25396 49308 25406 49364
rect 25554 49308 25564 49364
rect 25620 49308 27020 49364
rect 27076 49308 27086 49364
rect 30156 49308 30716 49364
rect 30772 49308 30782 49364
rect 30156 49252 30212 49308
rect 7970 49196 7980 49252
rect 8036 49196 8876 49252
rect 8932 49196 8942 49252
rect 12450 49196 12460 49252
rect 12516 49196 13468 49252
rect 13524 49196 13534 49252
rect 14466 49196 14476 49252
rect 14532 49196 14812 49252
rect 14868 49196 14878 49252
rect 19394 49196 19404 49252
rect 19460 49196 30212 49252
rect 30370 49196 30380 49252
rect 30436 49196 31164 49252
rect 31220 49196 33740 49252
rect 33796 49196 33806 49252
rect 16034 49084 16044 49140
rect 16100 49084 24892 49140
rect 24948 49084 25900 49140
rect 25956 49084 25966 49140
rect 10098 48972 10108 49028
rect 10164 48972 11228 49028
rect 11284 48972 11294 49028
rect 13794 48972 13804 49028
rect 13860 48972 14700 49028
rect 14756 48972 15932 49028
rect 15988 48972 15998 49028
rect 18610 48972 18620 49028
rect 18676 48972 22316 49028
rect 22372 48972 22382 49028
rect 30156 48916 30212 49196
rect 13010 48860 13020 48916
rect 13076 48860 14140 48916
rect 14196 48860 14206 48916
rect 23090 48860 23100 48916
rect 23156 48860 24108 48916
rect 24164 48860 24174 48916
rect 30156 48860 30604 48916
rect 30660 48860 34188 48916
rect 34244 48860 34254 48916
rect 34188 48804 34244 48860
rect 11890 48748 11900 48804
rect 11956 48748 12908 48804
rect 12964 48748 14252 48804
rect 14308 48748 14318 48804
rect 14914 48748 14924 48804
rect 14980 48748 15820 48804
rect 15876 48748 15886 48804
rect 21634 48748 21644 48804
rect 21700 48748 22652 48804
rect 22708 48748 25228 48804
rect 25284 48748 28252 48804
rect 28308 48748 28318 48804
rect 28802 48748 28812 48804
rect 28868 48748 29260 48804
rect 29316 48748 29326 48804
rect 34188 48748 34860 48804
rect 34916 48748 35196 48804
rect 35252 48748 35262 48804
rect 6850 48636 6860 48692
rect 6916 48636 8316 48692
rect 8372 48636 10444 48692
rect 10500 48636 10510 48692
rect 11414 48636 11452 48692
rect 11508 48636 11518 48692
rect 15092 48636 17052 48692
rect 17108 48636 17118 48692
rect 22754 48636 22764 48692
rect 22820 48636 23436 48692
rect 23492 48636 23660 48692
rect 23716 48636 23726 48692
rect 25778 48636 25788 48692
rect 25844 48636 27692 48692
rect 27748 48636 27758 48692
rect 34748 48636 35532 48692
rect 35588 48636 36204 48692
rect 36260 48636 36270 48692
rect 15092 48580 15148 48636
rect 19826 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20110 48636
rect 25788 48580 25844 48636
rect 9650 48524 9660 48580
rect 9716 48524 10220 48580
rect 10276 48524 15148 48580
rect 16258 48524 16268 48580
rect 16324 48524 19404 48580
rect 19460 48524 19470 48580
rect 21970 48524 21980 48580
rect 22036 48524 22316 48580
rect 22372 48524 24668 48580
rect 24724 48524 25844 48580
rect 26450 48524 26460 48580
rect 26516 48524 26796 48580
rect 26852 48524 26862 48580
rect 34748 48468 34804 48636
rect 13906 48412 13916 48468
rect 13972 48412 17388 48468
rect 17444 48412 17454 48468
rect 22978 48412 22988 48468
rect 23044 48412 23324 48468
rect 23380 48412 28028 48468
rect 28084 48412 28094 48468
rect 28578 48412 28588 48468
rect 28644 48412 29372 48468
rect 29428 48412 29438 48468
rect 33842 48412 33852 48468
rect 33908 48412 34748 48468
rect 34804 48412 34814 48468
rect 2930 48300 2940 48356
rect 2996 48300 3724 48356
rect 3780 48300 3790 48356
rect 15810 48300 15820 48356
rect 15876 48300 16492 48356
rect 16548 48300 16558 48356
rect 23650 48300 23660 48356
rect 23716 48300 31724 48356
rect 31780 48300 31790 48356
rect 14690 48188 14700 48244
rect 14756 48188 15372 48244
rect 15428 48188 15438 48244
rect 20514 48188 20524 48244
rect 20580 48188 21868 48244
rect 21924 48188 21934 48244
rect 22082 48188 22092 48244
rect 22148 48188 22652 48244
rect 22708 48188 22718 48244
rect 23874 48188 23884 48244
rect 23940 48188 27468 48244
rect 27524 48188 27534 48244
rect 5282 48076 5292 48132
rect 5348 48076 8876 48132
rect 8932 48076 9996 48132
rect 10052 48076 10062 48132
rect 10658 48076 10668 48132
rect 10724 48076 12348 48132
rect 12404 48076 13020 48132
rect 13076 48076 13086 48132
rect 23426 48076 23436 48132
rect 23492 48076 26124 48132
rect 26180 48076 26796 48132
rect 26852 48076 26862 48132
rect 30482 48076 30492 48132
rect 30548 48076 31388 48132
rect 31444 48076 32284 48132
rect 32340 48076 32350 48132
rect 8754 47964 8764 48020
rect 8820 47964 11676 48020
rect 11732 47964 12796 48020
rect 12852 47964 12862 48020
rect 12796 47908 12852 47964
rect 12796 47852 21644 47908
rect 21700 47852 26460 47908
rect 26516 47852 26526 47908
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 5058 47740 5068 47796
rect 5124 47740 5134 47796
rect 14802 47740 14812 47796
rect 14868 47740 15820 47796
rect 15876 47740 15886 47796
rect 5068 47236 5124 47740
rect 35522 47628 35532 47684
rect 35588 47628 36204 47684
rect 36260 47628 36270 47684
rect 13682 47516 13692 47572
rect 13748 47516 15596 47572
rect 15652 47516 15662 47572
rect 34066 47516 34076 47572
rect 34132 47516 34748 47572
rect 34804 47516 37548 47572
rect 37604 47516 37614 47572
rect 9426 47404 9436 47460
rect 9492 47404 10108 47460
rect 10164 47404 11788 47460
rect 28466 47404 28476 47460
rect 28532 47404 30828 47460
rect 30884 47404 31052 47460
rect 31108 47404 31836 47460
rect 31892 47404 31902 47460
rect 5282 47292 5292 47348
rect 5348 47292 6076 47348
rect 6132 47292 6142 47348
rect 11732 47236 11788 47404
rect 13122 47292 13132 47348
rect 13188 47292 15036 47348
rect 15092 47292 15102 47348
rect 15474 47292 15484 47348
rect 15540 47292 23660 47348
rect 23716 47292 23726 47348
rect 5068 47180 5740 47236
rect 5796 47180 7756 47236
rect 7812 47180 8316 47236
rect 8372 47180 8382 47236
rect 11732 47180 13580 47236
rect 13636 47180 13646 47236
rect 14354 47180 14364 47236
rect 14420 47180 15708 47236
rect 15764 47180 15774 47236
rect 16258 47180 16268 47236
rect 16324 47180 17164 47236
rect 17220 47180 19068 47236
rect 19124 47180 19134 47236
rect 20066 47180 20076 47236
rect 20132 47180 26908 47236
rect 26964 47180 26974 47236
rect 2258 47068 2268 47124
rect 2324 47068 5292 47124
rect 5348 47068 5358 47124
rect 20850 47068 20860 47124
rect 20916 47068 21532 47124
rect 21588 47068 22204 47124
rect 22260 47068 24276 47124
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 24220 47012 24276 47068
rect 28588 47012 28644 47404
rect 31490 47292 31500 47348
rect 31556 47292 32620 47348
rect 32676 47292 32686 47348
rect 36194 47292 36204 47348
rect 36260 47292 36988 47348
rect 37044 47292 37054 47348
rect 30930 47180 30940 47236
rect 30996 47180 31500 47236
rect 31556 47180 31566 47236
rect 24210 46956 24220 47012
rect 24276 46956 27244 47012
rect 27300 46956 27310 47012
rect 28578 46956 28588 47012
rect 28644 46956 28654 47012
rect 32050 46956 32060 47012
rect 32116 46956 33180 47012
rect 33236 46956 37212 47012
rect 37268 46956 37996 47012
rect 38052 46956 38062 47012
rect 11554 46844 11564 46900
rect 11620 46844 25228 46900
rect 25284 46844 25956 46900
rect 27906 46844 27916 46900
rect 27972 46844 28010 46900
rect 33394 46844 33404 46900
rect 33460 46844 35084 46900
rect 35140 46844 35150 46900
rect 18722 46732 18732 46788
rect 18788 46732 19964 46788
rect 20020 46732 20030 46788
rect 21074 46732 21084 46788
rect 21140 46732 23324 46788
rect 23380 46732 23660 46788
rect 23716 46732 24164 46788
rect 24322 46732 24332 46788
rect 24388 46732 25340 46788
rect 25396 46732 25406 46788
rect 24108 46676 24164 46732
rect 25900 46676 25956 46844
rect 26646 46732 26684 46788
rect 26740 46732 26750 46788
rect 36418 46732 36428 46788
rect 36484 46732 37436 46788
rect 37492 46732 37502 46788
rect 19506 46620 19516 46676
rect 19572 46620 21756 46676
rect 21812 46620 22092 46676
rect 22148 46620 22158 46676
rect 24098 46620 24108 46676
rect 24164 46620 24668 46676
rect 24724 46620 25844 46676
rect 25900 46620 28588 46676
rect 28644 46620 28654 46676
rect 25788 46564 25844 46620
rect 15586 46508 15596 46564
rect 15652 46508 16268 46564
rect 16324 46508 16334 46564
rect 18386 46508 18396 46564
rect 18452 46508 20860 46564
rect 20916 46508 20926 46564
rect 25554 46508 25564 46564
rect 25620 46508 25658 46564
rect 25788 46508 28140 46564
rect 28196 46508 28812 46564
rect 28868 46508 28878 46564
rect 18274 46396 18284 46452
rect 18340 46396 25732 46452
rect 26562 46396 26572 46452
rect 26628 46396 26908 46452
rect 26964 46396 28364 46452
rect 28420 46396 28430 46452
rect 29922 46396 29932 46452
rect 29988 46396 30604 46452
rect 30660 46396 31164 46452
rect 31220 46396 31230 46452
rect 35298 46396 35308 46452
rect 35364 46396 36988 46452
rect 37044 46396 37054 46452
rect 15922 46284 15932 46340
rect 15988 46284 18172 46340
rect 18228 46284 19404 46340
rect 19460 46284 19470 46340
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 25676 46228 25732 46396
rect 26198 46284 26236 46340
rect 26292 46284 26302 46340
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 6178 46172 6188 46228
rect 6244 46172 17500 46228
rect 17556 46172 23548 46228
rect 25676 46172 29148 46228
rect 29204 46172 30492 46228
rect 30548 46172 30558 46228
rect 23492 46116 23548 46172
rect 23492 46060 25452 46116
rect 25508 46060 29036 46116
rect 29092 46060 29102 46116
rect 30258 46060 30268 46116
rect 30324 46060 31164 46116
rect 31220 46060 31230 46116
rect 16370 45948 16380 46004
rect 16436 45948 19068 46004
rect 19124 45948 19134 46004
rect 23650 45948 23660 46004
rect 23716 45948 25564 46004
rect 25620 45948 25630 46004
rect 25778 45948 25788 46004
rect 25844 45948 27916 46004
rect 27972 45948 27982 46004
rect 28466 45948 28476 46004
rect 28532 45948 30604 46004
rect 30660 45948 30670 46004
rect 12898 45836 12908 45892
rect 12964 45836 13804 45892
rect 13860 45836 13870 45892
rect 16482 45836 16492 45892
rect 16548 45836 20524 45892
rect 20580 45836 21980 45892
rect 22036 45836 22046 45892
rect 22838 45836 22876 45892
rect 22932 45836 22942 45892
rect 24406 45836 24444 45892
rect 24500 45836 24510 45892
rect 25666 45836 25676 45892
rect 25732 45836 26684 45892
rect 26740 45836 26750 45892
rect 28326 45836 28364 45892
rect 28420 45836 28430 45892
rect 17602 45724 17612 45780
rect 17668 45724 18396 45780
rect 18452 45724 18462 45780
rect 19058 45724 19068 45780
rect 19124 45724 19852 45780
rect 19908 45724 20748 45780
rect 20804 45724 21084 45780
rect 21140 45724 21150 45780
rect 22082 45724 22092 45780
rect 22148 45724 22764 45780
rect 22820 45724 22830 45780
rect 23874 45724 23884 45780
rect 23940 45724 26796 45780
rect 26852 45724 26862 45780
rect 28130 45724 28140 45780
rect 28196 45724 29036 45780
rect 29092 45724 29102 45780
rect 22092 45668 22148 45724
rect 3266 45612 3276 45668
rect 3332 45612 3612 45668
rect 3668 45612 3678 45668
rect 12226 45612 12236 45668
rect 12292 45612 16940 45668
rect 16996 45612 17006 45668
rect 17500 45612 22148 45668
rect 34962 45612 34972 45668
rect 35028 45612 38108 45668
rect 38164 45612 38174 45668
rect 17500 45556 17556 45612
rect 16034 45500 16044 45556
rect 16100 45500 17388 45556
rect 17444 45500 17556 45556
rect 22866 45500 22876 45556
rect 22932 45500 24220 45556
rect 24276 45500 24286 45556
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 19394 45388 19404 45444
rect 19460 45388 19684 45444
rect 23174 45388 23212 45444
rect 23268 45388 23278 45444
rect 28214 45388 28252 45444
rect 28308 45388 28318 45444
rect 19628 45332 19684 45388
rect 4162 45276 4172 45332
rect 4228 45276 4956 45332
rect 5012 45276 5628 45332
rect 5684 45276 5694 45332
rect 14354 45276 14364 45332
rect 14420 45276 15148 45332
rect 15204 45276 15214 45332
rect 19628 45276 21980 45332
rect 22036 45276 22046 45332
rect 22194 45276 22204 45332
rect 22260 45276 23100 45332
rect 23156 45276 28476 45332
rect 28532 45276 28588 45332
rect 28644 45276 28654 45332
rect 21634 45164 21644 45220
rect 21700 45164 23772 45220
rect 23828 45164 23838 45220
rect 24770 45164 24780 45220
rect 24836 45164 26012 45220
rect 26068 45164 26078 45220
rect 26338 45164 26348 45220
rect 26404 45164 26572 45220
rect 26628 45164 26638 45220
rect 27570 45164 27580 45220
rect 27636 45164 28364 45220
rect 28420 45164 28588 45220
rect 28644 45164 28654 45220
rect 0 45108 400 45136
rect 26012 45108 26068 45164
rect 0 45052 3500 45108
rect 3556 45052 3566 45108
rect 14018 45052 14028 45108
rect 14084 45052 15372 45108
rect 15428 45052 16716 45108
rect 16772 45052 16782 45108
rect 21522 45052 21532 45108
rect 21588 45052 23436 45108
rect 23492 45052 23502 45108
rect 23650 45052 23660 45108
rect 23716 45052 24668 45108
rect 24724 45052 24734 45108
rect 26012 45052 26908 45108
rect 26964 45052 27356 45108
rect 27412 45052 27422 45108
rect 0 45024 400 45052
rect 11890 44940 11900 44996
rect 11956 44940 12460 44996
rect 12516 44940 12526 44996
rect 16818 44940 16828 44996
rect 16884 44940 17500 44996
rect 17556 44940 17566 44996
rect 7634 44828 7644 44884
rect 7700 44828 8316 44884
rect 8372 44828 8382 44884
rect 16258 44828 16268 44884
rect 16324 44828 17052 44884
rect 17108 44828 17118 44884
rect 18498 44828 18508 44884
rect 18564 44828 20748 44884
rect 20804 44828 21308 44884
rect 21364 44828 21374 44884
rect 24210 44828 24220 44884
rect 24276 44828 24892 44884
rect 24948 44828 25788 44884
rect 25844 44828 25854 44884
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 21158 44604 21196 44660
rect 21252 44604 21262 44660
rect 26562 44604 26572 44660
rect 26628 44604 27580 44660
rect 27636 44604 29036 44660
rect 29092 44604 30828 44660
rect 30884 44604 31948 44660
rect 32004 44604 32014 44660
rect 21494 44492 21532 44548
rect 21588 44492 21598 44548
rect 23538 44492 23548 44548
rect 23604 44492 30492 44548
rect 30548 44492 30558 44548
rect 17378 44380 17388 44436
rect 17444 44380 18732 44436
rect 18788 44380 18798 44436
rect 20290 44380 20300 44436
rect 20356 44380 21868 44436
rect 21924 44380 21934 44436
rect 22530 44380 22540 44436
rect 22596 44380 24108 44436
rect 24164 44380 24174 44436
rect 27346 44380 27356 44436
rect 27412 44380 29708 44436
rect 29764 44380 30156 44436
rect 30212 44380 30222 44436
rect 30902 44380 30940 44436
rect 30996 44380 31006 44436
rect 30156 44324 30212 44380
rect 2258 44268 2268 44324
rect 2324 44268 3612 44324
rect 3668 44268 3678 44324
rect 10546 44268 10556 44324
rect 10612 44268 21308 44324
rect 21364 44268 22876 44324
rect 22932 44268 22942 44324
rect 30156 44268 32396 44324
rect 32452 44268 32462 44324
rect 3602 44156 3612 44212
rect 3668 44156 4844 44212
rect 4900 44156 4910 44212
rect 15250 44156 15260 44212
rect 15316 44156 15932 44212
rect 15988 44156 16380 44212
rect 16436 44156 16446 44212
rect 17042 44156 17052 44212
rect 17108 44156 17724 44212
rect 17780 44156 17790 44212
rect 25554 44156 25564 44212
rect 25620 44156 29260 44212
rect 29316 44156 29326 44212
rect 30594 44156 30604 44212
rect 30660 44156 30828 44212
rect 30884 44156 30894 44212
rect 15586 44044 15596 44100
rect 15652 44044 16716 44100
rect 16772 44044 17836 44100
rect 17892 44044 17902 44100
rect 27906 44044 27916 44100
rect 27972 44044 30380 44100
rect 30436 44044 32844 44100
rect 32900 44044 35644 44100
rect 35700 44044 35710 44100
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 20402 43820 20412 43876
rect 20468 43820 21196 43876
rect 21252 43820 21262 43876
rect 23762 43820 23772 43876
rect 23828 43820 25564 43876
rect 25620 43820 25630 43876
rect 23202 43708 23212 43764
rect 23268 43708 27076 43764
rect 27020 43652 27076 43708
rect 3938 43596 3948 43652
rect 4004 43596 4844 43652
rect 4900 43596 4910 43652
rect 15138 43596 15148 43652
rect 15204 43596 16940 43652
rect 16996 43596 19068 43652
rect 19124 43596 19134 43652
rect 22642 43596 22652 43652
rect 22708 43596 23660 43652
rect 23716 43596 23726 43652
rect 26338 43596 26348 43652
rect 26404 43596 26796 43652
rect 26852 43596 26862 43652
rect 27010 43596 27020 43652
rect 27076 43596 27086 43652
rect 27346 43596 27356 43652
rect 27412 43596 27916 43652
rect 27972 43596 27982 43652
rect 33170 43596 33180 43652
rect 33236 43596 34972 43652
rect 35028 43596 35868 43652
rect 35924 43596 35934 43652
rect 5506 43484 5516 43540
rect 5572 43484 6188 43540
rect 6244 43484 6254 43540
rect 16146 43484 16156 43540
rect 16212 43484 21644 43540
rect 21700 43484 21710 43540
rect 22194 43484 22204 43540
rect 22260 43484 22540 43540
rect 22596 43484 22606 43540
rect 23426 43484 23436 43540
rect 23492 43484 24108 43540
rect 24164 43484 24174 43540
rect 26562 43484 26572 43540
rect 26628 43484 29484 43540
rect 29540 43484 29550 43540
rect 8978 43372 8988 43428
rect 9044 43372 10220 43428
rect 10276 43372 10286 43428
rect 16818 43372 16828 43428
rect 16884 43372 19852 43428
rect 19908 43372 21532 43428
rect 21588 43372 21598 43428
rect 25554 43372 25564 43428
rect 25620 43372 26460 43428
rect 26516 43372 26526 43428
rect 26852 43372 27132 43428
rect 27188 43372 27198 43428
rect 29586 43372 29596 43428
rect 29652 43372 30828 43428
rect 30884 43372 30894 43428
rect 33058 43372 33068 43428
rect 33124 43372 34636 43428
rect 34692 43372 34702 43428
rect 15474 43260 15484 43316
rect 15540 43260 21868 43316
rect 21924 43260 21934 43316
rect 15362 43148 15372 43204
rect 15428 43148 19068 43204
rect 19124 43148 20412 43204
rect 20468 43148 20478 43204
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 26852 43092 26908 43372
rect 27010 43260 27020 43316
rect 27076 43260 27524 43316
rect 30034 43260 30044 43316
rect 30100 43260 30716 43316
rect 30772 43260 30940 43316
rect 30996 43260 31006 43316
rect 27468 43204 27524 43260
rect 27458 43148 27468 43204
rect 27524 43148 31388 43204
rect 31444 43148 31454 43204
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 16370 43036 16380 43092
rect 16436 43036 16716 43092
rect 16772 43036 21196 43092
rect 21252 43036 22540 43092
rect 22596 43036 23212 43092
rect 23268 43036 23278 43092
rect 26674 43036 26684 43092
rect 26740 43036 29484 43092
rect 29540 43036 31500 43092
rect 31556 43036 32284 43092
rect 32340 43036 32350 43092
rect 6178 42924 6188 42980
rect 6244 42924 6636 42980
rect 6692 42924 6702 42980
rect 30930 42924 30940 42980
rect 30996 42924 31164 42980
rect 31220 42924 31230 42980
rect 35522 42924 35532 42980
rect 35588 42924 36876 42980
rect 36932 42924 36942 42980
rect 20710 42812 20748 42868
rect 20804 42812 21308 42868
rect 21364 42812 21374 42868
rect 29922 42812 29932 42868
rect 29988 42812 30604 42868
rect 30660 42812 30670 42868
rect 35858 42812 35868 42868
rect 35924 42812 36428 42868
rect 36484 42812 38220 42868
rect 38276 42812 38286 42868
rect 4834 42700 4844 42756
rect 4900 42700 5068 42756
rect 5124 42700 5852 42756
rect 5908 42700 5918 42756
rect 6290 42700 6300 42756
rect 6356 42700 6636 42756
rect 6692 42700 9884 42756
rect 9940 42700 9950 42756
rect 10322 42700 10332 42756
rect 10388 42700 11228 42756
rect 11284 42700 11294 42756
rect 28130 42700 28140 42756
rect 28196 42700 28364 42756
rect 28420 42700 34524 42756
rect 34580 42700 34590 42756
rect 9986 42588 9996 42644
rect 10052 42588 11060 42644
rect 11004 42532 11060 42588
rect 11788 42588 15036 42644
rect 15092 42588 16772 42644
rect 24658 42588 24668 42644
rect 24724 42588 25788 42644
rect 25844 42588 25854 42644
rect 36418 42588 36428 42644
rect 36484 42588 36988 42644
rect 37044 42588 37054 42644
rect 9314 42476 9324 42532
rect 9380 42476 10108 42532
rect 10164 42476 10174 42532
rect 10994 42476 11004 42532
rect 11060 42476 11452 42532
rect 11508 42476 11518 42532
rect 11788 42420 11844 42588
rect 16716 42532 16772 42588
rect 16706 42476 16716 42532
rect 16772 42476 16782 42532
rect 23762 42476 23772 42532
rect 23828 42476 25340 42532
rect 25396 42476 25406 42532
rect 31938 42476 31948 42532
rect 32004 42476 32396 42532
rect 32452 42476 33180 42532
rect 33236 42476 33246 42532
rect 5506 42364 5516 42420
rect 5572 42364 11844 42420
rect 20626 42364 20636 42420
rect 20692 42364 25676 42420
rect 25732 42364 26684 42420
rect 26740 42364 26750 42420
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 14354 42252 14364 42308
rect 14420 42252 15932 42308
rect 15988 42252 15998 42308
rect 23538 42252 23548 42308
rect 23604 42252 24332 42308
rect 24388 42252 26236 42308
rect 26292 42252 28924 42308
rect 28980 42252 29708 42308
rect 29764 42252 29774 42308
rect 14802 42140 14812 42196
rect 14868 42140 15484 42196
rect 15540 42140 16940 42196
rect 16996 42140 17006 42196
rect 19506 42140 19516 42196
rect 19572 42140 21868 42196
rect 21924 42140 21934 42196
rect 25442 42140 25452 42196
rect 25508 42140 26684 42196
rect 26740 42140 28476 42196
rect 28532 42140 28542 42196
rect 29922 42140 29932 42196
rect 29988 42140 30380 42196
rect 30436 42140 35308 42196
rect 35364 42140 35374 42196
rect 5842 42028 5852 42084
rect 5908 42028 9996 42084
rect 10052 42028 10062 42084
rect 10322 42028 10332 42084
rect 10388 42028 10398 42084
rect 20066 42028 20076 42084
rect 20132 42028 20748 42084
rect 20804 42028 20814 42084
rect 21494 42028 21532 42084
rect 21588 42028 21598 42084
rect 24322 42028 24332 42084
rect 24388 42028 26348 42084
rect 26404 42028 26414 42084
rect 30818 42028 30828 42084
rect 30884 42028 31276 42084
rect 31332 42028 31342 42084
rect 7308 41972 7364 42028
rect 10332 41972 10388 42028
rect 6066 41916 6076 41972
rect 6132 41916 6142 41972
rect 7298 41916 7308 41972
rect 7364 41916 7374 41972
rect 8082 41916 8092 41972
rect 8148 41916 10388 41972
rect 11666 41916 11676 41972
rect 11732 41916 13244 41972
rect 13300 41916 14588 41972
rect 14644 41916 14654 41972
rect 16930 41916 16940 41972
rect 16996 41916 18060 41972
rect 18116 41916 19180 41972
rect 19236 41916 19246 41972
rect 19506 41916 19516 41972
rect 19572 41916 20300 41972
rect 20356 41916 20748 41972
rect 20804 41916 20814 41972
rect 22390 41916 22428 41972
rect 22484 41916 22494 41972
rect 23986 41916 23996 41972
rect 24052 41916 24062 41972
rect 24994 41916 25004 41972
rect 25060 41916 25228 41972
rect 25284 41916 26236 41972
rect 26292 41916 26302 41972
rect 27234 41916 27244 41972
rect 27300 41916 27692 41972
rect 27748 41916 30492 41972
rect 30548 41916 30558 41972
rect 6076 41860 6132 41916
rect 6076 41804 7196 41860
rect 7252 41804 7262 41860
rect 6076 41748 6132 41804
rect 8092 41748 8148 41916
rect 23996 41860 24052 41916
rect 9762 41804 9772 41860
rect 9828 41804 11340 41860
rect 11396 41804 15036 41860
rect 5282 41692 5292 41748
rect 5348 41692 6132 41748
rect 6290 41692 6300 41748
rect 6356 41692 7420 41748
rect 7476 41692 8148 41748
rect 4946 41580 4956 41636
rect 5012 41580 6972 41636
rect 7028 41580 7644 41636
rect 7700 41580 7710 41636
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 15092 41412 15148 41860
rect 23996 41804 28252 41860
rect 28308 41804 28318 41860
rect 31490 41804 31500 41860
rect 31556 41804 32284 41860
rect 32340 41804 32350 41860
rect 39600 41748 40000 41776
rect 21634 41692 21644 41748
rect 21700 41692 22540 41748
rect 22596 41692 23324 41748
rect 23380 41692 23390 41748
rect 23538 41692 23548 41748
rect 23604 41692 26068 41748
rect 26226 41692 26236 41748
rect 26292 41692 29260 41748
rect 29316 41692 30940 41748
rect 30996 41692 31444 41748
rect 38210 41692 38220 41748
rect 38276 41692 40000 41748
rect 20626 41580 20636 41636
rect 20692 41580 22652 41636
rect 22708 41580 24220 41636
rect 24276 41580 24286 41636
rect 26012 41524 26068 41692
rect 31388 41636 31444 41692
rect 39600 41664 40000 41692
rect 31378 41580 31388 41636
rect 31444 41580 31454 41636
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 22082 41468 22092 41524
rect 22148 41468 22988 41524
rect 23044 41468 23054 41524
rect 23874 41468 23884 41524
rect 23940 41468 24780 41524
rect 24836 41468 24846 41524
rect 26012 41468 26236 41524
rect 26292 41468 26302 41524
rect 30902 41468 30940 41524
rect 30996 41468 31006 41524
rect 15092 41356 15372 41412
rect 15428 41356 15438 41412
rect 22642 41356 22652 41412
rect 22708 41356 28364 41412
rect 28420 41356 30492 41412
rect 30548 41356 31500 41412
rect 31556 41356 31566 41412
rect 32162 41356 32172 41412
rect 32228 41356 37436 41412
rect 37492 41356 37502 41412
rect 12898 41244 12908 41300
rect 12964 41244 15148 41300
rect 15204 41244 15214 41300
rect 21522 41244 21532 41300
rect 21588 41244 22876 41300
rect 22932 41244 24108 41300
rect 24164 41244 27468 41300
rect 27524 41244 27534 41300
rect 32722 41244 32732 41300
rect 32788 41244 35308 41300
rect 35364 41244 35756 41300
rect 35812 41244 36092 41300
rect 36148 41244 37100 41300
rect 37156 41244 37166 41300
rect 14802 41132 14812 41188
rect 14868 41132 16380 41188
rect 16436 41132 16446 41188
rect 21298 41132 21308 41188
rect 21364 41132 21868 41188
rect 21924 41132 22316 41188
rect 22372 41132 22382 41188
rect 22866 41132 22876 41188
rect 22932 41132 23212 41188
rect 23268 41132 23278 41188
rect 24434 41132 24444 41188
rect 24500 41132 25676 41188
rect 25732 41132 25742 41188
rect 15698 41020 15708 41076
rect 15764 41020 17836 41076
rect 17892 41020 17902 41076
rect 18498 41020 18508 41076
rect 18564 41020 19180 41076
rect 19236 41020 19516 41076
rect 19572 41020 22932 41076
rect 23762 41020 23772 41076
rect 23828 41020 24108 41076
rect 24164 41020 24174 41076
rect 26562 41020 26572 41076
rect 26628 41020 28140 41076
rect 28196 41020 28206 41076
rect 22876 40964 22932 41020
rect 15698 40908 15708 40964
rect 15764 40908 17052 40964
rect 17108 40908 17118 40964
rect 19180 40908 20076 40964
rect 20132 40908 20142 40964
rect 20850 40908 20860 40964
rect 20916 40908 22316 40964
rect 22372 40908 22382 40964
rect 22866 40908 22876 40964
rect 22932 40908 23548 40964
rect 27906 40908 27916 40964
rect 27972 40908 27982 40964
rect 19180 40852 19236 40908
rect 23492 40852 23548 40908
rect 6962 40796 6972 40852
rect 7028 40796 16492 40852
rect 16548 40796 16558 40852
rect 19170 40796 19180 40852
rect 19236 40796 19246 40852
rect 22194 40796 22204 40852
rect 22260 40796 22428 40852
rect 22484 40796 22494 40852
rect 23492 40796 24220 40852
rect 24276 40796 24286 40852
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 27916 40740 27972 40908
rect 16370 40684 16380 40740
rect 16436 40684 18508 40740
rect 18564 40684 18574 40740
rect 22082 40684 22092 40740
rect 22148 40684 23884 40740
rect 23940 40684 27972 40740
rect 4498 40572 4508 40628
rect 4564 40572 5740 40628
rect 5796 40572 5806 40628
rect 9986 40572 9996 40628
rect 10052 40572 13020 40628
rect 13076 40572 13692 40628
rect 13748 40572 13758 40628
rect 15362 40572 15372 40628
rect 15428 40572 22708 40628
rect 24210 40572 24220 40628
rect 24276 40572 24668 40628
rect 24724 40572 24734 40628
rect 25890 40572 25900 40628
rect 25956 40572 27804 40628
rect 27860 40572 27870 40628
rect 35410 40572 35420 40628
rect 35476 40572 36092 40628
rect 36148 40572 36158 40628
rect 22652 40516 22708 40572
rect 25900 40516 25956 40572
rect 3602 40460 3612 40516
rect 3668 40460 4284 40516
rect 4340 40460 4956 40516
rect 5012 40460 5022 40516
rect 13570 40460 13580 40516
rect 13636 40460 13646 40516
rect 13794 40460 13804 40516
rect 13860 40460 14364 40516
rect 14420 40460 16268 40516
rect 16324 40460 16334 40516
rect 16482 40460 16492 40516
rect 16548 40460 16828 40516
rect 16884 40460 16894 40516
rect 17602 40460 17612 40516
rect 17668 40460 18172 40516
rect 18228 40460 18238 40516
rect 18498 40460 18508 40516
rect 18564 40460 20300 40516
rect 20356 40460 20412 40516
rect 20468 40460 20478 40516
rect 22614 40460 22652 40516
rect 22708 40460 22718 40516
rect 22978 40460 22988 40516
rect 23044 40460 25956 40516
rect 13580 40404 13636 40460
rect 3154 40348 3164 40404
rect 3220 40348 3948 40404
rect 4004 40348 4014 40404
rect 5954 40348 5964 40404
rect 6020 40348 6972 40404
rect 7028 40348 7038 40404
rect 13580 40348 15596 40404
rect 15652 40348 15662 40404
rect 15922 40348 15932 40404
rect 15988 40348 17500 40404
rect 17556 40348 21756 40404
rect 21812 40348 23660 40404
rect 23716 40348 23726 40404
rect 29110 40348 29148 40404
rect 29204 40348 29214 40404
rect 5618 40236 5628 40292
rect 5684 40236 6524 40292
rect 6580 40236 6590 40292
rect 14914 40236 14924 40292
rect 14980 40236 17276 40292
rect 17332 40236 17342 40292
rect 22502 40236 22540 40292
rect 22596 40236 23436 40292
rect 23492 40236 23502 40292
rect 28578 40236 28588 40292
rect 28644 40236 30044 40292
rect 30100 40236 30110 40292
rect 34962 40236 34972 40292
rect 35028 40236 35644 40292
rect 35700 40236 35710 40292
rect 15698 40124 15708 40180
rect 15764 40124 17388 40180
rect 17444 40124 17454 40180
rect 26870 40124 26908 40180
rect 26964 40124 26974 40180
rect 35522 40124 35532 40180
rect 35588 40124 36204 40180
rect 36260 40124 36270 40180
rect 22194 40012 22204 40068
rect 22260 40012 22316 40068
rect 22372 40012 22382 40068
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 23986 39900 23996 39956
rect 24052 39900 24668 39956
rect 24724 39900 24734 39956
rect 24098 39788 24108 39844
rect 24164 39788 28308 39844
rect 30482 39788 30492 39844
rect 30548 39788 34300 39844
rect 34356 39788 34366 39844
rect 28252 39732 28308 39788
rect 5842 39676 5852 39732
rect 5908 39676 6748 39732
rect 6804 39676 6814 39732
rect 23650 39676 23660 39732
rect 23716 39676 24164 39732
rect 24434 39676 24444 39732
rect 24500 39676 25116 39732
rect 25172 39676 25182 39732
rect 28242 39676 28252 39732
rect 28308 39676 28318 39732
rect 31714 39676 31724 39732
rect 31780 39676 32508 39732
rect 32564 39676 32574 39732
rect 35186 39676 35196 39732
rect 35252 39676 35756 39732
rect 35812 39676 35822 39732
rect 5590 39564 5628 39620
rect 5684 39564 5694 39620
rect 11442 39564 11452 39620
rect 11508 39564 12908 39620
rect 12964 39564 15148 39620
rect 15204 39564 22204 39620
rect 22260 39564 22270 39620
rect 5170 39452 5180 39508
rect 5236 39452 6300 39508
rect 6356 39452 7196 39508
rect 7252 39452 7262 39508
rect 14028 39452 16156 39508
rect 16212 39452 16222 39508
rect 19506 39452 19516 39508
rect 19572 39452 21644 39508
rect 21700 39452 21710 39508
rect 14028 39396 14084 39452
rect 24108 39396 24164 39676
rect 25666 39564 25676 39620
rect 25732 39564 26460 39620
rect 26516 39564 26526 39620
rect 31938 39564 31948 39620
rect 32004 39564 33180 39620
rect 33236 39564 33740 39620
rect 33796 39564 33806 39620
rect 35298 39564 35308 39620
rect 35364 39564 36428 39620
rect 36484 39564 36494 39620
rect 24882 39452 24892 39508
rect 24948 39452 25340 39508
rect 25396 39452 25406 39508
rect 26002 39452 26012 39508
rect 26068 39452 27468 39508
rect 27524 39452 27534 39508
rect 3714 39340 3724 39396
rect 3780 39340 6076 39396
rect 6132 39340 6142 39396
rect 7970 39340 7980 39396
rect 8036 39340 12460 39396
rect 12516 39340 14028 39396
rect 14084 39340 14094 39396
rect 14914 39340 14924 39396
rect 14980 39340 20244 39396
rect 22194 39340 22204 39396
rect 22260 39340 22428 39396
rect 22484 39340 22494 39396
rect 24098 39340 24108 39396
rect 24164 39340 24174 39396
rect 24434 39340 24444 39396
rect 24500 39340 25900 39396
rect 25956 39340 25966 39396
rect 15026 39228 15036 39284
rect 15092 39228 15932 39284
rect 15988 39228 15998 39284
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 20188 39172 20244 39340
rect 27122 39228 27132 39284
rect 27188 39228 30492 39284
rect 30548 39228 30558 39284
rect 20188 39116 26460 39172
rect 26516 39116 26526 39172
rect 35252 39116 35532 39172
rect 35588 39116 35598 39172
rect 4610 39004 4620 39060
rect 4676 39004 5516 39060
rect 5572 39004 5852 39060
rect 5908 39004 5918 39060
rect 18386 39004 18396 39060
rect 18452 39004 19180 39060
rect 19236 39004 19246 39060
rect 20402 39004 20412 39060
rect 20468 39004 22092 39060
rect 22148 39004 22158 39060
rect 24406 39004 24444 39060
rect 24500 39004 24510 39060
rect 25778 39004 25788 39060
rect 25844 39004 26236 39060
rect 26292 39004 26302 39060
rect 35252 38948 35308 39116
rect 6850 38892 6860 38948
rect 6916 38892 16492 38948
rect 16548 38892 16558 38948
rect 21644 38892 23324 38948
rect 23380 38892 23390 38948
rect 27244 38892 30604 38948
rect 30660 38892 33180 38948
rect 33236 38892 35308 38948
rect 5170 38780 5180 38836
rect 5236 38780 5908 38836
rect 15922 38780 15932 38836
rect 15988 38780 16044 38836
rect 16100 38780 16110 38836
rect 16482 38780 16492 38836
rect 16548 38780 18620 38836
rect 18676 38780 18686 38836
rect 19170 38780 19180 38836
rect 19236 38780 19516 38836
rect 19572 38780 19582 38836
rect 5852 38724 5908 38780
rect 21644 38724 21700 38892
rect 27244 38836 27300 38892
rect 22194 38780 22204 38836
rect 22260 38780 22764 38836
rect 22820 38780 27244 38836
rect 27300 38780 27310 38836
rect 30482 38780 30492 38836
rect 30548 38780 32172 38836
rect 32228 38780 32238 38836
rect 1922 38668 1932 38724
rect 1988 38668 5628 38724
rect 5684 38668 5694 38724
rect 5852 38668 16212 38724
rect 16818 38668 16828 38724
rect 16884 38668 17612 38724
rect 17668 38668 18956 38724
rect 19012 38668 19022 38724
rect 20290 38668 20300 38724
rect 20356 38668 21644 38724
rect 21700 38668 21710 38724
rect 31378 38668 31388 38724
rect 31444 38668 31836 38724
rect 31892 38668 31902 38724
rect 4722 38556 4732 38612
rect 4788 38556 5964 38612
rect 6020 38556 6030 38612
rect 16156 38500 16212 38668
rect 16342 38556 16380 38612
rect 16436 38556 16446 38612
rect 22614 38556 22652 38612
rect 22708 38556 22718 38612
rect 30706 38556 30716 38612
rect 30772 38556 31612 38612
rect 31668 38556 31678 38612
rect 16156 38444 16828 38500
rect 16884 38444 16894 38500
rect 18274 38444 18284 38500
rect 18340 38444 19404 38500
rect 19460 38444 19470 38500
rect 22278 38444 22316 38500
rect 22372 38444 22382 38500
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 22418 38332 22428 38388
rect 22484 38332 22540 38388
rect 22596 38332 23436 38388
rect 23492 38332 23502 38388
rect 15250 38220 15260 38276
rect 15316 38220 24332 38276
rect 24388 38220 24398 38276
rect 4834 38108 4844 38164
rect 4900 38108 5404 38164
rect 5460 38108 7420 38164
rect 7476 38108 7486 38164
rect 13346 38108 13356 38164
rect 13412 38108 14812 38164
rect 14868 38108 15148 38164
rect 15922 38108 15932 38164
rect 15988 38108 16380 38164
rect 16436 38108 16446 38164
rect 23090 38108 23100 38164
rect 23156 38108 23660 38164
rect 23716 38108 24108 38164
rect 24164 38108 24174 38164
rect 15092 38052 15148 38108
rect 10210 37996 10220 38052
rect 10276 37996 11452 38052
rect 11508 37996 11518 38052
rect 15092 37996 15820 38052
rect 15876 37996 15886 38052
rect 20300 37996 20748 38052
rect 20804 37996 20814 38052
rect 36418 37996 36428 38052
rect 36484 37996 37772 38052
rect 37828 37996 37838 38052
rect 20300 37940 20356 37996
rect 9538 37884 9548 37940
rect 9604 37884 10668 37940
rect 10724 37884 10734 37940
rect 10994 37884 11004 37940
rect 11060 37884 20356 37940
rect 20514 37884 20524 37940
rect 20580 37884 21644 37940
rect 21700 37884 21710 37940
rect 21858 37884 21868 37940
rect 21924 37884 22204 37940
rect 22260 37884 23100 37940
rect 23156 37884 23166 37940
rect 36978 37884 36988 37940
rect 37044 37884 37548 37940
rect 37604 37884 37614 37940
rect 3266 37772 3276 37828
rect 3332 37772 4284 37828
rect 4340 37772 4350 37828
rect 4610 37772 4620 37828
rect 4676 37772 5068 37828
rect 5124 37772 9772 37828
rect 9828 37772 10556 37828
rect 10612 37772 13916 37828
rect 13972 37772 14588 37828
rect 14644 37772 14654 37828
rect 15558 37772 15596 37828
rect 15652 37772 15662 37828
rect 15894 37772 15932 37828
rect 15988 37772 15998 37828
rect 16482 37772 16492 37828
rect 16548 37772 16604 37828
rect 16660 37772 16670 37828
rect 17378 37772 17388 37828
rect 17444 37772 22148 37828
rect 25218 37772 25228 37828
rect 25284 37772 26012 37828
rect 26068 37772 26908 37828
rect 26964 37772 26974 37828
rect 33394 37772 33404 37828
rect 33460 37772 33852 37828
rect 33908 37772 33918 37828
rect 4620 37716 4676 37772
rect 3938 37660 3948 37716
rect 4004 37660 4676 37716
rect 16146 37660 16156 37716
rect 16212 37660 16716 37716
rect 16772 37660 16782 37716
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 22092 37604 22148 37772
rect 22092 37548 29148 37604
rect 29204 37548 29214 37604
rect 13020 37436 15372 37492
rect 15428 37436 15438 37492
rect 16370 37436 16380 37492
rect 16436 37436 16604 37492
rect 16660 37436 16670 37492
rect 16818 37436 16828 37492
rect 16884 37436 18284 37492
rect 18340 37436 18732 37492
rect 18788 37436 18798 37492
rect 19506 37436 19516 37492
rect 19572 37436 20300 37492
rect 20356 37436 22764 37492
rect 22820 37436 22830 37492
rect 23986 37436 23996 37492
rect 24052 37436 24668 37492
rect 24724 37436 25788 37492
rect 25844 37436 25854 37492
rect 28914 37436 28924 37492
rect 28980 37436 31052 37492
rect 31108 37436 31118 37492
rect 13020 37268 13076 37436
rect 16604 37380 16660 37436
rect 16604 37324 18620 37380
rect 18676 37324 18686 37380
rect 21746 37324 21756 37380
rect 21812 37324 22428 37380
rect 22484 37324 22494 37380
rect 27122 37324 27132 37380
rect 27188 37324 28140 37380
rect 28196 37324 28252 37380
rect 28308 37324 28318 37380
rect 3826 37212 3836 37268
rect 3892 37212 5180 37268
rect 5236 37212 5628 37268
rect 5684 37212 5694 37268
rect 12562 37212 12572 37268
rect 12628 37212 13076 37268
rect 20290 37212 20300 37268
rect 20356 37212 21084 37268
rect 21140 37212 21150 37268
rect 13020 37156 13076 37212
rect 6738 37100 6748 37156
rect 6804 37100 10220 37156
rect 10276 37100 10286 37156
rect 11666 37100 11676 37156
rect 11732 37100 12236 37156
rect 12292 37100 12302 37156
rect 13010 37100 13020 37156
rect 13076 37100 13086 37156
rect 17042 37100 17052 37156
rect 17108 37100 17724 37156
rect 17780 37100 17790 37156
rect 24546 37100 24556 37156
rect 24612 37100 25340 37156
rect 25396 37100 25788 37156
rect 25844 37100 25854 37156
rect 35298 37100 35308 37156
rect 35364 37100 35868 37156
rect 35924 37100 35934 37156
rect 36418 37100 36428 37156
rect 36484 37100 37436 37156
rect 37492 37100 37502 37156
rect 12674 36988 12684 37044
rect 12740 36988 19964 37044
rect 20020 36988 21084 37044
rect 21140 36988 21150 37044
rect 33842 36988 33852 37044
rect 33908 36988 35588 37044
rect 6514 36876 6524 36932
rect 6580 36876 6748 36932
rect 6804 36876 6814 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 17266 36764 17276 36820
rect 17332 36764 17836 36820
rect 17892 36764 17902 36820
rect 35532 36708 35588 36988
rect 4162 36652 4172 36708
rect 4228 36652 4508 36708
rect 4564 36652 6076 36708
rect 6132 36652 6142 36708
rect 20514 36652 20524 36708
rect 20580 36652 30268 36708
rect 30324 36652 30334 36708
rect 35522 36652 35532 36708
rect 35588 36652 35598 36708
rect 7522 36540 7532 36596
rect 7588 36540 8540 36596
rect 8596 36540 9100 36596
rect 9156 36540 9166 36596
rect 12002 36540 12012 36596
rect 12068 36540 15148 36596
rect 15204 36540 16828 36596
rect 16884 36540 17276 36596
rect 17332 36540 17342 36596
rect 17826 36540 17836 36596
rect 17892 36540 18508 36596
rect 18564 36540 18574 36596
rect 5842 36428 5852 36484
rect 5908 36428 6748 36484
rect 6804 36428 9772 36484
rect 9828 36428 10668 36484
rect 10724 36428 10734 36484
rect 19590 36428 19628 36484
rect 19684 36428 19694 36484
rect 22978 36428 22988 36484
rect 23044 36428 23996 36484
rect 24052 36428 24062 36484
rect 4274 36316 4284 36372
rect 4340 36316 5628 36372
rect 5684 36316 5694 36372
rect 22418 36316 22428 36372
rect 22484 36316 23604 36372
rect 24322 36316 24332 36372
rect 24388 36316 26012 36372
rect 26068 36316 26078 36372
rect 23548 36260 23604 36316
rect 9874 36204 9884 36260
rect 9940 36204 19628 36260
rect 19684 36204 19694 36260
rect 21522 36204 21532 36260
rect 21588 36204 22204 36260
rect 22260 36204 22270 36260
rect 22978 36204 22988 36260
rect 23044 36204 23212 36260
rect 23268 36204 23278 36260
rect 23538 36204 23548 36260
rect 23604 36204 25004 36260
rect 25060 36204 25070 36260
rect 28354 36204 28364 36260
rect 28420 36204 31836 36260
rect 31892 36204 32844 36260
rect 32900 36204 32910 36260
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 22194 35980 22204 36036
rect 22260 35980 24220 36036
rect 24276 35980 24286 36036
rect 9090 35868 9100 35924
rect 9156 35868 9884 35924
rect 9940 35868 9950 35924
rect 19954 35868 19964 35924
rect 20020 35868 20860 35924
rect 20916 35868 20926 35924
rect 28130 35868 28140 35924
rect 28196 35868 31052 35924
rect 31108 35868 31118 35924
rect 6402 35756 6412 35812
rect 6468 35756 17500 35812
rect 17556 35756 17566 35812
rect 26674 35756 26684 35812
rect 26740 35756 28924 35812
rect 28980 35756 28990 35812
rect 30594 35756 30604 35812
rect 30660 35756 32396 35812
rect 32452 35756 32462 35812
rect 35746 35756 35756 35812
rect 35812 35756 36988 35812
rect 37044 35756 37054 35812
rect 3602 35644 3612 35700
rect 3668 35644 4732 35700
rect 4788 35644 5516 35700
rect 5572 35644 5582 35700
rect 6178 35644 6188 35700
rect 6244 35644 6636 35700
rect 6692 35644 7196 35700
rect 7252 35644 10108 35700
rect 10164 35644 11116 35700
rect 11172 35644 11182 35700
rect 12898 35644 12908 35700
rect 12964 35644 15596 35700
rect 15652 35644 15662 35700
rect 17042 35644 17052 35700
rect 17108 35644 17948 35700
rect 18004 35644 18014 35700
rect 18582 35644 18620 35700
rect 18676 35644 18686 35700
rect 28466 35644 28476 35700
rect 28532 35644 29148 35700
rect 29204 35644 29214 35700
rect 17948 35588 18004 35644
rect 15810 35532 15820 35588
rect 15876 35532 17388 35588
rect 17444 35532 17454 35588
rect 17948 35532 18732 35588
rect 18788 35532 18798 35588
rect 19282 35532 19292 35588
rect 19348 35532 20076 35588
rect 20132 35532 20142 35588
rect 32162 35532 32172 35588
rect 32228 35532 32956 35588
rect 33012 35532 33022 35588
rect 36082 35532 36092 35588
rect 36148 35532 36764 35588
rect 36820 35532 37212 35588
rect 37268 35532 37278 35588
rect 14914 35420 14924 35476
rect 14980 35420 15372 35476
rect 15428 35420 15932 35476
rect 15988 35420 15998 35476
rect 18050 35420 18060 35476
rect 18116 35420 18126 35476
rect 18386 35420 18396 35476
rect 18452 35420 27356 35476
rect 27412 35420 27422 35476
rect 32834 35420 32844 35476
rect 32900 35420 36428 35476
rect 36484 35420 36494 35476
rect 18060 35364 18116 35420
rect 3602 35308 3612 35364
rect 3668 35308 3678 35364
rect 5506 35308 5516 35364
rect 5572 35308 7084 35364
rect 7140 35308 7150 35364
rect 18060 35308 18284 35364
rect 18340 35308 18350 35364
rect 19590 35308 19628 35364
rect 19684 35308 19694 35364
rect 22306 35308 22316 35364
rect 22372 35308 23772 35364
rect 23828 35308 23838 35364
rect 35970 35308 35980 35364
rect 36036 35308 36988 35364
rect 37044 35308 37054 35364
rect 0 35252 400 35280
rect 3612 35252 3668 35308
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 0 35196 3164 35252
rect 3220 35196 3230 35252
rect 3602 35196 3612 35252
rect 3668 35196 3678 35252
rect 6290 35196 6300 35252
rect 6356 35196 6524 35252
rect 6580 35196 6590 35252
rect 6738 35196 6748 35252
rect 6804 35196 7196 35252
rect 7252 35196 7262 35252
rect 31154 35196 31164 35252
rect 31220 35196 33740 35252
rect 33796 35196 33806 35252
rect 35606 35196 35644 35252
rect 35700 35196 35710 35252
rect 0 35168 400 35196
rect 17686 35084 17724 35140
rect 17780 35084 17790 35140
rect 17500 34972 18172 35028
rect 18228 34972 18238 35028
rect 18918 34972 18956 35028
rect 19012 34972 19022 35028
rect 35410 34972 35420 35028
rect 35476 34972 35644 35028
rect 35700 34972 35710 35028
rect 17500 34916 17556 34972
rect 5954 34860 5964 34916
rect 6020 34860 7420 34916
rect 7476 34860 7486 34916
rect 17490 34860 17500 34916
rect 17556 34860 17566 34916
rect 25218 34860 25228 34916
rect 25284 34860 25564 34916
rect 25620 34860 26684 34916
rect 26740 34860 26750 34916
rect 30258 34860 30268 34916
rect 30324 34860 30828 34916
rect 30884 34860 34076 34916
rect 34132 34860 35084 34916
rect 35140 34860 35868 34916
rect 35924 34860 35934 34916
rect 18162 34748 18172 34804
rect 18228 34748 19628 34804
rect 19684 34748 19694 34804
rect 31602 34748 31612 34804
rect 31668 34748 32732 34804
rect 32788 34748 32798 34804
rect 33730 34748 33740 34804
rect 33796 34748 35532 34804
rect 35588 34748 35644 34804
rect 35700 34748 35710 34804
rect 15138 34636 15148 34692
rect 15204 34636 15820 34692
rect 15876 34636 15886 34692
rect 18834 34636 18844 34692
rect 18900 34636 27020 34692
rect 27076 34636 27086 34692
rect 28242 34636 28252 34692
rect 28308 34636 34524 34692
rect 34580 34636 34590 34692
rect 17350 34524 17388 34580
rect 17444 34524 17454 34580
rect 18610 34524 18620 34580
rect 18676 34524 19180 34580
rect 19236 34524 19246 34580
rect 28690 34524 28700 34580
rect 28756 34524 30044 34580
rect 30100 34524 31948 34580
rect 32004 34524 32014 34580
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 6962 34300 6972 34356
rect 7028 34300 18060 34356
rect 18116 34300 18126 34356
rect 18946 34300 18956 34356
rect 19012 34300 19292 34356
rect 19348 34300 19358 34356
rect 30146 34300 30156 34356
rect 30212 34300 31948 34356
rect 32004 34300 32014 34356
rect 33394 34300 33404 34356
rect 33460 34300 34076 34356
rect 34132 34300 34142 34356
rect 35606 34300 35644 34356
rect 35700 34300 35710 34356
rect 36194 34300 36204 34356
rect 36260 34300 38220 34356
rect 38276 34300 38286 34356
rect 6738 34188 6748 34244
rect 6804 34188 7308 34244
rect 7364 34188 7374 34244
rect 35186 34188 35196 34244
rect 35252 34188 36876 34244
rect 36932 34188 36942 34244
rect 6178 34076 6188 34132
rect 6244 34076 7196 34132
rect 7252 34076 7756 34132
rect 7812 34076 7822 34132
rect 18386 34076 18396 34132
rect 18452 34076 18844 34132
rect 18900 34076 18910 34132
rect 22978 34076 22988 34132
rect 23044 34076 23548 34132
rect 23604 34076 23614 34132
rect 28130 34076 28140 34132
rect 28196 34076 31500 34132
rect 31556 34076 31566 34132
rect 4610 33964 4620 34020
rect 4676 33964 5852 34020
rect 5908 33964 5918 34020
rect 7410 33964 7420 34020
rect 7476 33964 9884 34020
rect 9940 33964 10108 34020
rect 10164 33964 10556 34020
rect 10612 33964 11564 34020
rect 11620 33964 11630 34020
rect 16146 33964 16156 34020
rect 16212 33964 17948 34020
rect 18004 33964 19852 34020
rect 19908 33964 19918 34020
rect 35522 33964 35532 34020
rect 35588 33964 36204 34020
rect 36260 33964 36270 34020
rect 6514 33852 6524 33908
rect 6580 33852 6860 33908
rect 6916 33852 6926 33908
rect 12226 33852 12236 33908
rect 12292 33852 12684 33908
rect 12740 33852 12750 33908
rect 16034 33852 16044 33908
rect 16100 33852 17612 33908
rect 17668 33852 19516 33908
rect 19572 33852 19582 33908
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 15810 33628 15820 33684
rect 15876 33628 22428 33684
rect 22484 33628 22494 33684
rect 23314 33628 23324 33684
rect 23380 33628 23548 33684
rect 23604 33628 23996 33684
rect 24052 33628 24062 33684
rect 11666 33516 11676 33572
rect 11732 33516 13580 33572
rect 13636 33516 13646 33572
rect 17378 33516 17388 33572
rect 17444 33516 17836 33572
rect 17892 33516 17902 33572
rect 19730 33516 19740 33572
rect 19796 33516 20748 33572
rect 20804 33516 21868 33572
rect 21924 33516 21934 33572
rect 27122 33516 27132 33572
rect 27188 33516 27692 33572
rect 27748 33516 27758 33572
rect 28578 33516 28588 33572
rect 28644 33516 29484 33572
rect 29540 33516 29550 33572
rect 31490 33516 31500 33572
rect 31556 33516 32172 33572
rect 32228 33516 32238 33572
rect 33058 33516 33068 33572
rect 33124 33516 33134 33572
rect 33068 33460 33124 33516
rect 17378 33404 17388 33460
rect 17444 33404 17612 33460
rect 17668 33404 17678 33460
rect 28466 33404 28476 33460
rect 28532 33404 33124 33460
rect 34290 33404 34300 33460
rect 34356 33404 34860 33460
rect 34916 33404 35308 33460
rect 35364 33404 35374 33460
rect 6178 33292 6188 33348
rect 6244 33292 6972 33348
rect 7028 33292 7038 33348
rect 28018 33292 28028 33348
rect 28084 33292 29260 33348
rect 29316 33292 29326 33348
rect 31490 33292 31500 33348
rect 31556 33292 34972 33348
rect 35028 33292 35532 33348
rect 35588 33292 36092 33348
rect 36148 33292 36158 33348
rect 36418 33292 36428 33348
rect 36484 33292 36876 33348
rect 36932 33292 36942 33348
rect 27346 33180 27356 33236
rect 27412 33180 28364 33236
rect 28420 33180 28430 33236
rect 35858 33180 35868 33236
rect 35924 33180 36988 33236
rect 37044 33180 37054 33236
rect 3938 33068 3948 33124
rect 4004 33068 4844 33124
rect 4900 33068 7420 33124
rect 7476 33068 7486 33124
rect 26450 33068 26460 33124
rect 26516 33068 27132 33124
rect 27188 33068 27198 33124
rect 25218 32956 25228 33012
rect 25284 32956 28812 33012
rect 28868 32956 28878 33012
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 14802 32844 14812 32900
rect 14868 32844 16828 32900
rect 16884 32844 17500 32900
rect 17556 32844 17836 32900
rect 17892 32844 17902 32900
rect 15586 32732 15596 32788
rect 15652 32732 17276 32788
rect 17332 32732 17342 32788
rect 7298 32620 7308 32676
rect 7364 32620 7756 32676
rect 7812 32620 8092 32676
rect 8148 32620 8158 32676
rect 31826 32620 31836 32676
rect 31892 32620 33068 32676
rect 33124 32620 33134 32676
rect 13570 32508 13580 32564
rect 13636 32508 15148 32564
rect 15204 32508 15214 32564
rect 2482 32396 2492 32452
rect 2548 32396 3948 32452
rect 4004 32396 4014 32452
rect 6402 32396 6412 32452
rect 6468 32396 6748 32452
rect 6804 32396 7084 32452
rect 7140 32396 7150 32452
rect 14690 32396 14700 32452
rect 14756 32396 15596 32452
rect 15652 32396 15662 32452
rect 17602 32284 17612 32340
rect 17668 32284 18060 32340
rect 18116 32284 30940 32340
rect 30996 32284 31006 32340
rect 35074 32284 35084 32340
rect 35140 32284 35868 32340
rect 35924 32284 35934 32340
rect 19170 32172 19180 32228
rect 19236 32172 19628 32228
rect 19684 32172 19694 32228
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 26898 31948 26908 32004
rect 26964 31948 29260 32004
rect 29316 31948 30044 32004
rect 30100 31948 30110 32004
rect 33842 31948 33852 32004
rect 33908 31948 35644 32004
rect 35700 31948 35710 32004
rect 9314 31836 9324 31892
rect 9380 31836 10556 31892
rect 10612 31836 10622 31892
rect 21410 31836 21420 31892
rect 21476 31836 23436 31892
rect 23492 31836 23502 31892
rect 5730 31724 5740 31780
rect 5796 31724 7308 31780
rect 7364 31724 7374 31780
rect 21298 31724 21308 31780
rect 21364 31724 21980 31780
rect 22036 31724 22046 31780
rect 24210 31724 24220 31780
rect 24276 31724 24668 31780
rect 24724 31724 25676 31780
rect 25732 31724 26684 31780
rect 26740 31724 26750 31780
rect 12226 31612 12236 31668
rect 12292 31612 15260 31668
rect 15316 31612 15820 31668
rect 15876 31612 26908 31668
rect 26964 31612 26974 31668
rect 36194 31612 36204 31668
rect 36260 31612 36988 31668
rect 37044 31612 37054 31668
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 7746 31164 7756 31220
rect 7812 31164 8988 31220
rect 9044 31164 10108 31220
rect 10164 31164 10174 31220
rect 23314 31164 23324 31220
rect 23380 31164 24220 31220
rect 24276 31164 24286 31220
rect 19506 31052 19516 31108
rect 19572 31052 19582 31108
rect 19516 30996 19572 31052
rect 15810 30940 15820 30996
rect 15876 30940 19852 30996
rect 19908 30940 19918 30996
rect 18946 30828 18956 30884
rect 19012 30828 19964 30884
rect 20020 30828 20030 30884
rect 30482 30828 30492 30884
rect 30548 30828 30716 30884
rect 30772 30828 31612 30884
rect 31668 30828 32396 30884
rect 32452 30828 32956 30884
rect 33012 30828 33022 30884
rect 33506 30828 33516 30884
rect 33572 30828 36428 30884
rect 36484 30828 38220 30884
rect 38276 30828 38286 30884
rect 10098 30716 10108 30772
rect 10164 30716 18060 30772
rect 18116 30716 18126 30772
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 13794 30380 13804 30436
rect 13860 30380 19404 30436
rect 19460 30380 19628 30436
rect 19684 30380 22876 30436
rect 22932 30380 23436 30436
rect 23492 30380 23502 30436
rect 18834 30268 18844 30324
rect 18900 30268 19180 30324
rect 19236 30268 19246 30324
rect 4722 30156 4732 30212
rect 4788 30156 5292 30212
rect 5348 30156 5358 30212
rect 7298 30156 7308 30212
rect 7364 30156 8092 30212
rect 8148 30156 8158 30212
rect 10546 30156 10556 30212
rect 10612 30156 11004 30212
rect 11060 30156 11070 30212
rect 18386 30156 18396 30212
rect 18452 30156 19964 30212
rect 20020 30156 20030 30212
rect 22754 30156 22764 30212
rect 22820 30156 23436 30212
rect 23492 30156 23502 30212
rect 31602 30156 31612 30212
rect 31668 30156 32732 30212
rect 32788 30156 32798 30212
rect 29810 30044 29820 30100
rect 29876 30044 30828 30100
rect 30884 30044 32060 30100
rect 32116 30044 32508 30100
rect 32564 30044 32574 30100
rect 20290 29932 20300 29988
rect 20356 29932 20366 29988
rect 22418 29932 22428 29988
rect 22484 29932 23100 29988
rect 23156 29932 23166 29988
rect 14242 29820 14252 29876
rect 14308 29820 15148 29876
rect 15204 29820 15932 29876
rect 15988 29820 19068 29876
rect 19124 29820 19134 29876
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 18498 29708 18508 29764
rect 18564 29708 18788 29764
rect 18732 29652 18788 29708
rect 3826 29596 3836 29652
rect 3892 29596 4732 29652
rect 4788 29596 4798 29652
rect 9874 29596 9884 29652
rect 9940 29596 10556 29652
rect 10612 29596 13244 29652
rect 13300 29596 13804 29652
rect 13860 29596 13870 29652
rect 16594 29596 16604 29652
rect 16660 29596 17388 29652
rect 17444 29596 17454 29652
rect 18722 29596 18732 29652
rect 18788 29596 18798 29652
rect 20300 29540 20356 29932
rect 23426 29596 23436 29652
rect 23492 29596 24108 29652
rect 24164 29596 24174 29652
rect 25890 29596 25900 29652
rect 25956 29596 27244 29652
rect 27300 29596 30716 29652
rect 30772 29596 31276 29652
rect 31332 29596 31342 29652
rect 33842 29596 33852 29652
rect 33908 29596 34748 29652
rect 34804 29596 34814 29652
rect 3938 29484 3948 29540
rect 4004 29484 4014 29540
rect 10770 29484 10780 29540
rect 10836 29484 11340 29540
rect 11396 29484 15484 29540
rect 15540 29484 15550 29540
rect 20290 29484 20300 29540
rect 20356 29484 20366 29540
rect 26562 29484 26572 29540
rect 26628 29484 26796 29540
rect 26852 29484 26862 29540
rect 3948 29316 4004 29484
rect 4610 29372 4620 29428
rect 4676 29372 5516 29428
rect 5572 29372 5582 29428
rect 14130 29372 14140 29428
rect 14196 29372 14700 29428
rect 14756 29372 14766 29428
rect 17042 29372 17052 29428
rect 17108 29372 17276 29428
rect 17332 29372 17342 29428
rect 19058 29372 19068 29428
rect 19124 29372 21196 29428
rect 21252 29372 21756 29428
rect 21812 29372 21822 29428
rect 26338 29372 26348 29428
rect 26404 29372 26684 29428
rect 26740 29372 29820 29428
rect 29876 29372 29886 29428
rect 3948 29260 4844 29316
rect 4900 29260 4910 29316
rect 24434 29260 24444 29316
rect 24500 29260 24780 29316
rect 24836 29260 24846 29316
rect 35298 29260 35308 29316
rect 35364 29260 35644 29316
rect 35700 29260 35710 29316
rect 26786 29148 26796 29204
rect 26852 29148 27804 29204
rect 27860 29148 27870 29204
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 12674 28812 12684 28868
rect 12740 28812 13468 28868
rect 13524 28812 13534 28868
rect 13692 28812 23772 28868
rect 23828 28812 23838 28868
rect 27458 28812 27468 28868
rect 27524 28812 30044 28868
rect 30100 28812 30716 28868
rect 30772 28812 31164 28868
rect 31220 28812 31230 28868
rect 13692 28756 13748 28812
rect 4620 28700 5292 28756
rect 5348 28700 5358 28756
rect 7970 28700 7980 28756
rect 8036 28700 8046 28756
rect 8194 28700 8204 28756
rect 8260 28700 13748 28756
rect 14018 28700 14028 28756
rect 14084 28700 18396 28756
rect 18452 28700 18462 28756
rect 4620 28644 4676 28700
rect 4162 28588 4172 28644
rect 4228 28588 4620 28644
rect 4676 28588 4686 28644
rect 4834 28588 4844 28644
rect 4900 28588 5012 28644
rect 6290 28588 6300 28644
rect 6356 28588 7084 28644
rect 7140 28588 7150 28644
rect 7298 28588 7308 28644
rect 7364 28588 7374 28644
rect 4956 28532 5012 28588
rect 7308 28532 7364 28588
rect 4956 28476 5740 28532
rect 5796 28476 5806 28532
rect 6066 28476 6076 28532
rect 6132 28476 6636 28532
rect 6692 28476 7364 28532
rect 7980 28308 8036 28700
rect 10098 28588 10108 28644
rect 10164 28588 13580 28644
rect 13636 28588 14140 28644
rect 14196 28588 15148 28644
rect 18582 28588 18620 28644
rect 18676 28588 18686 28644
rect 15092 28532 15148 28588
rect 15092 28476 16156 28532
rect 16212 28476 16222 28532
rect 17042 28476 17052 28532
rect 17108 28476 17948 28532
rect 18004 28476 20188 28532
rect 20244 28476 20524 28532
rect 20580 28476 20590 28532
rect 25442 28476 25452 28532
rect 25508 28476 26796 28532
rect 26852 28476 26862 28532
rect 7970 28252 7980 28308
rect 8036 28252 8046 28308
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 12898 28140 12908 28196
rect 12964 28140 17836 28196
rect 17892 28140 17902 28196
rect 21634 28140 21644 28196
rect 21700 28140 23996 28196
rect 24052 28140 24668 28196
rect 24724 28140 27468 28196
rect 27524 28140 27534 28196
rect 15092 28028 16268 28084
rect 16324 28028 16334 28084
rect 17602 28028 17612 28084
rect 17668 28028 18508 28084
rect 18564 28028 18574 28084
rect 29250 28028 29260 28084
rect 29316 28028 30156 28084
rect 30212 28028 30716 28084
rect 30772 28028 32844 28084
rect 32900 28028 32910 28084
rect 6178 27916 6188 27972
rect 6244 27916 6636 27972
rect 6692 27916 6702 27972
rect 6962 27804 6972 27860
rect 7028 27804 9884 27860
rect 9940 27804 10556 27860
rect 10612 27804 10622 27860
rect 15092 27748 15148 28028
rect 17714 27916 17724 27972
rect 17780 27916 25564 27972
rect 25620 27916 25630 27972
rect 16370 27804 16380 27860
rect 16436 27804 17388 27860
rect 17444 27804 17454 27860
rect 18610 27804 18620 27860
rect 18676 27804 20076 27860
rect 20132 27804 20142 27860
rect 10098 27692 10108 27748
rect 10164 27692 13468 27748
rect 13524 27692 15148 27748
rect 31490 27692 31500 27748
rect 31556 27692 32508 27748
rect 32564 27692 32574 27748
rect 8082 27580 8092 27636
rect 8148 27580 9548 27636
rect 9604 27580 9614 27636
rect 27458 27468 27468 27524
rect 27524 27468 28028 27524
rect 28084 27468 29260 27524
rect 29316 27468 29326 27524
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 16818 27356 16828 27412
rect 16884 27356 17500 27412
rect 17556 27356 17566 27412
rect 35298 27244 35308 27300
rect 35364 27244 36988 27300
rect 37044 27244 37054 27300
rect 36194 27132 36204 27188
rect 36260 27132 38220 27188
rect 38276 27132 38286 27188
rect 16258 27020 16268 27076
rect 16324 27020 16940 27076
rect 16996 27020 20300 27076
rect 20356 27020 20366 27076
rect 6514 26908 6524 26964
rect 6580 26908 6972 26964
rect 7028 26908 7038 26964
rect 15026 26908 15036 26964
rect 15092 26908 15596 26964
rect 15652 26908 15662 26964
rect 17154 26908 17164 26964
rect 17220 26908 17724 26964
rect 17780 26908 17790 26964
rect 23538 26908 23548 26964
rect 23604 26908 24332 26964
rect 24388 26908 25900 26964
rect 25956 26908 26908 26964
rect 26964 26908 30380 26964
rect 30436 26908 31388 26964
rect 31444 26908 31454 26964
rect 16706 26796 16716 26852
rect 16772 26796 25452 26852
rect 25508 26796 25518 26852
rect 17238 26684 17276 26740
rect 17332 26684 17342 26740
rect 26114 26684 26124 26740
rect 26180 26684 26572 26740
rect 26628 26684 26638 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 16594 26460 16604 26516
rect 16660 26460 17388 26516
rect 17444 26460 17454 26516
rect 22642 26460 22652 26516
rect 22708 26460 23436 26516
rect 23492 26460 23502 26516
rect 25666 26460 25676 26516
rect 25732 26460 26572 26516
rect 26628 26460 26638 26516
rect 22866 26348 22876 26404
rect 22932 26348 23772 26404
rect 23828 26348 23838 26404
rect 26338 26348 26348 26404
rect 26404 26348 27132 26404
rect 27188 26348 27198 26404
rect 14802 26236 14812 26292
rect 14868 26236 15820 26292
rect 15876 26236 15886 26292
rect 24770 26236 24780 26292
rect 24836 26236 25452 26292
rect 25508 26236 26460 26292
rect 26516 26236 26526 26292
rect 4498 26124 4508 26180
rect 4564 26124 5180 26180
rect 5236 26124 5246 26180
rect 22978 26124 22988 26180
rect 23044 26124 24444 26180
rect 24500 26124 24510 26180
rect 25900 26068 25956 26236
rect 3826 26012 3836 26068
rect 3892 26012 4844 26068
rect 4900 26012 4910 26068
rect 15474 26012 15484 26068
rect 15540 26012 16156 26068
rect 16212 26012 16222 26068
rect 17042 26012 17052 26068
rect 17108 26012 17724 26068
rect 17780 26012 17790 26068
rect 25890 26012 25900 26068
rect 25956 26012 25966 26068
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 26348 25676 27804 25732
rect 27860 25676 27870 25732
rect 26348 25620 26404 25676
rect 23090 25564 23100 25620
rect 23156 25564 26348 25620
rect 26404 25564 26414 25620
rect 1932 25452 3948 25508
rect 4004 25452 4014 25508
rect 25106 25452 25116 25508
rect 25172 25452 25676 25508
rect 25732 25452 25742 25508
rect 0 25396 400 25424
rect 1932 25396 1988 25452
rect 0 25340 1988 25396
rect 2594 25340 2604 25396
rect 2660 25340 3724 25396
rect 3780 25340 3790 25396
rect 12674 25340 12684 25396
rect 12740 25340 13244 25396
rect 13300 25340 15484 25396
rect 15540 25340 15550 25396
rect 19058 25340 19068 25396
rect 19124 25340 23100 25396
rect 23156 25340 23166 25396
rect 24210 25340 24220 25396
rect 24276 25340 26124 25396
rect 26180 25340 26190 25396
rect 35410 25340 35420 25396
rect 35476 25340 35868 25396
rect 35924 25340 36764 25396
rect 36820 25340 37548 25396
rect 37604 25340 37614 25396
rect 0 25312 400 25340
rect 4274 25228 4284 25284
rect 4340 25228 5628 25284
rect 5684 25228 5694 25284
rect 19618 25228 19628 25284
rect 19684 25228 23436 25284
rect 23492 25228 23502 25284
rect 26674 25228 26684 25284
rect 26740 25228 27020 25284
rect 27076 25228 27086 25284
rect 27794 25228 27804 25284
rect 27860 25228 30492 25284
rect 30548 25228 31052 25284
rect 31108 25228 31500 25284
rect 31556 25228 31566 25284
rect 39600 25172 40000 25200
rect 13010 25116 13020 25172
rect 13076 25116 13692 25172
rect 13748 25116 13758 25172
rect 26758 25116 26796 25172
rect 26852 25116 26862 25172
rect 30258 25116 30268 25172
rect 30324 25116 31164 25172
rect 31220 25116 31230 25172
rect 38210 25116 38220 25172
rect 38276 25116 40000 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 39600 25088 40000 25116
rect 24098 24892 24108 24948
rect 24164 24892 37884 24948
rect 37940 24892 37950 24948
rect 33394 24780 33404 24836
rect 33460 24780 35084 24836
rect 35140 24780 35150 24836
rect 27010 24668 27020 24724
rect 27076 24668 29708 24724
rect 29764 24668 29774 24724
rect 31490 24668 31500 24724
rect 31556 24668 32060 24724
rect 32116 24668 32126 24724
rect 9986 24556 9996 24612
rect 10052 24556 10332 24612
rect 10388 24556 10398 24612
rect 20738 24556 20748 24612
rect 20804 24556 22092 24612
rect 22148 24556 22158 24612
rect 30818 24556 30828 24612
rect 30884 24556 31388 24612
rect 31444 24556 31454 24612
rect 31826 24332 31836 24388
rect 31892 24332 32620 24388
rect 32676 24332 32686 24388
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 4050 24108 4060 24164
rect 4116 24108 5628 24164
rect 5684 24108 5694 24164
rect 12786 24108 12796 24164
rect 12852 24108 21980 24164
rect 22036 24108 22046 24164
rect 24434 24108 24444 24164
rect 24500 24108 25004 24164
rect 25060 24108 25070 24164
rect 29810 23996 29820 24052
rect 29876 23996 32172 24052
rect 32228 23996 32956 24052
rect 33012 23996 33022 24052
rect 2594 23884 2604 23940
rect 2660 23884 3948 23940
rect 4004 23884 4014 23940
rect 5170 23884 5180 23940
rect 5236 23884 5964 23940
rect 6020 23884 6030 23940
rect 6178 23884 6188 23940
rect 6244 23884 15484 23940
rect 15540 23884 15550 23940
rect 18834 23884 18844 23940
rect 18900 23884 19628 23940
rect 19684 23884 19694 23940
rect 24434 23884 24444 23940
rect 24500 23884 25564 23940
rect 25620 23884 25630 23940
rect 29698 23884 29708 23940
rect 29764 23884 33180 23940
rect 33236 23884 34636 23940
rect 34692 23884 35756 23940
rect 35812 23884 35822 23940
rect 23314 23772 23324 23828
rect 23380 23772 25228 23828
rect 25284 23772 25676 23828
rect 25732 23772 25742 23828
rect 30482 23772 30492 23828
rect 30548 23772 31164 23828
rect 31220 23772 31230 23828
rect 15810 23660 15820 23716
rect 15876 23660 16716 23716
rect 16772 23660 16782 23716
rect 18834 23660 18844 23716
rect 18900 23660 20412 23716
rect 20468 23660 20478 23716
rect 6738 23548 6748 23604
rect 6804 23548 7308 23604
rect 7364 23548 8428 23604
rect 8484 23548 9212 23604
rect 9268 23548 12348 23604
rect 12404 23548 12684 23604
rect 12740 23548 15148 23604
rect 16258 23548 16268 23604
rect 16324 23548 18284 23604
rect 18340 23548 18350 23604
rect 19618 23548 19628 23604
rect 19684 23548 19694 23604
rect 15092 23436 15148 23548
rect 15204 23436 18172 23492
rect 18228 23436 18238 23492
rect 19628 23380 19684 23548
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 25554 23492 25564 23548
rect 25620 23492 25630 23548
rect 23426 23436 23436 23492
rect 23492 23436 24108 23492
rect 24164 23436 24668 23492
rect 24724 23436 24734 23492
rect 25564 23436 29148 23492
rect 29204 23436 29214 23492
rect 34962 23436 34972 23492
rect 35028 23436 36540 23492
rect 36596 23436 36606 23492
rect 5842 23324 5852 23380
rect 5908 23324 6748 23380
rect 6804 23324 6814 23380
rect 9762 23324 9772 23380
rect 9828 23324 10556 23380
rect 10612 23324 18508 23380
rect 18564 23324 19068 23380
rect 19124 23324 19134 23380
rect 19628 23324 20300 23380
rect 20356 23324 20366 23380
rect 27906 23324 27916 23380
rect 27972 23324 29260 23380
rect 29316 23324 29326 23380
rect 19628 23268 19684 23324
rect 15092 23212 16716 23268
rect 16772 23212 17388 23268
rect 17444 23212 17454 23268
rect 17938 23212 17948 23268
rect 18004 23212 19684 23268
rect 28018 23212 28028 23268
rect 28084 23212 28588 23268
rect 28644 23212 28654 23268
rect 15092 23156 15148 23212
rect 5394 23100 5404 23156
rect 5460 23100 6300 23156
rect 6356 23100 6860 23156
rect 6916 23100 8764 23156
rect 8820 23100 11004 23156
rect 11060 23100 11070 23156
rect 13458 23100 13468 23156
rect 13524 23100 15148 23156
rect 34962 23100 34972 23156
rect 35028 23100 35532 23156
rect 35588 23100 35598 23156
rect 4722 22988 4732 23044
rect 4788 22988 5292 23044
rect 5348 22988 5358 23044
rect 12114 22988 12124 23044
rect 12180 22988 12348 23044
rect 12404 22988 16828 23044
rect 16884 22988 17612 23044
rect 17668 22988 18172 23044
rect 18228 22988 18238 23044
rect 25218 22988 25228 23044
rect 25284 22988 26012 23044
rect 26068 22988 26078 23044
rect 34178 22876 34188 22932
rect 34244 22876 35196 22932
rect 35252 22876 35262 22932
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 3332 22540 5068 22596
rect 5124 22540 5852 22596
rect 5908 22540 8652 22596
rect 8708 22540 9772 22596
rect 9828 22540 12796 22596
rect 12852 22540 13804 22596
rect 13860 22540 13870 22596
rect 18498 22540 18508 22596
rect 18564 22540 19964 22596
rect 20020 22540 20030 22596
rect 3332 22372 3388 22540
rect 4610 22428 4620 22484
rect 4676 22428 5628 22484
rect 5684 22428 5694 22484
rect 11442 22428 11452 22484
rect 11508 22428 12348 22484
rect 12404 22428 12414 22484
rect 13122 22428 13132 22484
rect 13188 22428 21532 22484
rect 21588 22428 22204 22484
rect 22260 22428 23324 22484
rect 23380 22428 23390 22484
rect 1810 22316 1820 22372
rect 1876 22316 3388 22372
rect 14914 22316 14924 22372
rect 14980 22316 15148 22372
rect 15204 22316 15214 22372
rect 15474 22316 15484 22372
rect 15540 22316 16156 22372
rect 16212 22316 16222 22372
rect 17378 22316 17388 22372
rect 17444 22316 19180 22372
rect 19236 22316 20412 22372
rect 20468 22316 20478 22372
rect 18498 22204 18508 22260
rect 18564 22204 19628 22260
rect 19684 22204 19694 22260
rect 6290 22092 6300 22148
rect 6356 22092 7308 22148
rect 7364 22092 7374 22148
rect 10994 22092 11004 22148
rect 11060 22092 15708 22148
rect 15764 22092 16828 22148
rect 16884 22092 16894 22148
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 16370 21756 16380 21812
rect 16436 21756 16716 21812
rect 16772 21756 19516 21812
rect 19572 21756 19582 21812
rect 20514 21644 20524 21700
rect 20580 21644 21532 21700
rect 21588 21644 21980 21700
rect 22036 21644 22046 21700
rect 10882 21532 10892 21588
rect 10948 21532 13468 21588
rect 13524 21532 14140 21588
rect 14196 21532 14206 21588
rect 32498 21532 32508 21588
rect 32564 21532 34524 21588
rect 34580 21532 37772 21588
rect 37828 21532 37838 21588
rect 4386 21420 4396 21476
rect 4452 21420 5852 21476
rect 5908 21420 5918 21476
rect 17378 21420 17388 21476
rect 17444 21420 17724 21476
rect 17780 21420 17790 21476
rect 22418 21420 22428 21476
rect 22484 21420 29596 21476
rect 29652 21420 29662 21476
rect 36082 21420 36092 21476
rect 36148 21420 36988 21476
rect 37044 21420 37054 21476
rect 31826 21308 31836 21364
rect 31892 21308 33068 21364
rect 33124 21308 33134 21364
rect 13682 21196 13692 21252
rect 13748 21196 15484 21252
rect 15540 21196 15550 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 7410 21084 7420 21140
rect 7476 21084 8204 21140
rect 8260 21084 8270 21140
rect 12002 20860 12012 20916
rect 12068 20860 13692 20916
rect 13748 20860 13758 20916
rect 5058 20748 5068 20804
rect 5124 20748 5964 20804
rect 6020 20748 7420 20804
rect 7476 20748 13132 20804
rect 13188 20748 13198 20804
rect 17378 20748 17388 20804
rect 17444 20748 18284 20804
rect 18340 20748 18350 20804
rect 26674 20524 26684 20580
rect 26740 20524 27244 20580
rect 27300 20524 29260 20580
rect 29316 20524 32732 20580
rect 32788 20524 33404 20580
rect 33460 20524 34860 20580
rect 34916 20524 34926 20580
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 6290 20188 6300 20244
rect 6356 20188 8092 20244
rect 8148 20188 8652 20244
rect 8708 20188 11116 20244
rect 11172 20188 11182 20244
rect 34178 20188 34188 20244
rect 34244 20188 34972 20244
rect 35028 20188 35038 20244
rect 34626 20076 34636 20132
rect 34692 20076 36316 20132
rect 36372 20076 36382 20132
rect 21186 19964 21196 20020
rect 21252 19964 23324 20020
rect 23380 19964 23884 20020
rect 23940 19964 26684 20020
rect 26740 19964 26750 20020
rect 33730 19964 33740 20020
rect 33796 19964 34076 20020
rect 34132 19964 34524 20020
rect 34580 19964 34590 20020
rect 34738 19964 34748 20020
rect 34804 19964 35532 20020
rect 35588 19964 35598 20020
rect 33618 19852 33628 19908
rect 33684 19852 35308 19908
rect 35364 19852 35374 19908
rect 11106 19740 11116 19796
rect 11172 19740 11788 19796
rect 11844 19740 12124 19796
rect 12180 19740 12190 19796
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 4162 19404 4172 19460
rect 4228 19404 4956 19460
rect 5012 19404 5022 19460
rect 22754 19404 22764 19460
rect 22820 19404 29708 19460
rect 29764 19404 30492 19460
rect 30548 19404 32844 19460
rect 32900 19404 33628 19460
rect 33684 19404 33694 19460
rect 34850 19404 34860 19460
rect 34916 19404 35756 19460
rect 35812 19404 35822 19460
rect 14242 19292 14252 19348
rect 14308 19292 17276 19348
rect 17332 19292 17342 19348
rect 29250 19292 29260 19348
rect 29316 19292 30828 19348
rect 30884 19292 32396 19348
rect 32452 19292 33292 19348
rect 33348 19292 34076 19348
rect 34132 19292 34142 19348
rect 13458 19180 13468 19236
rect 13524 19180 16828 19236
rect 16884 19180 16894 19236
rect 17042 19180 17052 19236
rect 17108 19180 17332 19236
rect 26674 19180 26684 19236
rect 26740 19180 27132 19236
rect 27188 19180 27198 19236
rect 17276 19124 17332 19180
rect 17266 19068 17276 19124
rect 17332 19068 17342 19124
rect 35186 18956 35196 19012
rect 35252 18956 36988 19012
rect 37044 18956 37054 19012
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 21074 18732 21084 18788
rect 21140 18732 31052 18788
rect 31108 18732 34300 18788
rect 34356 18732 34860 18788
rect 34916 18732 34926 18788
rect 20066 18620 20076 18676
rect 20132 18620 20636 18676
rect 20692 18620 20702 18676
rect 5058 18508 5068 18564
rect 5124 18508 5852 18564
rect 5908 18508 5918 18564
rect 34962 18508 34972 18564
rect 35028 18508 35756 18564
rect 35812 18508 35822 18564
rect 9314 18396 9324 18452
rect 9380 18396 10220 18452
rect 10276 18396 10286 18452
rect 18946 18396 18956 18452
rect 19012 18396 19964 18452
rect 20020 18396 20412 18452
rect 20468 18396 20478 18452
rect 34626 18396 34636 18452
rect 34692 18396 35980 18452
rect 36036 18396 36046 18452
rect 2594 18284 2604 18340
rect 2660 18284 5516 18340
rect 5572 18284 5582 18340
rect 15362 18284 15372 18340
rect 15428 18284 19740 18340
rect 19796 18284 19806 18340
rect 30482 18284 30492 18340
rect 30548 18284 30828 18340
rect 30884 18284 30894 18340
rect 31378 18284 31388 18340
rect 31444 18284 32060 18340
rect 32116 18284 32126 18340
rect 36642 18284 36652 18340
rect 36708 18284 37436 18340
rect 37492 18284 37502 18340
rect 16930 18172 16940 18228
rect 16996 18172 18060 18228
rect 18116 18172 18126 18228
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 16930 17948 16940 18004
rect 16996 17948 17388 18004
rect 17444 17948 17454 18004
rect 23986 17724 23996 17780
rect 24052 17724 25564 17780
rect 25620 17724 25630 17780
rect 27682 17724 27692 17780
rect 27748 17724 28588 17780
rect 28644 17724 29260 17780
rect 29316 17724 30044 17780
rect 30100 17724 30492 17780
rect 30548 17724 32508 17780
rect 32564 17724 32574 17780
rect 33282 17724 33292 17780
rect 33348 17724 34188 17780
rect 34244 17724 34254 17780
rect 20738 17612 20748 17668
rect 20804 17612 22652 17668
rect 22708 17612 22718 17668
rect 33170 17612 33180 17668
rect 33236 17612 35084 17668
rect 35140 17612 38108 17668
rect 38164 17612 38174 17668
rect 11778 17500 11788 17556
rect 11844 17500 13356 17556
rect 13412 17500 13422 17556
rect 12562 17388 12572 17444
rect 12628 17388 13468 17444
rect 13524 17388 13534 17444
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 5506 17052 5516 17108
rect 5572 17052 8652 17108
rect 8708 17052 10780 17108
rect 10836 17052 10846 17108
rect 16258 17052 16268 17108
rect 16324 17052 16940 17108
rect 16996 17052 17500 17108
rect 17556 17052 17566 17108
rect 26226 17052 26236 17108
rect 26292 17052 26908 17108
rect 26964 17052 30268 17108
rect 30324 17052 30334 17108
rect 32498 17052 32508 17108
rect 32564 17052 33180 17108
rect 33236 17052 33246 17108
rect 16706 16940 16716 16996
rect 16772 16940 17612 16996
rect 17668 16940 17948 16996
rect 18004 16940 18014 16996
rect 22642 16940 22652 16996
rect 22708 16940 23100 16996
rect 23156 16940 26684 16996
rect 26740 16940 27692 16996
rect 27748 16940 27758 16996
rect 14690 16828 14700 16884
rect 14756 16828 15596 16884
rect 15652 16828 15662 16884
rect 7522 16716 7532 16772
rect 7588 16716 12236 16772
rect 12292 16716 12302 16772
rect 16370 16716 16380 16772
rect 16436 16716 17388 16772
rect 17444 16716 17454 16772
rect 18722 16716 18732 16772
rect 18788 16716 19068 16772
rect 19124 16716 19134 16772
rect 25666 16716 25676 16772
rect 25732 16716 26796 16772
rect 26852 16716 28700 16772
rect 28756 16716 28766 16772
rect 14690 16492 14700 16548
rect 14756 16492 16156 16548
rect 16212 16492 16222 16548
rect 18274 16492 18284 16548
rect 18340 16492 19068 16548
rect 19124 16492 19134 16548
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 17826 16268 17836 16324
rect 17892 16268 19628 16324
rect 19684 16268 19694 16324
rect 21634 16268 21644 16324
rect 21700 16268 22092 16324
rect 22148 16268 22876 16324
rect 22932 16268 22942 16324
rect 10210 16156 10220 16212
rect 10276 16156 12124 16212
rect 12180 16156 12908 16212
rect 12964 16156 13804 16212
rect 13860 16156 15148 16212
rect 19730 16156 19740 16212
rect 19796 16156 21868 16212
rect 21924 16156 21934 16212
rect 30706 16156 30716 16212
rect 30772 16156 31052 16212
rect 31108 16156 31118 16212
rect 12002 16044 12012 16100
rect 12068 16044 14476 16100
rect 14532 16044 14542 16100
rect 15092 16044 15148 16156
rect 15204 16044 15214 16100
rect 20514 16044 20524 16100
rect 20580 16044 21420 16100
rect 21476 16044 21486 16100
rect 28690 16044 28700 16100
rect 28756 16044 29708 16100
rect 29764 16044 29774 16100
rect 34626 16044 34636 16100
rect 34692 16044 35196 16100
rect 35252 16044 35262 16100
rect 7074 15932 7084 15988
rect 7140 15932 7980 15988
rect 8036 15932 11788 15988
rect 11844 15932 11854 15988
rect 14242 15932 14252 15988
rect 14308 15932 19404 15988
rect 19460 15932 19470 15988
rect 11442 15820 11452 15876
rect 11508 15820 12236 15876
rect 12292 15820 12302 15876
rect 20402 15820 20412 15876
rect 20468 15820 28028 15876
rect 28084 15820 28094 15876
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 12674 15596 12684 15652
rect 12740 15596 15820 15652
rect 15876 15596 18956 15652
rect 19012 15596 19292 15652
rect 19348 15596 19358 15652
rect 0 15540 400 15568
rect 0 15484 8092 15540
rect 8148 15484 8158 15540
rect 8978 15484 8988 15540
rect 9044 15484 10220 15540
rect 10276 15484 10286 15540
rect 16482 15484 16492 15540
rect 16548 15484 18732 15540
rect 18788 15484 18798 15540
rect 23874 15484 23884 15540
rect 23940 15484 26012 15540
rect 26068 15484 26078 15540
rect 0 15456 400 15484
rect 12114 15372 12124 15428
rect 12180 15372 17836 15428
rect 17892 15372 17902 15428
rect 19282 15372 19292 15428
rect 19348 15372 20300 15428
rect 20356 15372 20366 15428
rect 24210 15372 24220 15428
rect 24276 15372 25340 15428
rect 25396 15372 26460 15428
rect 26516 15372 26526 15428
rect 6850 15260 6860 15316
rect 6916 15260 7532 15316
rect 7588 15260 7598 15316
rect 10434 15260 10444 15316
rect 10500 15260 11452 15316
rect 11508 15260 11518 15316
rect 11666 15260 11676 15316
rect 11732 15260 13132 15316
rect 13188 15260 14924 15316
rect 14980 15260 16492 15316
rect 16548 15260 16558 15316
rect 18162 15260 18172 15316
rect 18228 15260 24108 15316
rect 24164 15260 24174 15316
rect 30930 15260 30940 15316
rect 30996 15260 31836 15316
rect 31892 15260 31902 15316
rect 14578 15148 14588 15204
rect 14644 15148 16044 15204
rect 16100 15148 16110 15204
rect 18274 15148 18284 15204
rect 18340 15148 19404 15204
rect 19460 15148 19470 15204
rect 20850 15148 20860 15204
rect 20916 15148 21868 15204
rect 21924 15148 21934 15204
rect 31164 15148 34636 15204
rect 34692 15148 34702 15204
rect 18946 15036 18956 15092
rect 19012 15036 19180 15092
rect 19236 15036 19740 15092
rect 19796 15036 19806 15092
rect 31164 14980 31220 15148
rect 26450 14924 26460 14980
rect 26516 14924 27020 14980
rect 27076 14924 29484 14980
rect 29540 14924 30604 14980
rect 30660 14924 31220 14980
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 30594 14588 30604 14644
rect 30660 14588 31164 14644
rect 31220 14588 31230 14644
rect 21858 14476 21868 14532
rect 21924 14476 22764 14532
rect 22820 14476 22830 14532
rect 14466 14252 14476 14308
rect 14532 14252 15148 14308
rect 15204 14252 15214 14308
rect 31490 14252 31500 14308
rect 31556 14252 33292 14308
rect 33348 14252 33358 14308
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 8306 13804 8316 13860
rect 8372 13804 9548 13860
rect 9604 13804 9614 13860
rect 4722 13692 4732 13748
rect 4788 13692 7644 13748
rect 7700 13692 7980 13748
rect 8036 13692 8046 13748
rect 15138 13580 15148 13636
rect 15204 13580 17948 13636
rect 18004 13580 18620 13636
rect 18676 13580 18686 13636
rect 29026 13580 29036 13636
rect 29092 13580 30044 13636
rect 30100 13580 31500 13636
rect 31556 13580 31948 13636
rect 32004 13580 32014 13636
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 18610 13132 18620 13188
rect 18676 13132 24556 13188
rect 24612 13132 25228 13188
rect 25284 13132 30156 13188
rect 30212 13132 31164 13188
rect 31220 13132 31230 13188
rect 16146 13020 16156 13076
rect 16212 13020 17052 13076
rect 17108 13020 18284 13076
rect 18340 13020 18844 13076
rect 18900 13020 18910 13076
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 16594 12460 16604 12516
rect 16660 12460 17388 12516
rect 17444 12460 17454 12516
rect 6962 12348 6972 12404
rect 7028 12348 8092 12404
rect 8148 12348 9884 12404
rect 9940 12348 9950 12404
rect 11330 12348 11340 12404
rect 11396 12348 12236 12404
rect 12292 12348 13804 12404
rect 13860 12348 13870 12404
rect 15474 12348 15484 12404
rect 15540 12348 15932 12404
rect 15988 12348 16492 12404
rect 16548 12348 18956 12404
rect 19012 12348 19022 12404
rect 19170 12348 19180 12404
rect 19236 12348 19274 12404
rect 12002 12236 12012 12292
rect 12068 12236 13356 12292
rect 13412 12236 13422 12292
rect 19030 12236 19068 12292
rect 19124 12236 19134 12292
rect 23762 12236 23772 12292
rect 23828 12236 24220 12292
rect 24276 12236 25116 12292
rect 25172 12236 26908 12292
rect 26852 12180 26908 12236
rect 14354 12124 14364 12180
rect 14420 12124 14812 12180
rect 14868 12124 15932 12180
rect 15988 12124 15998 12180
rect 16258 12124 16268 12180
rect 16324 12124 17500 12180
rect 17556 12124 17566 12180
rect 18050 12124 18060 12180
rect 18116 12124 25228 12180
rect 25284 12124 25294 12180
rect 26852 12124 28588 12180
rect 28644 12124 29708 12180
rect 29764 12124 29774 12180
rect 4834 12012 4844 12068
rect 4900 12012 7644 12068
rect 7700 12012 8428 12068
rect 8484 12012 8494 12068
rect 8978 12012 8988 12068
rect 9044 12012 20188 12068
rect 20244 12012 20254 12068
rect 28018 12012 28028 12068
rect 28084 12012 28924 12068
rect 28980 12012 28990 12068
rect 17378 11900 17388 11956
rect 17444 11900 17836 11956
rect 17892 11900 18788 11956
rect 18946 11900 18956 11956
rect 19012 11900 19628 11956
rect 19684 11900 19694 11956
rect 18732 11844 18788 11900
rect 10994 11788 11004 11844
rect 11060 11788 17948 11844
rect 18004 11788 18014 11844
rect 18732 11788 19292 11844
rect 19348 11788 19740 11844
rect 19796 11788 19806 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 5730 11676 5740 11732
rect 5796 11676 7532 11732
rect 7588 11676 8988 11732
rect 9044 11676 10780 11732
rect 10836 11676 11676 11732
rect 11732 11676 12124 11732
rect 12180 11676 12190 11732
rect 19170 11676 19180 11732
rect 19236 11676 20244 11732
rect 20402 11676 20412 11732
rect 20468 11676 21196 11732
rect 21252 11676 21262 11732
rect 20188 11620 20244 11676
rect 12338 11564 12348 11620
rect 12404 11564 19740 11620
rect 19796 11564 19806 11620
rect 20150 11564 20188 11620
rect 20244 11564 20748 11620
rect 20804 11564 21756 11620
rect 21812 11564 21822 11620
rect 11778 11452 11788 11508
rect 11844 11452 12908 11508
rect 12964 11452 12974 11508
rect 17826 11452 17836 11508
rect 17892 11452 19852 11508
rect 19908 11452 19918 11508
rect 26226 11452 26236 11508
rect 26292 11452 30268 11508
rect 30324 11452 30334 11508
rect 20178 11340 20188 11396
rect 20244 11340 21420 11396
rect 21476 11340 21486 11396
rect 15698 11228 15708 11284
rect 15764 11228 16604 11284
rect 16660 11228 16670 11284
rect 19954 11228 19964 11284
rect 20020 11228 26796 11284
rect 26852 11228 26862 11284
rect 31378 11228 31388 11284
rect 31444 11228 32396 11284
rect 32452 11228 32462 11284
rect 12114 11116 12124 11172
rect 12180 11116 12460 11172
rect 12516 11116 13356 11172
rect 13412 11116 13422 11172
rect 14466 11116 14476 11172
rect 14532 11116 15148 11172
rect 15204 11116 15214 11172
rect 20514 11116 20524 11172
rect 20580 11116 21196 11172
rect 21252 11116 21262 11172
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 10770 10780 10780 10836
rect 10836 10780 11788 10836
rect 11844 10780 11854 10836
rect 15810 10780 15820 10836
rect 15876 10780 16156 10836
rect 16212 10780 16604 10836
rect 16660 10780 16670 10836
rect 17686 10780 17724 10836
rect 17780 10780 17790 10836
rect 18274 10780 18284 10836
rect 18340 10780 20636 10836
rect 20692 10780 20702 10836
rect 24210 10780 24220 10836
rect 24276 10780 25340 10836
rect 25396 10780 26348 10836
rect 26404 10780 26414 10836
rect 10098 10668 10108 10724
rect 10164 10668 10668 10724
rect 10724 10668 10734 10724
rect 19058 10668 19068 10724
rect 19124 10668 19740 10724
rect 19796 10668 19806 10724
rect 7186 10556 7196 10612
rect 7252 10556 10220 10612
rect 10276 10556 10286 10612
rect 10994 10556 11004 10612
rect 11060 10556 18508 10612
rect 18564 10556 18574 10612
rect 19058 10556 19068 10612
rect 19124 10556 19180 10612
rect 19236 10556 19246 10612
rect 19618 10556 19628 10612
rect 19684 10556 20524 10612
rect 20580 10556 20590 10612
rect 24658 10556 24668 10612
rect 24724 10556 25676 10612
rect 25732 10556 26012 10612
rect 26068 10556 26908 10612
rect 26964 10556 27468 10612
rect 27524 10556 27534 10612
rect 15810 10444 15820 10500
rect 15876 10444 16828 10500
rect 16884 10444 17500 10500
rect 17556 10444 17566 10500
rect 18946 10444 18956 10500
rect 19012 10444 19852 10500
rect 19908 10444 20188 10500
rect 20244 10444 20254 10500
rect 8530 10332 8540 10388
rect 8596 10332 9996 10388
rect 10052 10332 10444 10388
rect 10500 10332 10510 10388
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 19282 10108 19292 10164
rect 19348 10108 21868 10164
rect 21924 10108 21934 10164
rect 17686 9996 17724 10052
rect 17780 9996 17790 10052
rect 26338 9996 26348 10052
rect 26404 9996 27916 10052
rect 27972 9996 27982 10052
rect 4722 9884 4732 9940
rect 4788 9884 5516 9940
rect 5572 9884 5582 9940
rect 10658 9884 10668 9940
rect 10724 9884 11564 9940
rect 11620 9884 11630 9940
rect 16370 9884 16380 9940
rect 16436 9884 17164 9940
rect 17220 9884 17230 9940
rect 18610 9884 18620 9940
rect 18676 9884 26460 9940
rect 26516 9884 26526 9940
rect 26674 9884 26684 9940
rect 26740 9884 29148 9940
rect 29204 9884 31724 9940
rect 31780 9884 31790 9940
rect 17490 9772 17500 9828
rect 17556 9772 18396 9828
rect 18452 9772 26908 9828
rect 31490 9772 31500 9828
rect 31556 9772 32172 9828
rect 32228 9772 32238 9828
rect 26852 9716 26908 9772
rect 5058 9660 5068 9716
rect 5124 9660 7084 9716
rect 7140 9660 7150 9716
rect 26852 9660 29708 9716
rect 29764 9660 30828 9716
rect 30884 9660 37212 9716
rect 37268 9660 37278 9716
rect 17378 9548 17388 9604
rect 17444 9548 18172 9604
rect 18228 9548 18238 9604
rect 19954 9548 19964 9604
rect 20020 9548 21756 9604
rect 21812 9548 21822 9604
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 4274 9212 4284 9268
rect 4340 9212 8988 9268
rect 9044 9212 9884 9268
rect 9940 9212 10780 9268
rect 10836 9212 10846 9268
rect 16594 8764 16604 8820
rect 16660 8764 19740 8820
rect 19796 8764 19806 8820
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 39600 8596 40000 8624
rect 38322 8540 38332 8596
rect 38388 8540 40000 8596
rect 39600 8512 40000 8540
rect 25442 8428 25452 8484
rect 25508 8428 28700 8484
rect 28756 8428 29932 8484
rect 29988 8428 30156 8484
rect 30212 8428 31948 8484
rect 32004 8428 32014 8484
rect 27244 8260 27300 8428
rect 25554 8204 25564 8260
rect 25620 8204 27020 8260
rect 27076 8204 27086 8260
rect 27234 8204 27244 8260
rect 27300 8204 27310 8260
rect 15922 7980 15932 8036
rect 15988 7980 16604 8036
rect 16660 7980 16670 8036
rect 25106 7980 25116 8036
rect 25172 7980 26348 8036
rect 26404 7980 31276 8036
rect 31332 7980 31948 8036
rect 32004 7980 32014 8036
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 10658 7644 10668 7700
rect 10724 7644 11116 7700
rect 11172 7644 13468 7700
rect 13524 7644 14476 7700
rect 14532 7644 14542 7700
rect 30034 7644 30044 7700
rect 30100 7644 31388 7700
rect 31444 7644 31454 7700
rect 26898 7532 26908 7588
rect 26964 7532 27692 7588
rect 27748 7532 27758 7588
rect 6626 7308 6636 7364
rect 6692 7308 15148 7364
rect 19058 7308 19068 7364
rect 19124 7308 20412 7364
rect 20468 7308 20478 7364
rect 26562 7308 26572 7364
rect 26628 7308 30156 7364
rect 30212 7308 31500 7364
rect 31556 7308 31566 7364
rect 15092 7252 15148 7308
rect 5954 7196 5964 7252
rect 6020 7196 7420 7252
rect 7476 7196 8652 7252
rect 8708 7196 8718 7252
rect 15092 7196 15708 7252
rect 15764 7196 15774 7252
rect 8978 7084 8988 7140
rect 9044 7084 10332 7140
rect 10388 7084 10398 7140
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 10434 6860 10444 6916
rect 10500 6860 10780 6916
rect 10836 6860 11452 6916
rect 11508 6860 12124 6916
rect 12180 6860 13692 6916
rect 13748 6860 14364 6916
rect 14420 6860 14430 6916
rect 10098 6748 10108 6804
rect 10164 6748 10892 6804
rect 10948 6748 10958 6804
rect 14364 6692 14420 6860
rect 9986 6636 9996 6692
rect 10052 6636 10444 6692
rect 10500 6636 10510 6692
rect 14364 6636 15148 6692
rect 15204 6636 15214 6692
rect 16370 6636 16380 6692
rect 16436 6636 18284 6692
rect 18340 6636 18350 6692
rect 20402 6636 20412 6692
rect 20468 6636 21308 6692
rect 21364 6636 21374 6692
rect 25554 6636 25564 6692
rect 25620 6636 27356 6692
rect 27412 6636 27422 6692
rect 7298 6524 7308 6580
rect 7364 6524 9660 6580
rect 9716 6524 10668 6580
rect 10724 6524 10734 6580
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 13010 6076 13020 6132
rect 13076 6076 16268 6132
rect 16324 6076 16334 6132
rect 18946 5852 18956 5908
rect 19012 5852 22316 5908
rect 22372 5852 22382 5908
rect 23202 5852 23212 5908
rect 23268 5852 24220 5908
rect 24276 5852 24892 5908
rect 24948 5852 25564 5908
rect 25620 5852 25630 5908
rect 0 5684 400 5712
rect 0 5628 532 5684
rect 0 5600 400 5628
rect 476 5460 532 5628
rect 8642 5516 8652 5572
rect 8708 5516 9324 5572
rect 9380 5516 22204 5572
rect 22260 5516 22270 5572
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 252 5404 532 5460
rect 21532 5404 23100 5460
rect 23156 5404 25116 5460
rect 25172 5404 25182 5460
rect 27346 5404 27356 5460
rect 27412 5404 27422 5460
rect 252 5124 308 5404
rect 21532 5348 21588 5404
rect 20178 5292 20188 5348
rect 20244 5292 21532 5348
rect 21588 5292 21598 5348
rect 22306 5292 22316 5348
rect 22372 5292 22382 5348
rect 22316 5236 22372 5292
rect 27356 5236 27412 5404
rect 5282 5180 5292 5236
rect 5348 5180 6412 5236
rect 6468 5180 19740 5236
rect 19796 5180 20412 5236
rect 20468 5180 20478 5236
rect 22316 5180 23324 5236
rect 23380 5180 24220 5236
rect 24276 5180 26572 5236
rect 26628 5180 27692 5236
rect 27748 5180 27758 5236
rect 252 5068 3388 5124
rect 14914 5068 14924 5124
rect 14980 5068 15540 5124
rect 15698 5068 15708 5124
rect 15764 5068 16828 5124
rect 16884 5068 17724 5124
rect 17780 5068 17790 5124
rect 24434 5068 24444 5124
rect 24500 5068 25228 5124
rect 25284 5068 25294 5124
rect 3332 4900 3388 5068
rect 15484 5012 15540 5068
rect 15484 4956 16380 5012
rect 16436 4956 16446 5012
rect 3332 4844 5628 4900
rect 5684 4844 5694 4900
rect 19506 4844 19516 4900
rect 19572 4844 20076 4900
rect 20132 4844 20142 4900
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 8082 4508 8092 4564
rect 8148 4508 9772 4564
rect 9828 4508 10780 4564
rect 10836 4508 10846 4564
rect 12898 4396 12908 4452
rect 12964 4396 14140 4452
rect 14196 4396 14206 4452
rect 15092 4396 25228 4452
rect 25284 4396 25294 4452
rect 15092 4340 15148 4396
rect 10098 4284 10108 4340
rect 10164 4284 10556 4340
rect 10612 4284 10622 4340
rect 14018 4284 14028 4340
rect 14084 4284 15148 4340
rect 14476 4228 14532 4284
rect 14466 4172 14476 4228
rect 14532 4172 14542 4228
rect 8194 4060 8204 4116
rect 8260 4060 10556 4116
rect 10612 4060 10622 4116
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 7522 3500 7532 3556
rect 7588 3500 8316 3556
rect 8372 3500 8382 3556
rect 8754 3500 8764 3556
rect 8820 3500 10332 3556
rect 10388 3500 10398 3556
rect 6290 3388 6300 3444
rect 6356 3388 7420 3444
rect 7476 3388 7486 3444
rect 9090 3388 9100 3444
rect 9156 3388 10052 3444
rect 17826 3388 17836 3444
rect 17892 3388 18620 3444
rect 18676 3388 18686 3444
rect 32498 3388 32508 3444
rect 32564 3388 33628 3444
rect 33684 3388 33694 3444
rect 9996 3332 10052 3388
rect 9986 3276 9996 3332
rect 10052 3276 10062 3332
rect 11106 3276 11116 3332
rect 11172 3276 13468 3332
rect 13524 3276 13534 3332
rect 15138 3276 15148 3332
rect 15204 3276 16156 3332
rect 16212 3276 16222 3332
rect 25554 3276 25564 3332
rect 25620 3276 27020 3332
rect 27076 3276 27086 3332
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 34738 3052 34748 3108
rect 34804 3052 36652 3108
rect 36708 3052 36718 3108
rect 16370 2940 16380 2996
rect 16436 2940 19852 2996
rect 19908 2940 19918 2996
rect 34402 2940 34412 2996
rect 34468 2940 35980 2996
rect 36036 2940 36046 2996
rect 10882 2828 10892 2884
rect 10948 2828 11564 2884
rect 11620 2828 11630 2884
rect 14242 2828 14252 2884
rect 14308 2828 15260 2884
rect 15316 2828 15326 2884
rect 21410 2828 21420 2884
rect 21476 2828 22316 2884
rect 22372 2828 22382 2884
rect 25778 2828 25788 2884
rect 25844 2828 26796 2884
rect 26852 2828 26862 2884
rect 11890 2716 11900 2772
rect 11956 2716 12684 2772
rect 12740 2716 12750 2772
rect 16370 2716 16380 2772
rect 16436 2716 17612 2772
rect 17668 2716 18172 2772
rect 18228 2716 18238 2772
rect 23202 2716 23212 2772
rect 23268 2716 25228 2772
rect 25284 2716 25294 2772
rect 9762 2604 9772 2660
rect 9828 2604 10444 2660
rect 10500 2604 10510 2660
rect 11106 2604 11116 2660
rect 11172 2604 12908 2660
rect 12964 2604 20188 2660
rect 26562 2604 26572 2660
rect 26628 2604 27356 2660
rect 27412 2604 27422 2660
rect 34850 2604 34860 2660
rect 34916 2604 36092 2660
rect 36148 2604 36158 2660
rect 20132 2548 20188 2604
rect 10546 2492 10556 2548
rect 10612 2492 14476 2548
rect 14532 2492 14542 2548
rect 20132 2492 33180 2548
rect 33236 2492 33246 2548
rect 4466 2324 4476 2380
rect 4532 2324 4580 2380
rect 4636 2324 4684 2380
rect 4740 2324 4750 2380
rect 35186 2324 35196 2380
rect 35252 2324 35300 2380
rect 35356 2324 35404 2380
rect 35460 2324 35470 2380
rect 11554 2156 11564 2212
rect 11620 2156 13244 2212
rect 13300 2156 13310 2212
rect 21970 1932 21980 1988
rect 22036 1932 23660 1988
rect 23716 1932 23726 1988
rect 33730 1932 33740 1988
rect 33796 1932 35308 1988
rect 35364 1932 35374 1988
rect 3826 1820 3836 1876
rect 3892 1820 5852 1876
rect 5908 1820 5918 1876
rect 35186 1820 35196 1876
rect 35252 1820 36204 1876
rect 36260 1820 36270 1876
rect 5058 1708 5068 1764
rect 5124 1708 6748 1764
rect 6804 1708 6814 1764
rect 17266 1708 17276 1764
rect 17332 1708 18172 1764
rect 18228 1708 18238 1764
rect 27906 1708 27916 1764
rect 27972 1708 29148 1764
rect 29204 1708 29214 1764
rect 36082 1708 36092 1764
rect 36148 1708 36876 1764
rect 36932 1708 37436 1764
rect 37492 1708 37502 1764
rect 19826 1540 19836 1596
rect 19892 1540 19940 1596
rect 19996 1540 20044 1596
rect 20100 1540 20110 1596
<< via3 >>
rect 4476 97972 4532 98028
rect 4580 97972 4636 98028
rect 4684 97972 4740 98028
rect 35196 97972 35252 98028
rect 35300 97972 35356 98028
rect 35404 97972 35460 98028
rect 19836 97188 19892 97244
rect 19940 97188 19996 97244
rect 20044 97188 20100 97244
rect 4476 96404 4532 96460
rect 4580 96404 4636 96460
rect 4684 96404 4740 96460
rect 35196 96404 35252 96460
rect 35300 96404 35356 96460
rect 35404 96404 35460 96460
rect 19836 95620 19892 95676
rect 19940 95620 19996 95676
rect 20044 95620 20100 95676
rect 25116 95452 25172 95508
rect 4476 94836 4532 94892
rect 4580 94836 4636 94892
rect 4684 94836 4740 94892
rect 35196 94836 35252 94892
rect 35300 94836 35356 94892
rect 35404 94836 35460 94892
rect 19836 94052 19892 94108
rect 19940 94052 19996 94108
rect 20044 94052 20100 94108
rect 24444 93436 24500 93492
rect 4476 93268 4532 93324
rect 4580 93268 4636 93324
rect 4684 93268 4740 93324
rect 35196 93268 35252 93324
rect 35300 93268 35356 93324
rect 35404 93268 35460 93324
rect 19836 92484 19892 92540
rect 19940 92484 19996 92540
rect 20044 92484 20100 92540
rect 4476 91700 4532 91756
rect 4580 91700 4636 91756
rect 4684 91700 4740 91756
rect 35196 91700 35252 91756
rect 35300 91700 35356 91756
rect 35404 91700 35460 91756
rect 19836 90916 19892 90972
rect 19940 90916 19996 90972
rect 20044 90916 20100 90972
rect 24556 90636 24612 90692
rect 4476 90132 4532 90188
rect 4580 90132 4636 90188
rect 4684 90132 4740 90188
rect 35196 90132 35252 90188
rect 35300 90132 35356 90188
rect 35404 90132 35460 90188
rect 24556 89740 24612 89796
rect 27468 89516 27524 89572
rect 19836 89348 19892 89404
rect 19940 89348 19996 89404
rect 20044 89348 20100 89404
rect 4476 88564 4532 88620
rect 4580 88564 4636 88620
rect 4684 88564 4740 88620
rect 35196 88564 35252 88620
rect 35300 88564 35356 88620
rect 35404 88564 35460 88620
rect 19836 87780 19892 87836
rect 19940 87780 19996 87836
rect 20044 87780 20100 87836
rect 24556 87500 24612 87556
rect 4476 86996 4532 87052
rect 4580 86996 4636 87052
rect 4684 86996 4740 87052
rect 35196 86996 35252 87052
rect 35300 86996 35356 87052
rect 35404 86996 35460 87052
rect 24444 86828 24500 86884
rect 26012 86604 26068 86660
rect 19836 86212 19892 86268
rect 19940 86212 19996 86268
rect 20044 86212 20100 86268
rect 4476 85428 4532 85484
rect 4580 85428 4636 85484
rect 4684 85428 4740 85484
rect 35196 85428 35252 85484
rect 35300 85428 35356 85484
rect 35404 85428 35460 85484
rect 19836 84644 19892 84700
rect 19940 84644 19996 84700
rect 20044 84644 20100 84700
rect 25116 84140 25172 84196
rect 27356 84140 27412 84196
rect 4476 83860 4532 83916
rect 4580 83860 4636 83916
rect 4684 83860 4740 83916
rect 35196 83860 35252 83916
rect 35300 83860 35356 83916
rect 35404 83860 35460 83916
rect 26012 83244 26068 83300
rect 19836 83076 19892 83132
rect 19940 83076 19996 83132
rect 20044 83076 20100 83132
rect 27244 82348 27300 82404
rect 4476 82292 4532 82348
rect 4580 82292 4636 82348
rect 4684 82292 4740 82348
rect 35196 82292 35252 82348
rect 35300 82292 35356 82348
rect 35404 82292 35460 82348
rect 35644 81676 35700 81732
rect 19836 81508 19892 81564
rect 19940 81508 19996 81564
rect 20044 81508 20100 81564
rect 27356 81340 27412 81396
rect 4476 80724 4532 80780
rect 4580 80724 4636 80780
rect 4684 80724 4740 80780
rect 35196 80724 35252 80780
rect 35300 80724 35356 80780
rect 35404 80724 35460 80780
rect 34188 80668 34244 80724
rect 19836 79940 19892 79996
rect 19940 79940 19996 79996
rect 20044 79940 20100 79996
rect 30492 79212 30548 79268
rect 4476 79156 4532 79212
rect 4580 79156 4636 79212
rect 4684 79156 4740 79212
rect 35196 79156 35252 79212
rect 35300 79156 35356 79212
rect 35404 79156 35460 79212
rect 27020 79100 27076 79156
rect 27580 78988 27636 79044
rect 26908 78876 26964 78932
rect 26012 78652 26068 78708
rect 19836 78372 19892 78428
rect 19940 78372 19996 78428
rect 20044 78372 20100 78428
rect 25788 78092 25844 78148
rect 26124 78092 26180 78148
rect 25788 77868 25844 77924
rect 4476 77588 4532 77644
rect 4580 77588 4636 77644
rect 4684 77588 4740 77644
rect 35196 77588 35252 77644
rect 35300 77588 35356 77644
rect 35404 77588 35460 77644
rect 31052 77532 31108 77588
rect 35756 77532 35812 77588
rect 27020 77420 27076 77476
rect 26012 77196 26068 77252
rect 27468 76972 27524 77028
rect 19836 76804 19892 76860
rect 19940 76804 19996 76860
rect 20044 76804 20100 76860
rect 26908 76636 26964 76692
rect 27580 76524 27636 76580
rect 26124 76300 26180 76356
rect 35756 76300 35812 76356
rect 4476 76020 4532 76076
rect 4580 76020 4636 76076
rect 4684 76020 4740 76076
rect 35196 76020 35252 76076
rect 35300 76020 35356 76076
rect 35404 76020 35460 76076
rect 27244 75516 27300 75572
rect 35756 75404 35812 75460
rect 19836 75236 19892 75292
rect 19940 75236 19996 75292
rect 20044 75236 20100 75292
rect 30492 75180 30548 75236
rect 31052 75180 31108 75236
rect 35756 74620 35812 74676
rect 4476 74452 4532 74508
rect 4580 74452 4636 74508
rect 4684 74452 4740 74508
rect 35196 74452 35252 74508
rect 35300 74452 35356 74508
rect 35404 74452 35460 74508
rect 34412 74172 34468 74228
rect 35644 74172 35700 74228
rect 35756 73836 35812 73892
rect 19836 73668 19892 73724
rect 19940 73668 19996 73724
rect 20044 73668 20100 73724
rect 34412 73500 34468 73556
rect 4476 72884 4532 72940
rect 4580 72884 4636 72940
rect 4684 72884 4740 72940
rect 35196 72884 35252 72940
rect 35300 72884 35356 72940
rect 35404 72884 35460 72940
rect 36092 72268 36148 72324
rect 19836 72100 19892 72156
rect 19940 72100 19996 72156
rect 20044 72100 20100 72156
rect 4476 71316 4532 71372
rect 4580 71316 4636 71372
rect 4684 71316 4740 71372
rect 35196 71316 35252 71372
rect 35300 71316 35356 71372
rect 35404 71316 35460 71372
rect 29596 71148 29652 71204
rect 34188 71036 34244 71092
rect 36092 70588 36148 70644
rect 19836 70532 19892 70588
rect 19940 70532 19996 70588
rect 20044 70532 20100 70588
rect 29148 70364 29204 70420
rect 4476 69748 4532 69804
rect 4580 69748 4636 69804
rect 4684 69748 4740 69804
rect 35196 69748 35252 69804
rect 35300 69748 35356 69804
rect 35404 69748 35460 69804
rect 19836 68964 19892 69020
rect 19940 68964 19996 69020
rect 20044 68964 20100 69020
rect 21084 68684 21140 68740
rect 29596 68236 29652 68292
rect 4476 68180 4532 68236
rect 4580 68180 4636 68236
rect 4684 68180 4740 68236
rect 35196 68180 35252 68236
rect 35300 68180 35356 68236
rect 35404 68180 35460 68236
rect 19836 67396 19892 67452
rect 19940 67396 19996 67452
rect 20044 67396 20100 67452
rect 4476 66612 4532 66668
rect 4580 66612 4636 66668
rect 4684 66612 4740 66668
rect 35196 66612 35252 66668
rect 35300 66612 35356 66668
rect 35404 66612 35460 66668
rect 19836 65828 19892 65884
rect 19940 65828 19996 65884
rect 20044 65828 20100 65884
rect 4476 65044 4532 65100
rect 4580 65044 4636 65100
rect 4684 65044 4740 65100
rect 35196 65044 35252 65100
rect 35300 65044 35356 65100
rect 35404 65044 35460 65100
rect 29484 64876 29540 64932
rect 19836 64260 19892 64316
rect 19940 64260 19996 64316
rect 20044 64260 20100 64316
rect 4476 63476 4532 63532
rect 4580 63476 4636 63532
rect 4684 63476 4740 63532
rect 35196 63476 35252 63532
rect 35300 63476 35356 63532
rect 35404 63476 35460 63532
rect 19836 62692 19892 62748
rect 19940 62692 19996 62748
rect 20044 62692 20100 62748
rect 25676 62524 25732 62580
rect 29484 62300 29540 62356
rect 4476 61908 4532 61964
rect 4580 61908 4636 61964
rect 4684 61908 4740 61964
rect 35196 61908 35252 61964
rect 35300 61908 35356 61964
rect 35404 61908 35460 61964
rect 21084 61628 21140 61684
rect 29148 61404 29204 61460
rect 19836 61124 19892 61180
rect 19940 61124 19996 61180
rect 20044 61124 20100 61180
rect 4476 60340 4532 60396
rect 4580 60340 4636 60396
rect 4684 60340 4740 60396
rect 35196 60340 35252 60396
rect 35300 60340 35356 60396
rect 35404 60340 35460 60396
rect 19836 59556 19892 59612
rect 19940 59556 19996 59612
rect 20044 59556 20100 59612
rect 25676 59164 25732 59220
rect 21084 59052 21140 59108
rect 4476 58772 4532 58828
rect 4580 58772 4636 58828
rect 4684 58772 4740 58828
rect 35196 58772 35252 58828
rect 35300 58772 35356 58828
rect 35404 58772 35460 58828
rect 19836 57988 19892 58044
rect 19940 57988 19996 58044
rect 20044 57988 20100 58044
rect 16828 57708 16884 57764
rect 19628 57372 19684 57428
rect 4476 57204 4532 57260
rect 4580 57204 4636 57260
rect 4684 57204 4740 57260
rect 35196 57204 35252 57260
rect 35300 57204 35356 57260
rect 35404 57204 35460 57260
rect 18844 57036 18900 57092
rect 19292 57036 19348 57092
rect 19836 56420 19892 56476
rect 19940 56420 19996 56476
rect 20044 56420 20100 56476
rect 3948 55916 4004 55972
rect 4476 55636 4532 55692
rect 4580 55636 4636 55692
rect 4684 55636 4740 55692
rect 35196 55636 35252 55692
rect 35300 55636 35356 55692
rect 35404 55636 35460 55692
rect 21420 55020 21476 55076
rect 19836 54852 19892 54908
rect 19940 54852 19996 54908
rect 20044 54852 20100 54908
rect 11452 54796 11508 54852
rect 28476 54460 28532 54516
rect 4476 54068 4532 54124
rect 4580 54068 4636 54124
rect 4684 54068 4740 54124
rect 35196 54068 35252 54124
rect 35300 54068 35356 54124
rect 35404 54068 35460 54124
rect 3948 54012 4004 54068
rect 21644 53900 21700 53956
rect 19836 53284 19892 53340
rect 19940 53284 19996 53340
rect 20044 53284 20100 53340
rect 4956 53228 5012 53284
rect 21420 53116 21476 53172
rect 31500 52780 31556 52836
rect 18844 52556 18900 52612
rect 4476 52500 4532 52556
rect 4580 52500 4636 52556
rect 4684 52500 4740 52556
rect 35196 52500 35252 52556
rect 35300 52500 35356 52556
rect 35404 52500 35460 52556
rect 23324 52444 23380 52500
rect 4956 51996 5012 52052
rect 16828 51996 16884 52052
rect 19292 51884 19348 51940
rect 19836 51716 19892 51772
rect 19940 51716 19996 51772
rect 20044 51716 20100 51772
rect 19628 51660 19684 51716
rect 28476 51100 28532 51156
rect 4476 50932 4532 50988
rect 4580 50932 4636 50988
rect 4684 50932 4740 50988
rect 35196 50932 35252 50988
rect 35300 50932 35356 50988
rect 35404 50932 35460 50988
rect 19836 50148 19892 50204
rect 19940 50148 19996 50204
rect 20044 50148 20100 50204
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 11452 48636 11508 48692
rect 23436 48636 23492 48692
rect 19836 48580 19892 48636
rect 19940 48580 19996 48636
rect 20044 48580 20100 48636
rect 23324 48412 23380 48468
rect 23436 48076 23492 48132
rect 21644 47852 21700 47908
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 31500 47180 31556 47236
rect 28588 46956 28644 47012
rect 27916 46844 27972 46900
rect 24332 46732 24388 46788
rect 26684 46732 26740 46788
rect 25564 46508 25620 46564
rect 28140 46508 28196 46564
rect 26908 46396 26964 46452
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 26236 46284 26292 46340
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 29148 46172 29204 46228
rect 25564 45948 25620 46004
rect 27916 45948 27972 46004
rect 22876 45836 22932 45892
rect 24444 45836 24500 45892
rect 28364 45836 28420 45892
rect 20748 45724 20804 45780
rect 28140 45724 28196 45780
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 23212 45388 23268 45444
rect 28252 45388 28308 45444
rect 5628 45276 5684 45332
rect 28476 45276 28532 45332
rect 28588 45164 28644 45220
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 21196 44604 21252 44660
rect 21532 44492 21588 44548
rect 30940 44380 30996 44436
rect 3612 44156 3668 44212
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 21532 43372 21588 43428
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 21196 43036 21252 43092
rect 20748 42812 20804 42868
rect 28364 42700 28420 42756
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 15932 42252 15988 42308
rect 26684 42140 26740 42196
rect 20748 42028 20804 42084
rect 21532 42028 21588 42084
rect 22428 41916 22484 41972
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 22540 41692 22596 41748
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 30940 41468 30996 41524
rect 22876 41132 22932 41188
rect 28140 41020 28196 41076
rect 15708 40908 15764 40964
rect 22204 40796 22260 40852
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 20300 40460 20356 40516
rect 22652 40460 22708 40516
rect 29148 40348 29204 40404
rect 6524 40236 6580 40292
rect 22540 40236 22596 40292
rect 26908 40124 26964 40180
rect 22316 40012 22372 40068
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 28252 39676 28308 39732
rect 5628 39564 5684 39620
rect 22204 39564 22260 39620
rect 22428 39340 22484 39396
rect 15932 39228 15988 39284
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 24444 39004 24500 39060
rect 26236 39004 26292 39060
rect 16492 38892 16548 38948
rect 16044 38780 16100 38836
rect 16380 38556 16436 38612
rect 22652 38556 22708 38612
rect 22316 38444 22372 38500
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 22428 38332 22484 38388
rect 24332 38220 24388 38276
rect 22204 37884 22260 37940
rect 15596 37772 15652 37828
rect 15932 37772 15988 37828
rect 16492 37772 16548 37828
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 16380 37436 16436 37492
rect 20300 37436 20356 37492
rect 28252 37324 28308 37380
rect 6524 36876 6580 36932
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19628 36428 19684 36484
rect 23212 36204 23268 36260
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 18620 35644 18676 35700
rect 3612 35308 3668 35364
rect 19628 35308 19684 35364
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 35644 35196 35700 35252
rect 17724 35084 17780 35140
rect 18956 34972 19012 35028
rect 35644 34748 35700 34804
rect 17388 34524 17444 34580
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 35644 34300 35700 34356
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 17388 33404 17444 33460
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 18956 30828 19012 30884
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 26796 29484 26852 29540
rect 17276 29372 17332 29428
rect 35644 29260 35700 29316
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 18620 28588 18676 28644
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 17724 26908 17780 26964
rect 17276 26684 17332 26740
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 26796 25116 26852 25172
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 19180 12348 19236 12404
rect 19068 12236 19124 12292
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19180 11676 19236 11732
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 17724 10780 17780 10836
rect 19068 10556 19124 10612
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 17724 9996 17780 10052
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
rect 4476 2324 4532 2380
rect 4580 2324 4636 2380
rect 4684 2324 4740 2380
rect 35196 2324 35252 2380
rect 35300 2324 35356 2380
rect 35404 2324 35460 2380
rect 19836 1540 19892 1596
rect 19940 1540 19996 1596
rect 20044 1540 20100 1596
<< metal4 >>
rect 4448 98028 4768 98060
rect 4448 97972 4476 98028
rect 4532 97972 4580 98028
rect 4636 97972 4684 98028
rect 4740 97972 4768 98028
rect 4448 96460 4768 97972
rect 4448 96404 4476 96460
rect 4532 96404 4580 96460
rect 4636 96404 4684 96460
rect 4740 96404 4768 96460
rect 4448 94892 4768 96404
rect 4448 94836 4476 94892
rect 4532 94836 4580 94892
rect 4636 94836 4684 94892
rect 4740 94836 4768 94892
rect 4448 93324 4768 94836
rect 4448 93268 4476 93324
rect 4532 93268 4580 93324
rect 4636 93268 4684 93324
rect 4740 93268 4768 93324
rect 4448 91756 4768 93268
rect 4448 91700 4476 91756
rect 4532 91700 4580 91756
rect 4636 91700 4684 91756
rect 4740 91700 4768 91756
rect 4448 90188 4768 91700
rect 4448 90132 4476 90188
rect 4532 90132 4580 90188
rect 4636 90132 4684 90188
rect 4740 90132 4768 90188
rect 4448 88620 4768 90132
rect 4448 88564 4476 88620
rect 4532 88564 4580 88620
rect 4636 88564 4684 88620
rect 4740 88564 4768 88620
rect 4448 87052 4768 88564
rect 4448 86996 4476 87052
rect 4532 86996 4580 87052
rect 4636 86996 4684 87052
rect 4740 86996 4768 87052
rect 4448 85484 4768 86996
rect 4448 85428 4476 85484
rect 4532 85428 4580 85484
rect 4636 85428 4684 85484
rect 4740 85428 4768 85484
rect 4448 83916 4768 85428
rect 4448 83860 4476 83916
rect 4532 83860 4580 83916
rect 4636 83860 4684 83916
rect 4740 83860 4768 83916
rect 4448 82348 4768 83860
rect 4448 82292 4476 82348
rect 4532 82292 4580 82348
rect 4636 82292 4684 82348
rect 4740 82292 4768 82348
rect 4448 80780 4768 82292
rect 4448 80724 4476 80780
rect 4532 80724 4580 80780
rect 4636 80724 4684 80780
rect 4740 80724 4768 80780
rect 4448 79212 4768 80724
rect 4448 79156 4476 79212
rect 4532 79156 4580 79212
rect 4636 79156 4684 79212
rect 4740 79156 4768 79212
rect 4448 77644 4768 79156
rect 4448 77588 4476 77644
rect 4532 77588 4580 77644
rect 4636 77588 4684 77644
rect 4740 77588 4768 77644
rect 4448 76076 4768 77588
rect 4448 76020 4476 76076
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4740 76020 4768 76076
rect 4448 74508 4768 76020
rect 4448 74452 4476 74508
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4740 74452 4768 74508
rect 4448 72940 4768 74452
rect 4448 72884 4476 72940
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4740 72884 4768 72940
rect 4448 71372 4768 72884
rect 4448 71316 4476 71372
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4740 71316 4768 71372
rect 4448 69804 4768 71316
rect 4448 69748 4476 69804
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4740 69748 4768 69804
rect 4448 68236 4768 69748
rect 4448 68180 4476 68236
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4740 68180 4768 68236
rect 4448 66668 4768 68180
rect 4448 66612 4476 66668
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4740 66612 4768 66668
rect 4448 65100 4768 66612
rect 4448 65044 4476 65100
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4740 65044 4768 65100
rect 4448 63532 4768 65044
rect 4448 63476 4476 63532
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4740 63476 4768 63532
rect 4448 61964 4768 63476
rect 4448 61908 4476 61964
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4740 61908 4768 61964
rect 4448 60396 4768 61908
rect 4448 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4768 60396
rect 4448 58828 4768 60340
rect 4448 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4768 58828
rect 4448 57260 4768 58772
rect 19808 97244 20128 98060
rect 19808 97188 19836 97244
rect 19892 97188 19940 97244
rect 19996 97188 20044 97244
rect 20100 97188 20128 97244
rect 19808 95676 20128 97188
rect 19808 95620 19836 95676
rect 19892 95620 19940 95676
rect 19996 95620 20044 95676
rect 20100 95620 20128 95676
rect 19808 94108 20128 95620
rect 35168 98028 35488 98060
rect 35168 97972 35196 98028
rect 35252 97972 35300 98028
rect 35356 97972 35404 98028
rect 35460 97972 35488 98028
rect 35168 96460 35488 97972
rect 35168 96404 35196 96460
rect 35252 96404 35300 96460
rect 35356 96404 35404 96460
rect 35460 96404 35488 96460
rect 19808 94052 19836 94108
rect 19892 94052 19940 94108
rect 19996 94052 20044 94108
rect 20100 94052 20128 94108
rect 19808 92540 20128 94052
rect 25116 95508 25172 95518
rect 19808 92484 19836 92540
rect 19892 92484 19940 92540
rect 19996 92484 20044 92540
rect 20100 92484 20128 92540
rect 19808 90972 20128 92484
rect 19808 90916 19836 90972
rect 19892 90916 19940 90972
rect 19996 90916 20044 90972
rect 20100 90916 20128 90972
rect 19808 89404 20128 90916
rect 19808 89348 19836 89404
rect 19892 89348 19940 89404
rect 19996 89348 20044 89404
rect 20100 89348 20128 89404
rect 19808 87836 20128 89348
rect 19808 87780 19836 87836
rect 19892 87780 19940 87836
rect 19996 87780 20044 87836
rect 20100 87780 20128 87836
rect 19808 86268 20128 87780
rect 24444 93492 24500 93502
rect 24444 86884 24500 93436
rect 24556 90692 24612 90702
rect 24556 89796 24612 90636
rect 24556 87556 24612 89740
rect 24556 87490 24612 87500
rect 24444 86818 24500 86828
rect 19808 86212 19836 86268
rect 19892 86212 19940 86268
rect 19996 86212 20044 86268
rect 20100 86212 20128 86268
rect 19808 84700 20128 86212
rect 19808 84644 19836 84700
rect 19892 84644 19940 84700
rect 19996 84644 20044 84700
rect 20100 84644 20128 84700
rect 19808 83132 20128 84644
rect 25116 84196 25172 95452
rect 35168 94892 35488 96404
rect 35168 94836 35196 94892
rect 35252 94836 35300 94892
rect 35356 94836 35404 94892
rect 35460 94836 35488 94892
rect 35168 93324 35488 94836
rect 35168 93268 35196 93324
rect 35252 93268 35300 93324
rect 35356 93268 35404 93324
rect 35460 93268 35488 93324
rect 35168 91756 35488 93268
rect 35168 91700 35196 91756
rect 35252 91700 35300 91756
rect 35356 91700 35404 91756
rect 35460 91700 35488 91756
rect 35168 90188 35488 91700
rect 35168 90132 35196 90188
rect 35252 90132 35300 90188
rect 35356 90132 35404 90188
rect 35460 90132 35488 90188
rect 27468 89572 27524 89582
rect 25116 84130 25172 84140
rect 26012 86660 26068 86670
rect 26012 83300 26068 86604
rect 26012 83234 26068 83244
rect 27356 84196 27412 84206
rect 19808 83076 19836 83132
rect 19892 83076 19940 83132
rect 19996 83076 20044 83132
rect 20100 83076 20128 83132
rect 19808 81564 20128 83076
rect 19808 81508 19836 81564
rect 19892 81508 19940 81564
rect 19996 81508 20044 81564
rect 20100 81508 20128 81564
rect 19808 79996 20128 81508
rect 19808 79940 19836 79996
rect 19892 79940 19940 79996
rect 19996 79940 20044 79996
rect 20100 79940 20128 79996
rect 19808 78428 20128 79940
rect 27244 82404 27300 82414
rect 27020 79156 27076 79166
rect 26908 78932 26964 78942
rect 19808 78372 19836 78428
rect 19892 78372 19940 78428
rect 19996 78372 20044 78428
rect 20100 78372 20128 78428
rect 19808 76860 20128 78372
rect 26012 78708 26068 78718
rect 25788 78148 25844 78158
rect 25788 77924 25844 78092
rect 25788 77858 25844 77868
rect 26012 77252 26068 78652
rect 26012 77186 26068 77196
rect 26124 78148 26180 78158
rect 19808 76804 19836 76860
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 20100 76804 20128 76860
rect 19808 75292 20128 76804
rect 26124 76356 26180 78092
rect 26908 76692 26964 78876
rect 27020 77476 27076 79100
rect 27020 77410 27076 77420
rect 26908 76626 26964 76636
rect 26124 76290 26180 76300
rect 27244 75572 27300 82348
rect 27356 81396 27412 84140
rect 27356 81330 27412 81340
rect 27468 77028 27524 89516
rect 35168 88620 35488 90132
rect 35168 88564 35196 88620
rect 35252 88564 35300 88620
rect 35356 88564 35404 88620
rect 35460 88564 35488 88620
rect 35168 87052 35488 88564
rect 35168 86996 35196 87052
rect 35252 86996 35300 87052
rect 35356 86996 35404 87052
rect 35460 86996 35488 87052
rect 35168 85484 35488 86996
rect 35168 85428 35196 85484
rect 35252 85428 35300 85484
rect 35356 85428 35404 85484
rect 35460 85428 35488 85484
rect 35168 83916 35488 85428
rect 35168 83860 35196 83916
rect 35252 83860 35300 83916
rect 35356 83860 35404 83916
rect 35460 83860 35488 83916
rect 35168 82348 35488 83860
rect 35168 82292 35196 82348
rect 35252 82292 35300 82348
rect 35356 82292 35404 82348
rect 35460 82292 35488 82348
rect 35168 80780 35488 82292
rect 34188 80724 34244 80734
rect 30492 79268 30548 79278
rect 27468 76962 27524 76972
rect 27580 79044 27636 79054
rect 27580 76580 27636 78988
rect 27580 76514 27636 76524
rect 27244 75506 27300 75516
rect 19808 75236 19836 75292
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 20100 75236 20128 75292
rect 19808 73724 20128 75236
rect 30492 75236 30548 79212
rect 30492 75170 30548 75180
rect 31052 77588 31108 77598
rect 31052 75236 31108 77532
rect 31052 75170 31108 75180
rect 19808 73668 19836 73724
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 20100 73668 20128 73724
rect 19808 72156 20128 73668
rect 19808 72100 19836 72156
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 20100 72100 20128 72156
rect 19808 70588 20128 72100
rect 19808 70532 19836 70588
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 20100 70532 20128 70588
rect 19808 69020 20128 70532
rect 29596 71204 29652 71214
rect 19808 68964 19836 69020
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 20100 68964 20128 69020
rect 19808 67452 20128 68964
rect 29148 70420 29204 70430
rect 19808 67396 19836 67452
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 20100 67396 20128 67452
rect 19808 65884 20128 67396
rect 19808 65828 19836 65884
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 20100 65828 20128 65884
rect 19808 64316 20128 65828
rect 19808 64260 19836 64316
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 20100 64260 20128 64316
rect 19808 62748 20128 64260
rect 19808 62692 19836 62748
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 20100 62692 20128 62748
rect 19808 61180 20128 62692
rect 19808 61124 19836 61180
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 20100 61124 20128 61180
rect 19808 59612 20128 61124
rect 19808 59556 19836 59612
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 20100 59556 20128 59612
rect 19808 58044 20128 59556
rect 21084 68740 21140 68750
rect 21084 61684 21140 68684
rect 21084 59108 21140 61628
rect 25676 62580 25732 62590
rect 25676 59220 25732 62524
rect 29148 61460 29204 70364
rect 29596 68292 29652 71148
rect 34188 71092 34244 80668
rect 35168 80724 35196 80780
rect 35252 80724 35300 80780
rect 35356 80724 35404 80780
rect 35460 80724 35488 80780
rect 35168 79212 35488 80724
rect 35168 79156 35196 79212
rect 35252 79156 35300 79212
rect 35356 79156 35404 79212
rect 35460 79156 35488 79212
rect 35168 77644 35488 79156
rect 35168 77588 35196 77644
rect 35252 77588 35300 77644
rect 35356 77588 35404 77644
rect 35460 77588 35488 77644
rect 35168 76076 35488 77588
rect 35168 76020 35196 76076
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35460 76020 35488 76076
rect 35168 74508 35488 76020
rect 35168 74452 35196 74508
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35460 74452 35488 74508
rect 34412 74228 34468 74238
rect 34412 73556 34468 74172
rect 34412 73490 34468 73500
rect 34188 71026 34244 71036
rect 35168 72940 35488 74452
rect 35644 81732 35700 81742
rect 35644 74228 35700 81676
rect 35756 77588 35812 77598
rect 35756 76356 35812 77532
rect 35756 75460 35812 76300
rect 35756 75394 35812 75404
rect 35644 74162 35700 74172
rect 35756 74676 35812 74686
rect 35756 73892 35812 74620
rect 35756 73826 35812 73836
rect 35168 72884 35196 72940
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35460 72884 35488 72940
rect 35168 71372 35488 72884
rect 35168 71316 35196 71372
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35460 71316 35488 71372
rect 29596 68226 29652 68236
rect 35168 69804 35488 71316
rect 36092 72324 36148 72334
rect 36092 70644 36148 72268
rect 36092 70578 36148 70588
rect 35168 69748 35196 69804
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35460 69748 35488 69804
rect 35168 68236 35488 69748
rect 35168 68180 35196 68236
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35460 68180 35488 68236
rect 35168 66668 35488 68180
rect 35168 66612 35196 66668
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35460 66612 35488 66668
rect 35168 65100 35488 66612
rect 35168 65044 35196 65100
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35460 65044 35488 65100
rect 29484 64932 29540 64942
rect 29484 62356 29540 64876
rect 29484 62290 29540 62300
rect 35168 63532 35488 65044
rect 35168 63476 35196 63532
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35460 63476 35488 63532
rect 29148 61394 29204 61404
rect 35168 61964 35488 63476
rect 35168 61908 35196 61964
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35460 61908 35488 61964
rect 25676 59154 25732 59164
rect 35168 60396 35488 61908
rect 35168 60340 35196 60396
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35460 60340 35488 60396
rect 21084 59042 21140 59052
rect 19808 57988 19836 58044
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20100 57988 20128 58044
rect 4448 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4768 57260
rect 3948 55972 4004 55982
rect 3948 54068 4004 55916
rect 3948 54002 4004 54012
rect 4448 55692 4768 57204
rect 4448 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4768 55692
rect 4448 54124 4768 55636
rect 16828 57764 16884 57774
rect 4448 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4768 54124
rect 4448 52556 4768 54068
rect 11452 54852 11508 54862
rect 4448 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4768 52556
rect 4448 50988 4768 52500
rect 4956 53284 5012 53294
rect 4956 52052 5012 53228
rect 4956 51986 5012 51996
rect 4448 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4768 50988
rect 4448 49420 4768 50932
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 4448 47852 4768 49364
rect 11452 48692 11508 54796
rect 16828 52052 16884 57708
rect 19628 57428 19684 57438
rect 18844 57092 18900 57102
rect 18844 52612 18900 57036
rect 18844 52546 18900 52556
rect 19292 57092 19348 57102
rect 16828 51986 16884 51996
rect 19292 51940 19348 57036
rect 19292 51874 19348 51884
rect 19628 51716 19684 57372
rect 19628 51650 19684 51660
rect 19808 56476 20128 57988
rect 19808 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20128 56476
rect 19808 54908 20128 56420
rect 35168 58828 35488 60340
rect 35168 58772 35196 58828
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35460 58772 35488 58828
rect 35168 57260 35488 58772
rect 35168 57204 35196 57260
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35460 57204 35488 57260
rect 35168 55692 35488 57204
rect 35168 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35488 55692
rect 19808 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20128 54908
rect 19808 53340 20128 54852
rect 19808 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20128 53340
rect 19808 51772 20128 53284
rect 21420 55076 21476 55086
rect 21420 53172 21476 55020
rect 28476 54516 28532 54526
rect 21420 53106 21476 53116
rect 21644 53956 21700 53966
rect 19808 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20128 51772
rect 11452 48626 11508 48636
rect 19808 50204 20128 51716
rect 19808 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20128 50204
rect 19808 48636 20128 50148
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4448 46284 4768 47796
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 19808 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20128 48636
rect 19808 47068 20128 48580
rect 21644 47908 21700 53900
rect 23324 52500 23380 52510
rect 23324 48468 23380 52444
rect 28476 51156 28532 54460
rect 35168 54124 35488 55636
rect 35168 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35488 54124
rect 23324 48402 23380 48412
rect 23436 48692 23492 48702
rect 23436 48132 23492 48636
rect 23436 48066 23492 48076
rect 21644 47842 21700 47852
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 19808 45500 20128 47012
rect 27916 46900 27972 46910
rect 24332 46788 24388 46798
rect 22876 45892 22932 45902
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 3612 44212 3668 44222
rect 3612 35364 3668 44156
rect 3612 35298 3668 35308
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 5628 45332 5684 45342
rect 5628 39620 5684 45276
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 15932 42308 15988 42318
rect 15708 40964 15764 40974
rect 5628 39554 5684 39564
rect 6524 40292 6580 40302
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 6524 36932 6580 40236
rect 15708 38668 15764 40908
rect 15932 39284 15988 42252
rect 15932 39218 15988 39228
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 20748 45780 20804 45790
rect 20748 42868 20804 45724
rect 21196 44660 21252 44670
rect 21196 43092 21252 44604
rect 21196 43026 21252 43036
rect 21532 44548 21588 44558
rect 21532 43428 21588 44492
rect 20748 42084 20804 42812
rect 20748 42018 20804 42028
rect 21532 42084 21588 43372
rect 21532 42018 21588 42028
rect 22428 41972 22484 41982
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 22204 40852 22260 40862
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 16492 38948 16548 38958
rect 16044 38836 16100 38846
rect 16044 38668 16100 38780
rect 15596 38612 15764 38668
rect 15932 38612 16100 38668
rect 16380 38612 16436 38622
rect 15596 37828 15652 38612
rect 15596 37762 15652 37772
rect 15932 37828 15988 38612
rect 15932 37762 15988 37772
rect 16380 37492 16436 38556
rect 16492 37828 16548 38892
rect 16492 37762 16548 37772
rect 16380 37426 16436 37436
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 6524 36866 6580 36876
rect 4448 35308 4768 36820
rect 19628 36484 19684 36494
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 18620 35700 18676 35710
rect 17724 35140 17780 35150
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 17388 34580 17444 34590
rect 17388 33460 17444 34524
rect 17388 33394 17444 33404
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 17276 29428 17332 29438
rect 17276 26740 17332 29372
rect 17724 26964 17780 35084
rect 18620 28644 18676 35644
rect 19628 35364 19684 36428
rect 19628 35298 19684 35308
rect 19808 36092 20128 37604
rect 20300 40516 20356 40526
rect 20300 37492 20356 40460
rect 22204 39620 22260 40796
rect 22204 37940 22260 39564
rect 22316 40068 22372 40078
rect 22316 38500 22372 40012
rect 22316 38434 22372 38444
rect 22428 39396 22484 41916
rect 22540 41748 22596 41758
rect 22540 40292 22596 41692
rect 22876 41188 22932 45836
rect 22876 41122 22932 41132
rect 23212 45444 23268 45454
rect 22540 40226 22596 40236
rect 22652 40516 22708 40526
rect 22428 38388 22484 39340
rect 22652 38612 22708 40460
rect 22652 38546 22708 38556
rect 22428 38322 22484 38332
rect 22204 37874 22260 37884
rect 20300 37426 20356 37436
rect 23212 36260 23268 45388
rect 24332 38276 24388 46732
rect 26684 46788 26740 46798
rect 25564 46564 25620 46574
rect 25564 46004 25620 46508
rect 25564 45938 25620 45948
rect 26236 46340 26292 46350
rect 24444 45892 24500 45902
rect 24444 39060 24500 45836
rect 24444 38994 24500 39004
rect 26236 39060 26292 46284
rect 26684 42196 26740 46732
rect 26684 42130 26740 42140
rect 26908 46452 26964 46462
rect 26908 40180 26964 46396
rect 27916 46004 27972 46844
rect 27916 45938 27972 45948
rect 28140 46564 28196 46574
rect 28140 45780 28196 46508
rect 28140 41076 28196 45724
rect 28364 45892 28420 45902
rect 28140 41010 28196 41020
rect 28252 45444 28308 45454
rect 26908 40114 26964 40124
rect 26236 38994 26292 39004
rect 28252 39732 28308 45388
rect 28364 42756 28420 45836
rect 28476 45332 28532 51100
rect 31500 52836 31556 52846
rect 31500 47236 31556 52780
rect 31500 47170 31556 47180
rect 35168 52556 35488 54068
rect 35168 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35488 52556
rect 35168 50988 35488 52500
rect 35168 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35488 50988
rect 35168 49420 35488 50932
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 35168 47852 35488 49364
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 28476 45266 28532 45276
rect 28588 47012 28644 47022
rect 28588 45220 28644 46956
rect 35168 46284 35488 47796
rect 28588 45154 28644 45164
rect 29148 46228 29204 46238
rect 28364 42690 28420 42700
rect 29148 40404 29204 46172
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 30940 44436 30996 44446
rect 30940 41524 30996 44380
rect 30940 41458 30996 41468
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 29148 40338 29204 40348
rect 24332 38210 24388 38220
rect 28252 37380 28308 39676
rect 28252 37314 28308 37324
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 23212 36194 23268 36204
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 18956 35028 19012 35038
rect 18956 30884 19012 34972
rect 18956 30818 19012 30828
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 18620 28578 18676 28588
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 17724 26898 17780 26908
rect 19808 28252 20128 29764
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35644 35252 35700 35262
rect 35644 34804 35700 35196
rect 35644 34738 35700 34748
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 17276 26674 17332 26684
rect 19808 26684 20128 28196
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 26796 29540 26852 29550
rect 26796 25172 26852 29484
rect 26796 25106 26852 25116
rect 35168 29036 35488 30548
rect 35644 34356 35700 34366
rect 35644 29316 35700 34300
rect 35644 29250 35700 29260
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19180 12404 19236 12414
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 19068 12292 19124 12302
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 17724 10836 17780 10846
rect 17724 10052 17780 10780
rect 19068 10612 19124 12236
rect 19180 11732 19236 12348
rect 19180 11666 19236 11676
rect 19068 10546 19124 10556
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 17724 9986 17780 9996
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 2380 4768 3892
rect 4448 2324 4476 2380
rect 4532 2324 4580 2380
rect 4636 2324 4684 2380
rect 4740 2324 4768 2380
rect 4448 1508 4768 2324
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 1596 20128 3108
rect 19808 1540 19836 1596
rect 19892 1540 19940 1596
rect 19996 1540 20044 1596
rect 20100 1540 20128 1596
rect 19808 1508 20128 1540
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 2380 35488 3892
rect 35168 2324 35196 2380
rect 35252 2324 35300 2380
rect 35356 2324 35404 2380
rect 35460 2324 35488 2380
rect 35168 1508 35488 2324
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _0842_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 35056 0 1 81536
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0843_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29008 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0844_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 16016 0 -1 87808
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0845_
timestamp 1698431365
transform 1 0 20608 0 -1 89376
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0846_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21280 0 1 79968
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_4  _0847_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19824 0 1 83104
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _0848_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 19824 0 1 79968
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0849_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13888 0 1 83104
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0850_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14448 0 1 84672
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0851_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 19152 0 -1 87808
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0852_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29008 0 1 84672
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0853_
timestamp 1698431365
transform 1 0 30688 0 -1 87808
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0854_
timestamp 1698431365
transform 1 0 32928 0 -1 86240
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _0855_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 34160 0 1 84672
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _0856_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 35168 0 -1 84672
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _0857_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18704 0 -1 79968
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  _0858_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21168 0 1 75264
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0859_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 30912 0 1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0860_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 30240 0 1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_12  _0861_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 16128 0 1 75264
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_8  _0862_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22848 0 -1 62720
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  _0863_
timestamp 1698431365
transform 1 0 29792 0 1 64288
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0864_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 37184 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_12  _0865_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21952 0 1 68992
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _0866_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21168 0 1 62720
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _0867_
timestamp 1698431365
transform 1 0 18704 0 -1 72128
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_12  _0868_
timestamp 1698431365
transform 1 0 14112 0 1 73696
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _0869_
timestamp 1698431365
transform 1 0 21168 0 1 45472
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__and2_4  _0870_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 19824 0 -1 47040
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  _0871_
timestamp 1698431365
transform 1 0 21616 0 1 61152
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0872_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 26544 0 1 42336
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  _0873_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 23184 0 -1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _0874_
timestamp 1698431365
transform 1 0 14672 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _0875_
timestamp 1698431365
transform 1 0 20160 0 -1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0876_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19264 0 -1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _0877_
timestamp 1698431365
transform -1 0 23184 0 1 50176
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0878_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 30128 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0879_
timestamp 1698431365
transform 1 0 29344 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _0880_
timestamp 1698431365
transform 1 0 22960 0 1 54880
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _0881_
timestamp 1698431365
transform -1 0 23520 0 -1 64288
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__and3_2  _0882_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26992 0 1 43904
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0883_
timestamp 1698431365
transform 1 0 30464 0 -1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _0884_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17360 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0885_
timestamp 1698431365
transform 1 0 17248 0 -1 48608
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0886_
timestamp 1698431365
transform 1 0 18144 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  _0887_
timestamp 1698431365
transform 1 0 17920 0 -1 51744
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0888_
timestamp 1698431365
transform 1 0 29904 0 1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__inv_4  _0889_
timestamp 1698431365
transform 1 0 21840 0 1 59584
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0890_
timestamp 1698431365
transform -1 0 26992 0 1 43904
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0891_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26656 0 -1 29792
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  _0892_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 24080 0 1 70560
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0893_
timestamp 1698431365
transform 1 0 26208 0 -1 28224
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0894_
timestamp 1698431365
transform 1 0 27440 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0895_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 30800 0 -1 34496
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _0896_
timestamp 1698431365
transform 1 0 17920 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _0897_
timestamp 1698431365
transform 1 0 17248 0 -1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__or2_4  _0898_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15008 0 -1 45472
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0899_
timestamp 1698431365
transform 1 0 16800 0 1 40768
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0900_
timestamp 1698431365
transform 1 0 15232 0 1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _0901_
timestamp 1698431365
transform -1 0 16800 0 1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0902_
timestamp 1698431365
transform 1 0 16352 0 1 42336
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0903_
timestamp 1698431365
transform 1 0 5264 0 -1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0904_
timestamp 1698431365
transform 1 0 16800 0 1 50176
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _0905_
timestamp 1698431365
transform 1 0 17248 0 -1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0906_
timestamp 1698431365
transform 1 0 4816 0 -1 53312
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0907_
timestamp 1698431365
transform 1 0 15792 0 1 43904
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0908_
timestamp 1698431365
transform -1 0 22512 0 -1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _0909_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 17024 0 -1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0910_
timestamp 1698431365
transform -1 0 7056 0 1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0911_
timestamp 1698431365
transform -1 0 20944 0 1 48608
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__and3_2  _0912_
timestamp 1698431365
transform 1 0 21504 0 -1 42336
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0913_
timestamp 1698431365
transform 1 0 5488 0 1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0914_
timestamp 1698431365
transform 1 0 5712 0 -1 39200
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0915_
timestamp 1698431365
transform -1 0 20608 0 1 53312
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0916_
timestamp 1698431365
transform 1 0 13328 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0917_
timestamp 1698431365
transform -1 0 24752 0 -1 64288
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0918_
timestamp 1698431365
transform -1 0 26656 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0919_
timestamp 1698431365
transform 1 0 18480 0 -1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0920_
timestamp 1698431365
transform 1 0 14336 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _0921_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 18368 0 1 65856
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0922_
timestamp 1698431365
transform 1 0 13776 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0923_
timestamp 1698431365
transform 1 0 21168 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _0924_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 16464 0 1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0925_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14896 0 -1 64288
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0926_
timestamp 1698431365
transform 1 0 17248 0 -1 64288
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0927_
timestamp 1698431365
transform 1 0 17696 0 -1 43904
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0928_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19152 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_2  _0929_
timestamp 1698431365
transform 1 0 21168 0 1 42336
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _0930_
timestamp 1698431365
transform 1 0 23072 0 -1 45472
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0931_
timestamp 1698431365
transform -1 0 24640 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and3_2  _0932_
timestamp 1698431365
transform -1 0 16576 0 1 45472
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0933_
timestamp 1698431365
transform 1 0 16576 0 1 45472
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0934_
timestamp 1698431365
transform 1 0 11648 0 1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0935_
timestamp 1698431365
transform 1 0 17360 0 -1 42336
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _0936_
timestamp 1698431365
transform 1 0 16576 0 1 39200
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0937_
timestamp 1698431365
transform 1 0 15904 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0938_
timestamp 1698431365
transform -1 0 18480 0 -1 15680
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0939_
timestamp 1698431365
transform 1 0 16240 0 1 37632
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0940_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29008 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0941_
timestamp 1698431365
transform 1 0 29120 0 1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _0942_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 28672 0 -1 65856
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0943_
timestamp 1698431365
transform 1 0 29008 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0944_
timestamp 1698431365
transform 1 0 33264 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0945_
timestamp 1698431365
transform -1 0 34496 0 -1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0946_
timestamp 1698431365
transform 1 0 33488 0 -1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0947_
timestamp 1698431365
transform 1 0 30688 0 1 29792
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0948_
timestamp 1698431365
transform 1 0 30800 0 1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0949_
timestamp 1698431365
transform 1 0 31696 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0950_
timestamp 1698431365
transform -1 0 34272 0 1 32928
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0951_
timestamp 1698431365
transform 1 0 15344 0 -1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0952_
timestamp 1698431365
transform 1 0 5488 0 1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0953_
timestamp 1698431365
transform 1 0 4256 0 1 58016
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0954_
timestamp 1698431365
transform 1 0 5040 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0955_
timestamp 1698431365
transform 1 0 4256 0 1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0956_
timestamp 1698431365
transform 1 0 5264 0 -1 37632
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0957_
timestamp 1698431365
transform 1 0 9856 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0958_
timestamp 1698431365
transform -1 0 24416 0 -1 65856
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0959_
timestamp 1698431365
transform -1 0 18368 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0960_
timestamp 1698431365
transform 1 0 18144 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _0961_
timestamp 1698431365
transform 1 0 17248 0 -1 67424
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0962_
timestamp 1698431365
transform -1 0 14448 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _0963_
timestamp 1698431365
transform -1 0 16464 0 1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0964_
timestamp 1698431365
transform 1 0 14784 0 -1 65856
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0965_
timestamp 1698431365
transform 1 0 17248 0 -1 65856
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0966_
timestamp 1698431365
transform 1 0 20384 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0967_
timestamp 1698431365
transform -1 0 26096 0 -1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0968_
timestamp 1698431365
transform 1 0 10080 0 -1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0969_
timestamp 1698431365
transform 1 0 15792 0 -1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0970_
timestamp 1698431365
transform -1 0 18480 0 -1 12544
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0971_
timestamp 1698431365
transform 1 0 17248 0 -1 36064
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0972_
timestamp 1698431365
transform 1 0 27216 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0973_
timestamp 1698431365
transform 1 0 29120 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _0974_
timestamp 1698431365
transform -1 0 32032 0 -1 61152
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0975_
timestamp 1698431365
transform -1 0 28784 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0976_
timestamp 1698431365
transform 1 0 34160 0 -1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0977_
timestamp 1698431365
transform -1 0 36288 0 1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0978_
timestamp 1698431365
transform -1 0 35952 0 1 47040
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0979_
timestamp 1698431365
transform 1 0 32368 0 1 29792
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0980_
timestamp 1698431365
transform 1 0 31920 0 -1 28224
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0981_
timestamp 1698431365
transform 1 0 32928 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0982_
timestamp 1698431365
transform -1 0 35728 0 -1 34496
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0983_
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0984_
timestamp 1698431365
transform 1 0 5600 0 1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _0985_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 7280 0 -1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0986_
timestamp 1698431365
transform 1 0 5600 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0987_
timestamp 1698431365
transform 1 0 5488 0 -1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0988_
timestamp 1698431365
transform 1 0 5824 0 -1 34496
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0989_
timestamp 1698431365
transform 1 0 10752 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0990_
timestamp 1698431365
transform -1 0 25312 0 1 64288
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0991_
timestamp 1698431365
transform -1 0 19936 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0992_
timestamp 1698431365
transform -1 0 21392 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _0993_
timestamp 1698431365
transform 1 0 18368 0 1 65856
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0994_
timestamp 1698431365
transform 1 0 14448 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _0995_
timestamp 1698431365
transform -1 0 17472 0 1 62720
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0996_
timestamp 1698431365
transform -1 0 16576 0 -1 62720
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0997_
timestamp 1698431365
transform 1 0 16800 0 1 64288
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0998_
timestamp 1698431365
transform 1 0 19488 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0999_
timestamp 1698431365
transform -1 0 27216 0 1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1000_
timestamp 1698431365
transform 1 0 10304 0 1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1001_
timestamp 1698431365
transform 1 0 17024 0 1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1002_
timestamp 1698431365
transform -1 0 19040 0 -1 10976
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1003_
timestamp 1698431365
transform 1 0 17696 0 1 34496
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1004_
timestamp 1698431365
transform 1 0 26880 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1005_
timestamp 1698431365
transform 1 0 28672 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1006_
timestamp 1698431365
transform -1 0 32480 0 1 59584
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1007_
timestamp 1698431365
transform -1 0 30128 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1008_
timestamp 1698431365
transform 1 0 34384 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1009_
timestamp 1698431365
transform -1 0 36512 0 1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1010_
timestamp 1698431365
transform -1 0 35952 0 1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1011_
timestamp 1698431365
transform 1 0 31808 0 -1 39200
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1012_
timestamp 1698431365
transform 1 0 32032 0 1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1013_
timestamp 1698431365
transform 1 0 32928 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1014_
timestamp 1698431365
transform -1 0 35504 0 1 39200
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1015_
timestamp 1698431365
transform 1 0 19152 0 -1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1016_
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1017_
timestamp 1698431365
transform 1 0 6608 0 1 58016
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1018_
timestamp 1698431365
transform -1 0 9184 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1019_
timestamp 1698431365
transform 1 0 9632 0 1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1020_
timestamp 1698431365
transform 1 0 8736 0 1 36064
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1021_
timestamp 1698431365
transform 1 0 8960 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1022_
timestamp 1698431365
transform -1 0 24416 0 1 59584
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1023_
timestamp 1698431365
transform -1 0 20384 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1024_
timestamp 1698431365
transform -1 0 22064 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _1025_
timestamp 1698431365
transform 1 0 18368 0 1 59584
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1026_
timestamp 1698431365
transform -1 0 16352 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1027_
timestamp 1698431365
transform 1 0 17248 0 -1 58016
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1028_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1029_
timestamp 1698431365
transform 1 0 18816 0 -1 59584
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1030_
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1031_
timestamp 1698431365
transform -1 0 27328 0 -1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1032_
timestamp 1698431365
transform 1 0 11872 0 -1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1033_
timestamp 1698431365
transform 1 0 18480 0 -1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1034_
timestamp 1698431365
transform -1 0 20384 0 1 10976
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1035_
timestamp 1698431365
transform 1 0 19376 0 -1 36064
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1036_
timestamp 1698431365
transform -1 0 30800 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1037_
timestamp 1698431365
transform 1 0 29792 0 1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1038_
timestamp 1698431365
transform -1 0 33152 0 1 58016
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1039_
timestamp 1698431365
transform -1 0 30352 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1040_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19376 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1041_
timestamp 1698431365
transform 1 0 12544 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1042_
timestamp 1698431365
transform 1 0 28784 0 -1 42336
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1043_
timestamp 1698431365
transform 1 0 20608 0 -1 50176
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1044_
timestamp 1698431365
transform -1 0 23072 0 -1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1045_
timestamp 1698431365
transform -1 0 25536 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1046_
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1047_
timestamp 1698431365
transform -1 0 26880 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1048_
timestamp 1698431365
transform -1 0 25872 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1049_
timestamp 1698431365
transform -1 0 34832 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1050_
timestamp 1698431365
transform 1 0 26544 0 -1 45472
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1051_
timestamp 1698431365
transform 1 0 26096 0 -1 42336
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1052_
timestamp 1698431365
transform -1 0 20944 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1053_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 28560 0 1 42336
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1054_
timestamp 1698431365
transform -1 0 25872 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1055_
timestamp 1698431365
transform 1 0 25088 0 -1 45472
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1056_
timestamp 1698431365
transform 1 0 25312 0 -1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1057_
timestamp 1698431365
transform 1 0 13664 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1058_
timestamp 1698431365
transform 1 0 25088 0 -1 39200
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1059_
timestamp 1698431365
transform -1 0 28784 0 1 39200
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1060_
timestamp 1698431365
transform -1 0 14896 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1061_
timestamp 1698431365
transform 1 0 14000 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1062_
timestamp 1698431365
transform 1 0 14896 0 1 47040
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1063_
timestamp 1698431365
transform -1 0 16688 0 -1 50176
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1064_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22512 0 -1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1065_
timestamp 1698431365
transform -1 0 20944 0 1 51744
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1066_
timestamp 1698431365
transform 1 0 19712 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1067_
timestamp 1698431365
transform -1 0 21728 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1068_
timestamp 1698431365
transform 1 0 18928 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1069_
timestamp 1698431365
transform -1 0 22624 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1070_
timestamp 1698431365
transform -1 0 24416 0 -1 43904
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1071_
timestamp 1698431365
transform -1 0 10416 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1072_
timestamp 1698431365
transform 1 0 21728 0 -1 53312
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1073_
timestamp 1698431365
transform 1 0 19824 0 -1 47040
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1074_
timestamp 1698431365
transform -1 0 22176 0 1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1075_
timestamp 1698431365
transform 1 0 7168 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1076_
timestamp 1698431365
transform 1 0 20048 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1077_
timestamp 1698431365
transform -1 0 24864 0 -1 51744
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1078_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29008 0 1 56448
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1079_
timestamp 1698431365
transform 1 0 27888 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1080_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29120 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1081_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 30352 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1082_
timestamp 1698431365
transform 1 0 15568 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1083_
timestamp 1698431365
transform -1 0 16128 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1084_
timestamp 1698431365
transform 1 0 16128 0 1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1085_
timestamp 1698431365
transform -1 0 17920 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1086_
timestamp 1698431365
transform 1 0 15456 0 1 51744
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1087_
timestamp 1698431365
transform 1 0 9856 0 -1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1088_
timestamp 1698431365
transform 1 0 15456 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1089_
timestamp 1698431365
transform 1 0 14448 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1090_
timestamp 1698431365
transform 1 0 25200 0 1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1091_
timestamp 1698431365
transform 1 0 15456 0 1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1092_
timestamp 1698431365
transform 1 0 15008 0 -1 48608
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1093_
timestamp 1698431365
transform -1 0 20160 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1094_
timestamp 1698431365
transform -1 0 23632 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1095_
timestamp 1698431365
transform -1 0 17024 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1096_
timestamp 1698431365
transform -1 0 16352 0 1 42336
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1097_
timestamp 1698431365
transform 1 0 16352 0 1 47040
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1098_
timestamp 1698431365
transform 1 0 21504 0 1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1099_
timestamp 1698431365
transform 1 0 21504 0 1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1100_
timestamp 1698431365
transform 1 0 22512 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1101_
timestamp 1698431365
transform 1 0 20048 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1102_
timestamp 1698431365
transform -1 0 11984 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1103_
timestamp 1698431365
transform -1 0 22624 0 1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1104_
timestamp 1698431365
transform 1 0 23520 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1105_
timestamp 1698431365
transform 1 0 25088 0 -1 42336
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1106_
timestamp 1698431365
transform 1 0 23744 0 -1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1107_
timestamp 1698431365
transform 1 0 24304 0 1 40768
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1108_
timestamp 1698431365
transform 1 0 25088 0 -1 47040
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1109_
timestamp 1698431365
transform 1 0 30016 0 1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1110_
timestamp 1698431365
transform 1 0 23408 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1111_
timestamp 1698431365
transform -1 0 28112 0 1 45472
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1112_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29008 0 1 54880
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1113_
timestamp 1698431365
transform 1 0 27440 0 -1 59584
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1114_
timestamp 1698431365
transform -1 0 19824 0 1 83104
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1115_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 31024 0 -1 83104
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1116_
timestamp 1698431365
transform 1 0 31024 0 1 81536
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1117_
timestamp 1698431365
transform 1 0 29680 0 -1 83104
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1118_
timestamp 1698431365
transform 1 0 21168 0 1 83104
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1119_
timestamp 1698431365
transform 1 0 25088 0 -1 83104
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1120_
timestamp 1698431365
transform -1 0 23184 0 -1 84672
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1121_
timestamp 1698431365
transform -1 0 22848 0 1 86240
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1122_
timestamp 1698431365
transform -1 0 22400 0 -1 87808
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1123_
timestamp 1698431365
transform 1 0 25088 0 1 86240
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1124_
timestamp 1698431365
transform -1 0 25312 0 1 87808
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1125_
timestamp 1698431365
transform -1 0 24080 0 1 89376
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1126_
timestamp 1698431365
transform 1 0 21392 0 1 87808
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1127_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 24080 0 1 89376
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  _1128_
timestamp 1698431365
transform -1 0 38416 0 -1 89376
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _1129_
timestamp 1698431365
transform -1 0 27216 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1130_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 38416 0 1 70560
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1131_
timestamp 1698431365
transform 1 0 25984 0 -1 70560
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1132_
timestamp 1698431365
transform -1 0 27888 0 -1 83104
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1133_
timestamp 1698431365
transform 1 0 26544 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1134_
timestamp 1698431365
transform -1 0 28560 0 1 72128
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1135_
timestamp 1698431365
transform -1 0 26544 0 -1 73696
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1136_
timestamp 1698431365
transform -1 0 29568 0 1 73696
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1137_
timestamp 1698431365
transform 1 0 26544 0 -1 73696
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1138_
timestamp 1698431365
transform -1 0 28672 0 1 70560
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1139_
timestamp 1698431365
transform -1 0 32144 0 1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1140_
timestamp 1698431365
transform 1 0 29344 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _1141_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 30128 0 1 68992
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__and3_2  _1142_
timestamp 1698431365
transform 1 0 30240 0 -1 70560
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1143_
timestamp 1698431365
transform -1 0 34608 0 -1 70560
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1144_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 31920 0 1 70560
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1145_
timestamp 1698431365
transform 1 0 31248 0 1 78400
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1146_
timestamp 1698431365
transform -1 0 31248 0 1 78400
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1147_
timestamp 1698431365
transform -1 0 31920 0 1 70560
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1148_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29456 0 1 79968
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1149_
timestamp 1698431365
transform -1 0 29008 0 -1 81536
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1150_
timestamp 1698431365
transform 1 0 27552 0 1 68992
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1151_
timestamp 1698431365
transform -1 0 31024 0 1 72128
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1152_
timestamp 1698431365
transform 1 0 27888 0 1 81536
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1153_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 27552 0 -1 81536
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1154_
timestamp 1698431365
transform 1 0 28784 0 -1 83104
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1155_
timestamp 1698431365
transform 1 0 29008 0 1 83104
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1156_
timestamp 1698431365
transform -1 0 27888 0 -1 84672
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1157_
timestamp 1698431365
transform 1 0 28448 0 -1 64288
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1158_
timestamp 1698431365
transform -1 0 31584 0 -1 64288
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1159_
timestamp 1698431365
transform 1 0 31024 0 1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1160_
timestamp 1698431365
transform -1 0 30912 0 -1 78400
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1161_
timestamp 1698431365
transform 1 0 29344 0 1 81536
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1162_
timestamp 1698431365
transform 1 0 27888 0 -1 83104
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1163_
timestamp 1698431365
transform 1 0 27552 0 -1 81536
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1164_
timestamp 1698431365
transform 1 0 25536 0 1 78400
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _1165_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 28560 0 1 73696
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1166_
timestamp 1698431365
transform 1 0 27888 0 -1 84672
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1167_
timestamp 1698431365
transform 1 0 29008 0 -1 84672
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1168_
timestamp 1698431365
transform -1 0 23408 0 -1 87808
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1169_
timestamp 1698431365
transform -1 0 23968 0 1 86240
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1170_
timestamp 1698431365
transform -1 0 24640 0 -1 84672
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1171_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 22512 0 1 84672
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1172_
timestamp 1698431365
transform 1 0 23968 0 1 86240
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1173_
timestamp 1698431365
transform 1 0 24864 0 1 95648
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1174_
timestamp 1698431365
transform 1 0 28112 0 -1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1175_
timestamp 1698431365
transform 1 0 29120 0 1 61152
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1176_
timestamp 1698431365
transform 1 0 31920 0 1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1177_
timestamp 1698431365
transform -1 0 29904 0 -1 78400
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1178_
timestamp 1698431365
transform 1 0 29680 0 -1 81536
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1179_
timestamp 1698431365
transform -1 0 29904 0 1 78400
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1180_
timestamp 1698431365
transform -1 0 29456 0 -1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1181_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 28672 0 1 79968
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1182_
timestamp 1698431365
transform 1 0 23184 0 -1 79968
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1183_
timestamp 1698431365
transform 1 0 22400 0 1 89376
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1184_
timestamp 1698431365
transform -1 0 18704 0 -1 79968
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1185_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20944 0 1 79968
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1186_
timestamp 1698431365
transform -1 0 17808 0 1 79968
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1187_
timestamp 1698431365
transform 1 0 23744 0 1 95648
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1188_
timestamp 1698431365
transform 1 0 29008 0 -1 64288
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1189_
timestamp 1698431365
transform 1 0 29456 0 1 62720
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1190_
timestamp 1698431365
transform 1 0 31696 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1191_
timestamp 1698431365
transform -1 0 30800 0 1 75264
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1192_
timestamp 1698431365
transform 1 0 29344 0 -1 76832
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1193_
timestamp 1698431365
transform -1 0 28560 0 1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1194_
timestamp 1698431365
transform -1 0 27552 0 -1 76832
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1195_
timestamp 1698431365
transform 1 0 25088 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1196_
timestamp 1698431365
transform 1 0 26768 0 1 86240
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1197_
timestamp 1698431365
transform -1 0 24640 0 1 78400
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1198_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21616 0 -1 79968
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1199_
timestamp 1698431365
transform -1 0 25984 0 -1 78400
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1200_
timestamp 1698431365
transform 1 0 24640 0 1 78400
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1201_
timestamp 1698431365
transform 1 0 25536 0 1 95648
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1202_
timestamp 1698431365
transform 1 0 29232 0 1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1203_
timestamp 1698431365
transform -1 0 32144 0 -1 59584
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1204_
timestamp 1698431365
transform 1 0 31024 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1205_
timestamp 1698431365
transform 1 0 30912 0 -1 78400
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1206_
timestamp 1698431365
transform 1 0 30688 0 -1 79968
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1207_
timestamp 1698431365
transform -1 0 28784 0 1 78400
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1208_
timestamp 1698431365
transform -1 0 27888 0 1 78400
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1209_
timestamp 1698431365
transform -1 0 26880 0 -1 78400
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1210_
timestamp 1698431365
transform -1 0 26432 0 1 89376
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1211_
timestamp 1698431365
transform 1 0 26768 0 1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1212_
timestamp 1698431365
transform 1 0 26880 0 -1 78400
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1213_
timestamp 1698431365
transform 1 0 26320 0 1 95648
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1214_
timestamp 1698431365
transform 1 0 31696 0 -1 70560
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1215_
timestamp 1698431365
transform -1 0 32368 0 1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1216_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 30240 0 1 65856
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1217_
timestamp 1698431365
transform -1 0 28784 0 -1 68992
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1218_
timestamp 1698431365
transform 1 0 29456 0 -1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1219_
timestamp 1698431365
transform 1 0 26544 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1220_
timestamp 1698431365
transform 1 0 29008 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1221_
timestamp 1698431365
transform 1 0 27216 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1222_
timestamp 1698431365
transform -1 0 28112 0 -1 76832
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1223_
timestamp 1698431365
transform 1 0 24304 0 -1 75264
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1224_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25424 0 -1 72128
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1225_
timestamp 1698431365
transform -1 0 25984 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1226_
timestamp 1698431365
transform 1 0 27664 0 1 86240
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _1227_
timestamp 1698431365
transform 1 0 22288 0 -1 81536
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1228_
timestamp 1698431365
transform -1 0 28560 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1229_
timestamp 1698431365
transform -1 0 30800 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _1230_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 27328 0 -1 58016
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1231_
timestamp 1698431365
transform 1 0 30800 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1232_
timestamp 1698431365
transform -1 0 29344 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_2  _1233_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 28784 0 -1 75264
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1234_
timestamp 1698431365
transform -1 0 28784 0 -1 75264
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1235_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26768 0 1 81536
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1236_
timestamp 1698431365
transform -1 0 24864 0 -1 89376
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1237_
timestamp 1698431365
transform 1 0 25088 0 -1 84672
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1238_
timestamp 1698431365
transform 1 0 29008 0 -1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1239_
timestamp 1698431365
transform -1 0 29344 0 -1 70560
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1240_
timestamp 1698431365
transform 1 0 25088 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1241_
timestamp 1698431365
transform -1 0 22288 0 -1 81536
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1242_
timestamp 1698431365
transform 1 0 25088 0 -1 81536
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1243_
timestamp 1698431365
transform 1 0 23408 0 -1 87808
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1244_
timestamp 1698431365
transform 1 0 20272 0 1 84672
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1245_
timestamp 1698431365
transform -1 0 20944 0 1 86240
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  _1246_
timestamp 1698431365
transform 1 0 4480 0 -1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  _1247_
timestamp 1698431365
transform 1 0 6944 0 1 78400
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1248_
timestamp 1698431365
transform 1 0 6048 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1249_
timestamp 1698431365
transform 1 0 6720 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1250_
timestamp 1698431365
transform 1 0 15904 0 1 3136
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1251_
timestamp 1698431365
transform 1 0 19600 0 -1 3136
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1252_
timestamp 1698431365
transform 1 0 9968 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1253_
timestamp 1698431365
transform -1 0 11200 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1254_
timestamp 1698431365
transform 1 0 12544 0 -1 3136
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1255_
timestamp 1698431365
transform 1 0 12992 0 1 1568
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1256_
timestamp 1698431365
transform 1 0 30912 0 1 3136
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1257_
timestamp 1698431365
transform 1 0 33712 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1258_
timestamp 1698431365
transform 1 0 32928 0 -1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1259_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26768 0 1 3136
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1260_
timestamp 1698431365
transform 1 0 25088 0 -1 3136
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1261_
timestamp 1698431365
transform -1 0 26096 0 -1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1262_
timestamp 1698431365
transform -1 0 14784 0 -1 4704
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1263_
timestamp 1698431365
transform -1 0 10416 0 -1 81536
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1264_
timestamp 1698431365
transform 1 0 10640 0 1 81536
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1265_
timestamp 1698431365
transform 1 0 4704 0 1 81536
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1266_
timestamp 1698431365
transform -1 0 21504 0 -1 84672
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1267_
timestamp 1698431365
transform -1 0 6832 0 1 81536
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1268_
timestamp 1698431365
transform 1 0 5824 0 -1 79968
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1269_
timestamp 1698431365
transform -1 0 20944 0 1 78400
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1270_
timestamp 1698431365
transform -1 0 6720 0 1 78400
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1271_
timestamp 1698431365
transform 1 0 6496 0 1 73696
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1272_
timestamp 1698431365
transform -1 0 23184 0 1 78400
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1273_
timestamp 1698431365
transform -1 0 8400 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1274_
timestamp 1698431365
transform 1 0 5600 0 1 73696
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1275_
timestamp 1698431365
transform -1 0 22288 0 1 78400
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1276_
timestamp 1698431365
transform -1 0 6608 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1277_
timestamp 1698431365
transform -1 0 10864 0 1 78400
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1278_
timestamp 1698431365
transform -1 0 10080 0 -1 78400
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1279_
timestamp 1698431365
transform -1 0 10416 0 -1 76832
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1280_
timestamp 1698431365
transform -1 0 9184 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1281_
timestamp 1698431365
transform -1 0 10416 0 -1 83104
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1282_
timestamp 1698431365
transform -1 0 8624 0 1 83104
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1283_
timestamp 1698431365
transform -1 0 5264 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  _1284_
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1285_
timestamp 1698431365
transform 1 0 8512 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1286_
timestamp 1698431365
transform 1 0 9856 0 -1 3136
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1287_
timestamp 1698431365
transform -1 0 8512 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1288_
timestamp 1698431365
transform -1 0 37744 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1289_
timestamp 1698431365
transform 1 0 36848 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1290_
timestamp 1698431365
transform 1 0 26880 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1291_
timestamp 1698431365
transform 1 0 27552 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1292_
timestamp 1698431365
transform 1 0 28000 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  _1293_
timestamp 1698431365
transform 1 0 11200 0 -1 75264
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1294_
timestamp 1698431365
transform 1 0 29232 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1295_
timestamp 1698431365
transform -1 0 28672 0 1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1296_
timestamp 1698431365
transform -1 0 28112 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1297_
timestamp 1698431365
transform 1 0 26544 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  _1298_
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1299_
timestamp 1698431365
transform -1 0 12768 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1300_
timestamp 1698431365
transform -1 0 11984 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1301_
timestamp 1698431365
transform -1 0 13328 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1302_
timestamp 1698431365
transform 1 0 12320 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1303_
timestamp 1698431365
transform 1 0 15456 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1304_
timestamp 1698431365
transform 1 0 16128 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1305_
timestamp 1698431365
transform 1 0 7280 0 -1 61152
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1306_
timestamp 1698431365
transform 1 0 19040 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1307_
timestamp 1698431365
transform 1 0 19936 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1308_
timestamp 1698431365
transform -1 0 14224 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1309_
timestamp 1698431365
transform 1 0 12432 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1310_
timestamp 1698431365
transform -1 0 10976 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1311_
timestamp 1698431365
transform -1 0 10080 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1312_
timestamp 1698431365
transform -1 0 7280 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1313_
timestamp 1698431365
transform -1 0 6496 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1314_
timestamp 1698431365
transform -1 0 7392 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1315_
timestamp 1698431365
transform 1 0 5824 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1316_
timestamp 1698431365
transform -1 0 10304 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1317_
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1318_
timestamp 1698431365
transform -1 0 12096 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1319_
timestamp 1698431365
transform -1 0 11760 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1320_
timestamp 1698431365
transform -1 0 12096 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1321_
timestamp 1698431365
transform -1 0 10752 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1322_
timestamp 1698431365
transform -1 0 7056 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1323_
timestamp 1698431365
transform -1 0 4368 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1324_
timestamp 1698431365
transform -1 0 4368 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1325_
timestamp 1698431365
transform -1 0 3360 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1326_
timestamp 1698431365
transform -1 0 4144 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1327_
timestamp 1698431365
transform -1 0 3360 0 1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1328_
timestamp 1698431365
transform -1 0 4592 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1329_
timestamp 1698431365
transform -1 0 4816 0 1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1330_
timestamp 1698431365
transform -1 0 6944 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1331_
timestamp 1698431365
transform 1 0 6272 0 1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1332_
timestamp 1698431365
transform 1 0 9408 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1333_
timestamp 1698431365
transform -1 0 10080 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1334_
timestamp 1698431365
transform -1 0 11088 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1335_
timestamp 1698431365
transform -1 0 10528 0 -1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1336_
timestamp 1698431365
transform 1 0 10864 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1337_
timestamp 1698431365
transform -1 0 12096 0 1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1338_
timestamp 1698431365
transform -1 0 14224 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1339_
timestamp 1698431365
transform -1 0 14000 0 1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1340_
timestamp 1698431365
transform 1 0 14448 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1341_
timestamp 1698431365
transform -1 0 16016 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1342_
timestamp 1698431365
transform 1 0 16800 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1343_
timestamp 1698431365
transform 1 0 17360 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1344_
timestamp 1698431365
transform -1 0 22064 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1345_
timestamp 1698431365
transform 1 0 20944 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1346_
timestamp 1698431365
transform 1 0 23072 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1347_
timestamp 1698431365
transform 1 0 23968 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1348_
timestamp 1698431365
transform 1 0 27104 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1349_
timestamp 1698431365
transform -1 0 28672 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1350_
timestamp 1698431365
transform -1 0 31136 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1351_
timestamp 1698431365
transform -1 0 30688 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1352_
timestamp 1698431365
transform 1 0 31472 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1353_
timestamp 1698431365
transform 1 0 32032 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1354_
timestamp 1698431365
transform -1 0 27328 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1355_
timestamp 1698431365
transform 1 0 26880 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1356_
timestamp 1698431365
transform -1 0 26992 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1357_
timestamp 1698431365
transform -1 0 25872 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1358_
timestamp 1698431365
transform -1 0 26096 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1359_
timestamp 1698431365
transform -1 0 25872 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1360_
timestamp 1698431365
transform 1 0 16016 0 -1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1361_
timestamp 1698431365
transform 1 0 17472 0 1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1362_
timestamp 1698431365
transform -1 0 21840 0 1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1363_
timestamp 1698431365
transform -1 0 19712 0 -1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1364_
timestamp 1698431365
transform -1 0 19600 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1365_
timestamp 1698431365
transform -1 0 16800 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1366_
timestamp 1698431365
transform -1 0 7056 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1367_
timestamp 1698431365
transform -1 0 3920 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1368_
timestamp 1698431365
transform -1 0 4368 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1369_
timestamp 1698431365
transform -1 0 3360 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1370_
timestamp 1698431365
transform 1 0 4144 0 -1 68992
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1371_
timestamp 1698431365
transform -1 0 4144 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1372_
timestamp 1698431365
transform -1 0 3360 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1373_
timestamp 1698431365
transform 1 0 4144 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1374_
timestamp 1698431365
transform -1 0 6160 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1375_
timestamp 1698431365
transform -1 0 7280 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1376_
timestamp 1698431365
transform -1 0 7168 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1377_
timestamp 1698431365
transform 1 0 7840 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1378_
timestamp 1698431365
transform -1 0 10080 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1379_
timestamp 1698431365
transform -1 0 8400 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1380_
timestamp 1698431365
transform -1 0 3696 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1381_
timestamp 1698431365
transform -1 0 4368 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1382_
timestamp 1698431365
transform -1 0 3472 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1383_
timestamp 1698431365
transform -1 0 4368 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1384_
timestamp 1698431365
transform 1 0 2128 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1385_
timestamp 1698431365
transform 1 0 5488 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1386_
timestamp 1698431365
transform 1 0 6496 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1387_
timestamp 1698431365
transform 1 0 35056 0 1 54880
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1388_
timestamp 1698431365
transform 1 0 9408 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1389_
timestamp 1698431365
transform 1 0 10416 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1390_
timestamp 1698431365
transform 1 0 15008 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1391_
timestamp 1698431365
transform 1 0 17248 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1392_
timestamp 1698431365
transform 1 0 22288 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1393_
timestamp 1698431365
transform 1 0 23856 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1394_
timestamp 1698431365
transform 1 0 31136 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1395_
timestamp 1698431365
transform 1 0 32928 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1396_
timestamp 1698431365
transform 1 0 35504 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1397_
timestamp 1698431365
transform 1 0 36848 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1398_
timestamp 1698431365
transform 1 0 36848 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1399_
timestamp 1698431365
transform 1 0 36848 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1400_
timestamp 1698431365
transform 1 0 35728 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1401_
timestamp 1698431365
transform 1 0 36848 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1402_
timestamp 1698431365
transform 1 0 30240 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1403_
timestamp 1698431365
transform 1 0 31024 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1404_
timestamp 1698431365
transform 1 0 31136 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1405_
timestamp 1698431365
transform 1 0 31248 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1406_
timestamp 1698431365
transform -1 0 32592 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1407_
timestamp 1698431365
transform 1 0 31136 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1408_
timestamp 1698431365
transform 1 0 35168 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1409_
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1410_
timestamp 1698431365
transform -1 0 37184 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1411_
timestamp 1698431365
transform 1 0 35952 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1412_
timestamp 1698431365
transform -1 0 35728 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1413_
timestamp 1698431365
transform 1 0 34384 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1414_
timestamp 1698431365
transform -1 0 28672 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1415_
timestamp 1698431365
transform -1 0 30352 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1416_
timestamp 1698431365
transform -1 0 30016 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1417_
timestamp 1698431365
transform -1 0 32480 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1418_
timestamp 1698431365
transform 1 0 31024 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1419_
timestamp 1698431365
transform -1 0 37744 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1420_
timestamp 1698431365
transform 1 0 35952 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1421_
timestamp 1698431365
transform 1 0 36848 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1422_
timestamp 1698431365
transform 1 0 36848 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1423_
timestamp 1698431365
transform -1 0 35392 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1424_
timestamp 1698431365
transform -1 0 34160 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1425_
timestamp 1698431365
transform 1 0 23520 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1426_
timestamp 1698431365
transform 1 0 25088 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1427_
timestamp 1698431365
transform 1 0 25760 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1428_
timestamp 1698431365
transform 1 0 26656 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1429_
timestamp 1698431365
transform 1 0 30016 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1430_
timestamp 1698431365
transform 1 0 30688 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1431_
timestamp 1698431365
transform -1 0 33824 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1432_
timestamp 1698431365
transform -1 0 33712 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1433_
timestamp 1698431365
transform 1 0 35168 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1434_
timestamp 1698431365
transform 1 0 35840 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1435_
timestamp 1698431365
transform -1 0 37744 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1436_
timestamp 1698431365
transform 1 0 36848 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1437_
timestamp 1698431365
transform 1 0 11648 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1438_
timestamp 1698431365
transform -1 0 14000 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1439_
timestamp 1698431365
transform -1 0 11984 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1440_
timestamp 1698431365
transform 1 0 10416 0 -1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1441_
timestamp 1698431365
transform -1 0 8624 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1442_
timestamp 1698431365
transform -1 0 7616 0 -1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1443_
timestamp 1698431365
transform -1 0 9184 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1444_
timestamp 1698431365
transform -1 0 8400 0 1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1445_
timestamp 1698431365
transform -1 0 10304 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1446_
timestamp 1698431365
transform -1 0 4032 0 -1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1447_
timestamp 1698431365
transform -1 0 6384 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1448_
timestamp 1698431365
transform 1 0 5488 0 1 70560
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1449_
timestamp 1698431365
transform 1 0 8400 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1450_
timestamp 1698431365
transform -1 0 9072 0 -1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1451_
timestamp 1698431365
transform 1 0 9968 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1452_
timestamp 1698431365
transform 1 0 11088 0 1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1453_
timestamp 1698431365
transform 1 0 15456 0 -1 70560
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1454_
timestamp 1698431365
transform 1 0 18032 0 -1 70560
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1455_
timestamp 1698431365
transform 1 0 20384 0 1 67424
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1456_
timestamp 1698431365
transform 1 0 21168 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1457_
timestamp 1698431365
transform -1 0 23072 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1458_
timestamp 1698431365
transform 1 0 20720 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1459_
timestamp 1698431365
transform -1 0 19376 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1460_
timestamp 1698431365
transform -1 0 16240 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1461_
timestamp 1698431365
transform 1 0 30464 0 1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1462_
timestamp 1698431365
transform -1 0 15008 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1463_
timestamp 1698431365
transform -1 0 14000 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1464_
timestamp 1698431365
transform -1 0 15568 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1465_
timestamp 1698431365
transform 1 0 14896 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1466_
timestamp 1698431365
transform 1 0 17696 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1467_
timestamp 1698431365
transform -1 0 19152 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1468_
timestamp 1698431365
transform 1 0 5600 0 -1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1469_
timestamp 1698431365
transform -1 0 22064 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1470_
timestamp 1698431365
transform 1 0 20944 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1471_
timestamp 1698431365
transform 1 0 22064 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1472_
timestamp 1698431365
transform -1 0 22960 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1473_
timestamp 1698431365
transform -1 0 24304 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1474_
timestamp 1698431365
transform 1 0 22960 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1475_
timestamp 1698431365
transform -1 0 24976 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1476_
timestamp 1698431365
transform -1 0 24640 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1477_
timestamp 1698431365
transform 1 0 25984 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1478_
timestamp 1698431365
transform 1 0 26432 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1479_
timestamp 1698431365
transform -1 0 31696 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1480_
timestamp 1698431365
transform 1 0 30352 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1481_
timestamp 1698431365
transform -1 0 31920 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1482_
timestamp 1698431365
transform 1 0 30912 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1483_
timestamp 1698431365
transform -1 0 26656 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1484_
timestamp 1698431365
transform -1 0 26432 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1485_
timestamp 1698431365
transform -1 0 21504 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1486_
timestamp 1698431365
transform -1 0 11200 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1487_
timestamp 1698431365
transform -1 0 5040 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1488_
timestamp 1698431365
transform -1 0 3472 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1489_
timestamp 1698431365
transform -1 0 4368 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1490_
timestamp 1698431365
transform -1 0 3472 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1491_
timestamp 1698431365
transform 1 0 5824 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1492_
timestamp 1698431365
transform 1 0 6832 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1493_
timestamp 1698431365
transform 1 0 9408 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1494_
timestamp 1698431365
transform 1 0 9968 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1495_
timestamp 1698431365
transform -1 0 13328 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1496_
timestamp 1698431365
transform -1 0 12880 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1497_
timestamp 1698431365
transform -1 0 14224 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1498_
timestamp 1698431365
transform -1 0 12656 0 -1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1499_
timestamp 1698431365
transform -1 0 14560 0 1 64288
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1500_
timestamp 1698431365
transform 1 0 13328 0 1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1501_
timestamp 1698431365
transform -1 0 14896 0 1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1502_
timestamp 1698431365
transform -1 0 14896 0 1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1503_
timestamp 1698431365
transform 1 0 13328 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1504_
timestamp 1698431365
transform 1 0 14000 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1505_
timestamp 1698431365
transform -1 0 14896 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1506_
timestamp 1698431365
transform -1 0 14000 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1507_
timestamp 1698431365
transform 1 0 14112 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1508_
timestamp 1698431365
transform -1 0 15680 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1509_
timestamp 1698431365
transform -1 0 17024 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1510_
timestamp 1698431365
transform 1 0 15232 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1511_
timestamp 1698431365
transform -1 0 18368 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1512_
timestamp 1698431365
transform 1 0 17248 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1513_
timestamp 1698431365
transform -1 0 16576 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1514_
timestamp 1698431365
transform 1 0 14560 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1515_
timestamp 1698431365
transform -1 0 10304 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1516_
timestamp 1698431365
transform 1 0 7840 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1517_
timestamp 1698431365
transform -1 0 6384 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1518_
timestamp 1698431365
transform -1 0 4480 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1519_
timestamp 1698431365
transform -1 0 5488 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1520_
timestamp 1698431365
transform -1 0 4368 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1521_
timestamp 1698431365
transform 1 0 5600 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1522_
timestamp 1698431365
transform 1 0 6496 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1523_
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1524_
timestamp 1698431365
transform 1 0 9520 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1525_
timestamp 1698431365
transform 1 0 12880 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1526_
timestamp 1698431365
transform 1 0 13440 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1527_
timestamp 1698431365
transform 1 0 18144 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1528_
timestamp 1698431365
transform 1 0 20272 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1529_
timestamp 1698431365
transform 1 0 25984 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1530_
timestamp 1698431365
transform 1 0 26880 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1531_
timestamp 1698431365
transform 1 0 30128 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1532_
timestamp 1698431365
transform -1 0 31696 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1533_
timestamp 1698431365
transform 1 0 31696 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1534_
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1535_
timestamp 1698431365
transform -1 0 30016 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1536_
timestamp 1698431365
transform -1 0 28112 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1537_
timestamp 1698431365
transform -1 0 26320 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1538_
timestamp 1698431365
transform 1 0 24192 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1539_
timestamp 1698431365
transform 1 0 26880 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1540_
timestamp 1698431365
transform 1 0 27664 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1541_
timestamp 1698431365
transform 1 0 30688 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1542_
timestamp 1698431365
transform -1 0 32256 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1543_
timestamp 1698431365
transform -1 0 34384 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1544_
timestamp 1698431365
transform 1 0 33264 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1545_
timestamp 1698431365
transform 1 0 34496 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1546_
timestamp 1698431365
transform 1 0 36848 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1547_
timestamp 1698431365
transform -1 0 33824 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1548_
timestamp 1698431365
transform -1 0 32032 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1549_
timestamp 1698431365
transform -1 0 22624 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1550_
timestamp 1698431365
transform 1 0 21616 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1551_
timestamp 1698431365
transform -1 0 22176 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1552_
timestamp 1698431365
transform -1 0 21168 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1553_
timestamp 1698431365
transform 1 0 19936 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1554_
timestamp 1698431365
transform 1 0 20048 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1555_
timestamp 1698431365
transform -1 0 20832 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1556_
timestamp 1698431365
transform 1 0 19152 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1557_
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1558_
timestamp 1698431365
transform -1 0 22736 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1559_
timestamp 1698431365
transform 1 0 22064 0 -1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1560_
timestamp 1698431365
transform 1 0 21728 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1561_
timestamp 1698431365
transform 1 0 22064 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1562_
timestamp 1698431365
transform -1 0 22064 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1563_
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1564_
timestamp 1698431365
transform 1 0 21728 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1565_
timestamp 1698431365
transform 1 0 22176 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1566_
timestamp 1698431365
transform -1 0 24640 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1567_
timestamp 1698431365
transform 1 0 23296 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1568_
timestamp 1698431365
transform -1 0 25984 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1569_
timestamp 1698431365
transform 1 0 24192 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1570_
timestamp 1698431365
transform -1 0 27776 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1571_
timestamp 1698431365
transform 1 0 25312 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1572_
timestamp 1698431365
transform -1 0 28224 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1573_
timestamp 1698431365
transform 1 0 27552 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1574_
timestamp 1698431365
transform 1 0 26656 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1575_
timestamp 1698431365
transform 1 0 26880 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1576_
timestamp 1698431365
transform -1 0 29904 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1577_
timestamp 1698431365
transform 1 0 29120 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1578_
timestamp 1698431365
transform 1 0 30800 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1579_
timestamp 1698431365
transform -1 0 33600 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1580_
timestamp 1698431365
transform 1 0 34832 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1581_
timestamp 1698431365
transform 1 0 36176 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1582_
timestamp 1698431365
transform 1 0 35392 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1583_
timestamp 1698431365
transform 1 0 35616 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1584_
timestamp 1698431365
transform 1 0 35392 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1585_
timestamp 1698431365
transform -1 0 36288 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1586_
timestamp 1698431365
transform 1 0 23184 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1587_
timestamp 1698431365
transform 1 0 24080 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1588_
timestamp 1698431365
transform -1 0 24640 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1589_
timestamp 1698431365
transform 1 0 23408 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1590_
timestamp 1698431365
transform -1 0 23744 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1591_
timestamp 1698431365
transform -1 0 23184 0 -1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1592_
timestamp 1698431365
transform 1 0 25088 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1593_
timestamp 1698431365
transform 1 0 25088 0 1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1594_
timestamp 1698431365
transform 1 0 25312 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1595_
timestamp 1698431365
transform 1 0 25424 0 -1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1596_
timestamp 1698431365
transform -1 0 24864 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1597_
timestamp 1698431365
transform 1 0 24080 0 -1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1598_
timestamp 1698431365
transform 1 0 23968 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1599_
timestamp 1698431365
transform -1 0 24528 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1600_
timestamp 1698431365
transform -1 0 8512 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1601_
timestamp 1698431365
transform -1 0 5488 0 -1 10976
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1602_
timestamp 1698431365
transform -1 0 5600 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1603_
timestamp 1698431365
transform -1 0 3808 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1604_
timestamp 1698431365
transform -1 0 4592 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1605_
timestamp 1698431365
transform -1 0 3808 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1606_
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1607_
timestamp 1698431365
transform -1 0 7056 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1608_
timestamp 1698431365
transform 1 0 8288 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1609_
timestamp 1698431365
transform -1 0 10080 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1610_
timestamp 1698431365
transform -1 0 12544 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1611_
timestamp 1698431365
transform -1 0 12096 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1612_
timestamp 1698431365
transform -1 0 12208 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1613_
timestamp 1698431365
transform -1 0 10864 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1614_
timestamp 1698431365
transform -1 0 10640 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1615_
timestamp 1698431365
transform -1 0 10080 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1616_
timestamp 1698431365
transform -1 0 10304 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1617_
timestamp 1698431365
transform -1 0 9072 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1618_
timestamp 1698431365
transform -1 0 11200 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1619_
timestamp 1698431365
transform 1 0 9744 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1620_
timestamp 1698431365
transform -1 0 12544 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1621_
timestamp 1698431365
transform -1 0 12432 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1622_
timestamp 1698431365
transform -1 0 14224 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1623_
timestamp 1698431365
transform -1 0 14000 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1624_
timestamp 1698431365
transform -1 0 15792 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1625_
timestamp 1698431365
transform -1 0 14672 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1626_
timestamp 1698431365
transform -1 0 14784 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1627_
timestamp 1698431365
transform -1 0 14784 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1628_
timestamp 1698431365
transform -1 0 16128 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1629_
timestamp 1698431365
transform -1 0 16352 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1630_
timestamp 1698431365
transform -1 0 18144 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1631_
timestamp 1698431365
transform -1 0 17920 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1632_
timestamp 1698431365
transform -1 0 18480 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1633_
timestamp 1698431365
transform 1 0 17696 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1634_
timestamp 1698431365
transform 1 0 17808 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1635_
timestamp 1698431365
transform -1 0 20160 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1636_
timestamp 1698431365
transform -1 0 6384 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1637_
timestamp 1698431365
transform -1 0 4256 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1638_
timestamp 1698431365
transform -1 0 4592 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1639_
timestamp 1698431365
transform -1 0 3584 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1640_
timestamp 1698431365
transform -1 0 5712 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1641_
timestamp 1698431365
transform -1 0 4032 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1642_
timestamp 1698431365
transform -1 0 7392 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1643_
timestamp 1698431365
transform 1 0 6272 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1644_
timestamp 1698431365
transform -1 0 8736 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1645_
timestamp 1698431365
transform -1 0 7952 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1646_
timestamp 1698431365
transform -1 0 8176 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1647_
timestamp 1698431365
transform -1 0 7280 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1648_
timestamp 1698431365
transform -1 0 5488 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1649_
timestamp 1698431365
transform -1 0 4256 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1650_
timestamp 1698431365
transform -1 0 4704 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1651_
timestamp 1698431365
transform -1 0 3472 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1652_
timestamp 1698431365
transform 1 0 4368 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1653_
timestamp 1698431365
transform -1 0 5488 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1654_
timestamp 1698431365
transform 1 0 6944 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1655_
timestamp 1698431365
transform 1 0 7504 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1656_
timestamp 1698431365
transform 1 0 9744 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1657_
timestamp 1698431365
transform 1 0 10528 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1658_
timestamp 1698431365
transform -1 0 18144 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1659_
timestamp 1698431365
transform 1 0 16352 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1660_
timestamp 1698431365
transform -1 0 20608 0 -1 84672
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1661_
timestamp 1698431365
transform -1 0 19040 0 -1 83104
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1662_
timestamp 1698431365
transform 1 0 16240 0 1 79968
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1663_
timestamp 1698431365
transform -1 0 17024 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1664_
timestamp 1698431365
transform -1 0 18144 0 -1 78400
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1665_
timestamp 1698431365
transform -1 0 15344 0 1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1666_
timestamp 1698431365
transform 1 0 14448 0 1 78400
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1667_
timestamp 1698431365
transform 1 0 13552 0 1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1668_
timestamp 1698431365
transform 1 0 12208 0 1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1669_
timestamp 1698431365
transform -1 0 18144 0 -1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1670_
timestamp 1698431365
transform 1 0 17248 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1671_
timestamp 1698431365
transform 1 0 19712 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1672_
timestamp 1698431365
transform 1 0 17808 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1673_
timestamp 1698431365
transform -1 0 23296 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1674_
timestamp 1698431365
transform 1 0 23296 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1675_
timestamp 1698431365
transform 1 0 20496 0 -1 81536
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1676_
timestamp 1698431365
transform -1 0 19488 0 -1 84672
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1677_
timestamp 1698431365
transform -1 0 20048 0 1 87808
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1678_
timestamp 1698431365
transform -1 0 18704 0 1 83104
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1679_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 13776 0 -1 81536
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1680_
timestamp 1698431365
transform -1 0 12656 0 1 78400
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1681_
timestamp 1698431365
transform -1 0 12096 0 1 79968
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1682_
timestamp 1698431365
transform 1 0 13664 0 1 81536
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1683_
timestamp 1698431365
transform 1 0 15008 0 1 83104
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1684_
timestamp 1698431365
transform -1 0 14672 0 -1 86240
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1685_
timestamp 1698431365
transform -1 0 14448 0 1 84672
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1686_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 16016 0 1 87808
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1687_
timestamp 1698431365
transform -1 0 14560 0 1 87808
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1688_
timestamp 1698431365
transform 1 0 15456 0 -1 87808
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1689_
timestamp 1698431365
transform -1 0 18032 0 1 86240
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1690_
timestamp 1698431365
transform -1 0 17024 0 -1 89376
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1691_
timestamp 1698431365
transform -1 0 27776 0 1 89376
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1692_
timestamp 1698431365
transform -1 0 24864 0 -1 87808
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1693_
timestamp 1698431365
transform -1 0 31024 0 1 89376
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1694_
timestamp 1698431365
transform -1 0 30464 0 -1 90944
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1695_
timestamp 1698431365
transform 1 0 31136 0 -1 86240
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1696_
timestamp 1698431365
transform 1 0 31472 0 1 84672
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1697_
timestamp 1698431365
transform 1 0 32368 0 1 84672
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1698_
timestamp 1698431365
transform -1 0 33824 0 -1 87808
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1699_
timestamp 1698431365
transform 1 0 34608 0 -1 86240
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1700_
timestamp 1698431365
transform -1 0 35840 0 1 87808
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1701_
timestamp 1698431365
transform 1 0 35728 0 1 84672
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1702_
timestamp 1698431365
transform 1 0 35056 0 1 83104
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1703_
timestamp 1698431365
transform 1 0 36848 0 1 83104
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1704_
timestamp 1698431365
transform -1 0 37856 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1705_
timestamp 1698431365
transform -1 0 35056 0 1 83104
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1706_
timestamp 1698431365
transform 1 0 35168 0 1 84672
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1707_
timestamp 1698431365
transform 1 0 36064 0 -1 86240
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1708_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 10640 0 1 81536
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1709_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 6832 0 -1 81536
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1710_
timestamp 1698431365
transform -1 0 6720 0 -1 78400
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1711_
timestamp 1698431365
transform -1 0 7504 0 -1 75264
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1712_
timestamp 1698431365
transform -1 0 5264 0 1 73696
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1713_
timestamp 1698431365
transform -1 0 10416 0 1 76832
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1714_
timestamp 1698431365
transform -1 0 10752 0 1 75264
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1715_
timestamp 1698431365
transform -1 0 9184 0 -1 83104
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1716_
timestamp 1698431365
transform -1 0 8736 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1717_
timestamp 1698431365
transform -1 0 38416 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1718_
timestamp 1698431365
transform 1 0 25536 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1719_
timestamp 1698431365
transform 1 0 26656 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1720_
timestamp 1698431365
transform 1 0 27104 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1721_
timestamp 1698431365
transform 1 0 29008 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1722_
timestamp 1698431365
transform 1 0 26544 0 -1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1723_
timestamp 1698431365
transform -1 0 28336 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1724_
timestamp 1698431365
transform 1 0 9856 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1725_
timestamp 1698431365
transform 1 0 11648 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1726_
timestamp 1698431365
transform 1 0 15792 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1727_
timestamp 1698431365
transform -1 0 21504 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1728_
timestamp 1698431365
transform -1 0 14448 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1729_
timestamp 1698431365
transform -1 0 11088 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1730_
timestamp 1698431365
transform 1 0 4480 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1731_
timestamp 1698431365
transform 1 0 5488 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1732_
timestamp 1698431365
transform 1 0 8960 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1733_
timestamp 1698431365
transform 1 0 9856 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1734_
timestamp 1698431365
transform -1 0 11424 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1735_
timestamp 1698431365
transform 1 0 1792 0 1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1736_
timestamp 1698431365
transform 1 0 1568 0 1 59584
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1737_
timestamp 1698431365
transform 1 0 1568 0 -1 67424
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1738_
timestamp 1698431365
transform 1 0 2688 0 -1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1739_
timestamp 1698431365
transform 1 0 5600 0 -1 62720
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1740_
timestamp 1698431365
transform 1 0 8176 0 1 58016
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1741_
timestamp 1698431365
transform 1 0 8848 0 1 62720
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1742_
timestamp 1698431365
transform 1 0 9856 0 1 70560
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1743_
timestamp 1698431365
transform 1 0 11760 0 -1 70560
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1744_
timestamp 1698431365
transform 1 0 13776 0 1 58016
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1745_
timestamp 1698431365
transform 1 0 17248 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1746_
timestamp 1698431365
transform 1 0 21168 0 1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1747_
timestamp 1698431365
transform 1 0 23856 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1748_
timestamp 1698431365
transform 1 0 27216 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1749_
timestamp 1698431365
transform 1 0 29456 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1750_
timestamp 1698431365
transform -1 0 33600 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1751_
timestamp 1698431365
transform -1 0 28672 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1752_
timestamp 1698431365
transform 1 0 23744 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1753_
timestamp 1698431365
transform 1 0 24304 0 1 62720
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1754_
timestamp 1698431365
transform 1 0 14672 0 1 68992
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1755_
timestamp 1698431365
transform 1 0 17248 0 -1 68992
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1756_
timestamp 1698431365
transform 1 0 17696 0 1 62720
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1757_
timestamp 1698431365
transform 1 0 17696 0 1 58016
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1758_
timestamp 1698431365
transform -1 0 16128 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1759_
timestamp 1698431365
transform 1 0 1568 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1760_
timestamp 1698431365
transform 1 0 1568 0 -1 58016
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1761_
timestamp 1698431365
transform 1 0 1568 0 -1 62720
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1762_
timestamp 1698431365
transform 1 0 3696 0 -1 59584
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1763_
timestamp 1698431365
transform 1 0 5600 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1764_
timestamp 1698431365
transform 1 0 5936 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1765_
timestamp 1698431365
transform 1 0 1568 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1766_
timestamp 1698431365
transform 1 0 1568 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1767_
timestamp 1698431365
transform 1 0 2016 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1768_
timestamp 1698431365
transform 1 0 6384 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1769_
timestamp 1698431365
transform 1 0 9856 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1770_
timestamp 1698431365
transform 1 0 17472 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1771_
timestamp 1698431365
transform 1 0 25088 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1772_
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1773_
timestamp 1698431365
transform -1 0 38416 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1774_
timestamp 1698431365
transform -1 0 38416 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1775_
timestamp 1698431365
transform -1 0 38416 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1776_
timestamp 1698431365
transform -1 0 32704 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1777_
timestamp 1698431365
transform -1 0 33488 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1778_
timestamp 1698431365
transform 1 0 31808 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1779_
timestamp 1698431365
transform -1 0 38416 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1780_
timestamp 1698431365
transform -1 0 38416 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1781_
timestamp 1698431365
transform -1 0 36176 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1782_
timestamp 1698431365
transform 1 0 27328 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1783_
timestamp 1698431365
transform 1 0 28336 0 -1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1784_
timestamp 1698431365
transform 1 0 31696 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1785_
timestamp 1698431365
transform -1 0 38416 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1786_
timestamp 1698431365
transform -1 0 38416 0 -1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1787_
timestamp 1698431365
transform -1 0 34832 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1788_
timestamp 1698431365
transform -1 0 28000 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1789_
timestamp 1698431365
transform 1 0 26768 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1790_
timestamp 1698431365
transform 1 0 30352 0 1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1791_
timestamp 1698431365
transform 1 0 32256 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1792_
timestamp 1698431365
transform 1 0 35168 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1793_
timestamp 1698431365
transform -1 0 38416 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1794_
timestamp 1698431365
transform 1 0 9856 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1795_
timestamp 1698431365
transform -1 0 12208 0 1 59584
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1796_
timestamp 1698431365
transform 1 0 5600 0 1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1797_
timestamp 1698431365
transform 1 0 5936 0 -1 68992
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1798_
timestamp 1698431365
transform 1 0 2016 0 1 68992
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1799_
timestamp 1698431365
transform 1 0 5264 0 -1 70560
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1800_
timestamp 1698431365
transform 1 0 6608 0 1 70560
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1801_
timestamp 1698431365
transform 1 0 10864 0 -1 72128
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1802_
timestamp 1698431365
transform 1 0 14784 0 1 70560
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1803_
timestamp 1698431365
transform 1 0 18704 0 -1 70560
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1804_
timestamp 1698431365
transform 1 0 19824 0 -1 67424
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1805_
timestamp 1698431365
transform 1 0 21168 0 1 58016
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1806_
timestamp 1698431365
transform -1 0 22624 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1807_
timestamp 1698431365
transform -1 0 16464 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1808_
timestamp 1698431365
transform 1 0 11872 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1809_
timestamp 1698431365
transform 1 0 14336 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1810_
timestamp 1698431365
transform 1 0 17696 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1811_
timestamp 1698431365
transform -1 0 24416 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1812_
timestamp 1698431365
transform 1 0 21392 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1813_
timestamp 1698431365
transform 1 0 22512 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1814_
timestamp 1698431365
transform 1 0 22960 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1815_
timestamp 1698431365
transform 1 0 27104 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1816_
timestamp 1698431365
transform -1 0 32256 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1817_
timestamp 1698431365
transform -1 0 33376 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1818_
timestamp 1698431365
transform -1 0 26880 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1819_
timestamp 1698431365
transform -1 0 10528 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1820_
timestamp 1698431365
transform 1 0 1568 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1821_
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1822_
timestamp 1698431365
transform 1 0 6608 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1823_
timestamp 1698431365
transform 1 0 9744 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1824_
timestamp 1698431365
transform 1 0 11200 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1825_
timestamp 1698431365
transform 1 0 10752 0 -1 59584
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1826_
timestamp 1698431365
transform 1 0 11200 0 -1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1827_
timestamp 1698431365
transform 1 0 11536 0 -1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1828_
timestamp 1698431365
transform 1 0 13328 0 1 59584
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1829_
timestamp 1698431365
transform 1 0 12096 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1830_
timestamp 1698431365
transform 1 0 11424 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1831_
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1832_
timestamp 1698431365
transform 1 0 11984 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1833_
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1834_
timestamp 1698431365
transform 1 0 15680 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1835_
timestamp 1698431365
transform -1 0 19040 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1836_
timestamp 1698431365
transform -1 0 16576 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1837_
timestamp 1698431365
transform -1 0 9408 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1838_
timestamp 1698431365
transform 1 0 1680 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1839_
timestamp 1698431365
transform 1 0 2352 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1840_
timestamp 1698431365
transform 1 0 5824 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1841_
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1842_
timestamp 1698431365
transform 1 0 13216 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1843_
timestamp 1698431365
transform 1 0 21168 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1844_
timestamp 1698431365
transform 1 0 26880 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1845_
timestamp 1698431365
transform 1 0 29568 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1846_
timestamp 1698431365
transform -1 0 36064 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1847_
timestamp 1698431365
transform -1 0 28336 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1848_
timestamp 1698431365
transform 1 0 24080 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1849_
timestamp 1698431365
transform 1 0 27440 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1850_
timestamp 1698431365
transform 1 0 30240 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1851_
timestamp 1698431365
transform 1 0 32928 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1852_
timestamp 1698431365
transform -1 0 38416 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1853_
timestamp 1698431365
transform -1 0 32704 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1854_
timestamp 1698431365
transform -1 0 23632 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1855_
timestamp 1698431365
transform -1 0 20944 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1856_
timestamp 1698431365
transform -1 0 22176 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1857_
timestamp 1698431365
transform 1 0 18704 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1858_
timestamp 1698431365
transform -1 0 23072 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1859_
timestamp 1698431365
transform -1 0 23968 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1860_
timestamp 1698431365
transform -1 0 22848 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1861_
timestamp 1698431365
transform 1 0 21616 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1862_
timestamp 1698431365
transform 1 0 22960 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1863_
timestamp 1698431365
transform 1 0 23968 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1864_
timestamp 1698431365
transform 1 0 25200 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1865_
timestamp 1698431365
transform -1 0 29904 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1866_
timestamp 1698431365
transform -1 0 28784 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1867_
timestamp 1698431365
transform 1 0 28784 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1868_
timestamp 1698431365
transform 1 0 31696 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1869_
timestamp 1698431365
transform -1 0 38416 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1870_
timestamp 1698431365
transform -1 0 37968 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1871_
timestamp 1698431365
transform 1 0 34832 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1872_
timestamp 1698431365
transform -1 0 25312 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1873_
timestamp 1698431365
transform -1 0 25200 0 1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1874_
timestamp 1698431365
transform 1 0 21840 0 1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1875_
timestamp 1698431365
transform -1 0 27216 0 1 67424
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1876_
timestamp 1698431365
transform -1 0 27552 0 1 61152
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1877_
timestamp 1698431365
transform -1 0 28448 0 1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1878_
timestamp 1698431365
transform -1 0 26208 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1879_
timestamp 1698431365
transform -1 0 9184 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1880_
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1881_
timestamp 1698431365
transform 1 0 2016 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1882_
timestamp 1698431365
transform 1 0 5152 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1883_
timestamp 1698431365
transform 1 0 8400 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1884_
timestamp 1698431365
transform 1 0 10640 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1885_
timestamp 1698431365
transform 1 0 8400 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1886_
timestamp 1698431365
transform 1 0 7392 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1887_
timestamp 1698431365
transform 1 0 7056 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1888_
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1889_
timestamp 1698431365
transform 1 0 10976 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1890_
timestamp 1698431365
transform 1 0 11648 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1891_
timestamp 1698431365
transform 1 0 12992 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1892_
timestamp 1698431365
transform 1 0 12768 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1893_
timestamp 1698431365
transform 1 0 14784 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1894_
timestamp 1698431365
transform 1 0 16128 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1895_
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1896_
timestamp 1698431365
transform -1 0 19488 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1897_
timestamp 1698431365
transform 1 0 1680 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1898_
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1899_
timestamp 1698431365
transform 1 0 2240 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1900_
timestamp 1698431365
transform 1 0 5936 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1901_
timestamp 1698431365
transform 1 0 5936 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1902_
timestamp 1698431365
transform 1 0 5824 0 -1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1903_
timestamp 1698431365
transform 1 0 2016 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1904_
timestamp 1698431365
transform 1 0 1568 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1905_
timestamp 1698431365
transform 1 0 3696 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1906_
timestamp 1698431365
transform 1 0 7056 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1907_
timestamp 1698431365
transform 1 0 9856 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1908_
timestamp 1698431365
transform 1 0 16800 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1909_
timestamp 1698431365
transform 1 0 16016 0 1 78400
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1910_
timestamp 1698431365
transform 1 0 13104 0 -1 78400
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1911_
timestamp 1698431365
transform 1 0 11312 0 -1 76832
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1912_
timestamp 1698431365
transform -1 0 17024 0 -1 73696
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1913_
timestamp 1698431365
transform 1 0 18816 0 -1 75264
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1914_
timestamp 1698431365
transform 1 0 21616 0 -1 72128
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1915_
timestamp 1698431365
transform 1 0 17248 0 -1 81536
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1916_
timestamp 1698431365
transform 1 0 17360 0 -1 89376
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1917_
timestamp 1698431365
transform 1 0 17248 0 1 81536
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1918_
timestamp 1698431365
transform 1 0 10416 0 -1 79968
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1919_
timestamp 1698431365
transform 1 0 11760 0 -1 83104
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1920_
timestamp 1698431365
transform -1 0 15680 0 -1 84672
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1921_
timestamp 1698431365
transform 1 0 13104 0 -1 89376
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1922_
timestamp 1698431365
transform 1 0 16016 0 1 87808
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1923_
timestamp 1698431365
transform -1 0 28784 0 1 87808
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1924_
timestamp 1698431365
transform 1 0 29008 0 1 87808
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1925_
timestamp 1698431365
transform -1 0 32704 0 1 86240
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1926_
timestamp 1698431365
transform -1 0 35952 0 1 86240
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1927_
timestamp 1698431365
transform 1 0 34720 0 -1 87808
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1928_
timestamp 1698431365
transform 1 0 35168 0 -1 84672
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1929_
timestamp 1698431365
transform 1 0 34832 0 -1 83104
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0842__I open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 36176 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0843__I
timestamp 1698431365
transform 1 0 30800 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0846__I
timestamp 1698431365
transform -1 0 24528 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0848__A2
timestamp 1698431365
transform -1 0 17024 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0849__A1
timestamp 1698431365
transform -1 0 13104 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0849__A2
timestamp 1698431365
transform 1 0 16128 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0849__A3
timestamp 1698431365
transform 1 0 16576 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0850__A1
timestamp 1698431365
transform 1 0 15568 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0851__A1
timestamp 1698431365
transform 1 0 17472 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0851__A2
timestamp 1698431365
transform 1 0 19152 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0855__A1
timestamp 1698431365
transform -1 0 37744 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0855__A2
timestamp 1698431365
transform 1 0 37072 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0858__I
timestamp 1698431365
transform 1 0 19040 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0859__A1
timestamp 1698431365
transform 1 0 30016 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0859__A2
timestamp 1698431365
transform 1 0 31360 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0862__I
timestamp 1698431365
transform 1 0 23856 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0863__I
timestamp 1698431365
transform 1 0 31808 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0866__A1
timestamp 1698431365
transform 1 0 25760 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0866__A2
timestamp 1698431365
transform 1 0 19040 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0866__A3
timestamp 1698431365
transform 1 0 20720 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0869__A1
timestamp 1698431365
transform 1 0 16800 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0869__A2
timestamp 1698431365
transform 1 0 15120 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0870__A1
timestamp 1698431365
transform 1 0 15904 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0871__I
timestamp 1698431365
transform 1 0 21392 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0872__A1
timestamp 1698431365
transform 1 0 31360 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0872__A2
timestamp 1698431365
transform -1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0872__A3
timestamp 1698431365
transform 1 0 23296 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0872__A4
timestamp 1698431365
transform 1 0 24192 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0873__A1
timestamp 1698431365
transform 1 0 28000 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0874__I
timestamp 1698431365
transform -1 0 14896 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0876__A1
timestamp 1698431365
transform 1 0 23632 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0876__A2
timestamp 1698431365
transform 1 0 18144 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0876__A3
timestamp 1698431365
transform 1 0 18592 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0876__A4
timestamp 1698431365
transform 1 0 23184 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0877__A1
timestamp 1698431365
transform 1 0 25312 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0877__A2
timestamp 1698431365
transform 1 0 23856 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0878__A2
timestamp 1698431365
transform 1 0 29232 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0878__B1
timestamp 1698431365
transform 1 0 29680 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0879__A1
timestamp 1698431365
transform 1 0 32256 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0880__A1
timestamp 1698431365
transform 1 0 22512 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0880__A2
timestamp 1698431365
transform 1 0 22064 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0881__A1
timestamp 1698431365
transform 1 0 26656 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0881__A2
timestamp 1698431365
transform 1 0 22064 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0882__A1
timestamp 1698431365
transform 1 0 31696 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0882__A2
timestamp 1698431365
transform 1 0 32368 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0882__A3
timestamp 1698431365
transform 1 0 31920 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0883__B1
timestamp 1698431365
transform 1 0 30240 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0884__A1
timestamp 1698431365
transform 1 0 15232 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0884__A2
timestamp 1698431365
transform -1 0 15456 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0885__A1
timestamp 1698431365
transform 1 0 24640 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0885__A2
timestamp 1698431365
transform 1 0 26992 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0885__A3
timestamp 1698431365
transform -1 0 14000 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0886__A1
timestamp 1698431365
transform 1 0 19264 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0886__A2
timestamp 1698431365
transform 1 0 17920 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0887__A1
timestamp 1698431365
transform 1 0 16800 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0888__A2
timestamp 1698431365
transform 1 0 30688 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0888__B1
timestamp 1698431365
transform 1 0 31136 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0889__I
timestamp 1698431365
transform 1 0 21616 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0890__A1
timestamp 1698431365
transform -1 0 22624 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0890__A2
timestamp 1698431365
transform -1 0 22176 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0890__A3
timestamp 1698431365
transform 1 0 24416 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0890__A4
timestamp 1698431365
transform 1 0 22848 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0891__A1
timestamp 1698431365
transform -1 0 25984 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0891__A3
timestamp 1698431365
transform 1 0 26208 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0892__I
timestamp 1698431365
transform 1 0 24304 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0893__A1
timestamp 1698431365
transform 1 0 26880 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0893__A3
timestamp 1698431365
transform 1 0 26320 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0896__A1
timestamp 1698431365
transform 1 0 18480 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0896__A2
timestamp 1698431365
transform 1 0 16800 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0897__A1
timestamp 1698431365
transform -1 0 18480 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0898__A1
timestamp 1698431365
transform -1 0 14112 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0898__A2
timestamp 1698431365
transform 1 0 14336 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0899__A1
timestamp 1698431365
transform 1 0 26544 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0899__A2
timestamp 1698431365
transform -1 0 21952 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0899__A3
timestamp 1698431365
transform -1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0900__B2
timestamp 1698431365
transform 1 0 15344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0901__A1
timestamp 1698431365
transform 1 0 16352 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0902__A2
timestamp 1698431365
transform 1 0 20272 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0902__A3
timestamp 1698431365
transform -1 0 20048 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0903__A2
timestamp 1698431365
transform 1 0 6944 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0903__B1
timestamp 1698431365
transform 1 0 6496 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0904__A1
timestamp 1698431365
transform 1 0 16576 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0904__A2
timestamp 1698431365
transform 1 0 19376 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0904__A3
timestamp 1698431365
transform 1 0 23408 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0905__A1
timestamp 1698431365
transform 1 0 14784 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0906__A2
timestamp 1698431365
transform 1 0 5824 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0906__B1
timestamp 1698431365
transform 1 0 6048 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0907__A1
timestamp 1698431365
transform 1 0 20384 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0907__A2
timestamp 1698431365
transform 1 0 15568 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0907__A3
timestamp 1698431365
transform 1 0 15120 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0908__A1
timestamp 1698431365
transform 1 0 20720 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0908__A2
timestamp 1698431365
transform 1 0 27552 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0909__A1
timestamp 1698431365
transform 1 0 15456 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0909__A2
timestamp 1698431365
transform 1 0 16352 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0909__A3
timestamp 1698431365
transform 1 0 15904 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0910__A2
timestamp 1698431365
transform 1 0 7056 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0910__B1
timestamp 1698431365
transform 1 0 7280 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0911__A1
timestamp 1698431365
transform 1 0 20720 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0911__A2
timestamp 1698431365
transform 1 0 24640 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0911__A3
timestamp 1698431365
transform 1 0 24192 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0912__A1
timestamp 1698431365
transform 1 0 16800 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0912__A2
timestamp 1698431365
transform 1 0 27888 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0912__A3
timestamp 1698431365
transform 1 0 27776 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0913__A2
timestamp 1698431365
transform 1 0 7168 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0913__B1
timestamp 1698431365
transform 1 0 6720 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0915__A1
timestamp 1698431365
transform 1 0 21840 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0915__A2
timestamp 1698431365
transform 1 0 21392 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0915__A3
timestamp 1698431365
transform 1 0 20608 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0916__A2
timestamp 1698431365
transform 1 0 14224 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0917__A1
timestamp 1698431365
transform 1 0 25312 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0917__A3
timestamp 1698431365
transform 1 0 27104 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0917__A4
timestamp 1698431365
transform 1 0 26208 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0919__A1
timestamp 1698431365
transform 1 0 23184 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0919__A2
timestamp 1698431365
transform 1 0 22736 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0919__A3
timestamp 1698431365
transform 1 0 22288 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0921__A1
timestamp 1698431365
transform 1 0 18592 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0921__A3
timestamp 1698431365
transform -1 0 17472 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0923__A1
timestamp 1698431365
transform 1 0 29232 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0923__A2
timestamp 1698431365
transform 1 0 26096 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0923__A3
timestamp 1698431365
transform 1 0 28224 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0924__A1
timestamp 1698431365
transform 1 0 17024 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0924__A2
timestamp 1698431365
transform 1 0 14448 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0924__A4
timestamp 1698431365
transform 1 0 16128 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0925__A2
timestamp 1698431365
transform 1 0 16688 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0927__A2
timestamp 1698431365
transform -1 0 23520 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0927__A3
timestamp 1698431365
transform -1 0 23968 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0928__A2
timestamp 1698431365
transform 1 0 20272 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0928__B
timestamp 1698431365
transform 1 0 18928 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0929__A1
timestamp 1698431365
transform -1 0 23072 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0930__A1
timestamp 1698431365
transform 1 0 29232 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0930__A2
timestamp 1698431365
transform 1 0 23296 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0930__A3
timestamp 1698431365
transform 1 0 24640 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0931__A2
timestamp 1698431365
transform 1 0 23408 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0931__B1
timestamp 1698431365
transform 1 0 25312 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0932__A1
timestamp 1698431365
transform -1 0 14896 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0933__A1
timestamp 1698431365
transform 1 0 20720 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0933__A2
timestamp 1698431365
transform -1 0 16576 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0933__A3
timestamp 1698431365
transform -1 0 17696 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0934__A2
timestamp 1698431365
transform 1 0 12656 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0934__B1
timestamp 1698431365
transform 1 0 14448 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0935__A1
timestamp 1698431365
transform 1 0 22736 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0935__A2
timestamp 1698431365
transform 1 0 23296 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0935__A3
timestamp 1698431365
transform 1 0 24640 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0936__A1
timestamp 1698431365
transform 1 0 19488 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0937__A2
timestamp 1698431365
transform 1 0 17920 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0937__B1
timestamp 1698431365
transform 1 0 17472 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0939__A3
timestamp 1698431365
transform -1 0 18368 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0939__A4
timestamp 1698431365
transform 1 0 17696 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0940__A1
timestamp 1698431365
transform 1 0 32816 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0940__A2
timestamp 1698431365
transform 1 0 28896 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0941__A2
timestamp 1698431365
transform -1 0 27888 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0942__A1
timestamp 1698431365
transform -1 0 28672 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0944__A2
timestamp 1698431365
transform 1 0 32368 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0944__B1
timestamp 1698431365
transform 1 0 32816 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0945__B1
timestamp 1698431365
transform -1 0 33488 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0946__A2
timestamp 1698431365
transform -1 0 33488 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0946__B1
timestamp 1698431365
transform 1 0 34720 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0947__A1
timestamp 1698431365
transform 1 0 30464 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0947__A3
timestamp 1698431365
transform 1 0 29792 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0948__A1
timestamp 1698431365
transform 1 0 30352 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0948__A3
timestamp 1698431365
transform 1 0 29904 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0952__A2
timestamp 1698431365
transform 1 0 7168 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0952__B1
timestamp 1698431365
transform 1 0 6720 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0953__A2
timestamp 1698431365
transform 1 0 6160 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0953__B1
timestamp 1698431365
transform 1 0 5712 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0954__A2
timestamp 1698431365
transform 1 0 6720 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0954__B1
timestamp 1698431365
transform 1 0 6272 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0955__A2
timestamp 1698431365
transform -1 0 5264 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0955__B1
timestamp 1698431365
transform 1 0 5488 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0956__A2
timestamp 1698431365
transform -1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0957__A2
timestamp 1698431365
transform 1 0 10752 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0958__A1
timestamp 1698431365
transform 1 0 24640 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0958__A3
timestamp 1698431365
transform -1 0 24864 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0958__A4
timestamp 1698431365
transform -1 0 23520 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0961__A1
timestamp 1698431365
transform 1 0 20160 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0961__A3
timestamp 1698431365
transform -1 0 19488 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0963__A1
timestamp 1698431365
transform -1 0 17024 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0963__A2
timestamp 1698431365
transform 1 0 15568 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0963__A4
timestamp 1698431365
transform -1 0 16576 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0964__A2
timestamp 1698431365
transform -1 0 16128 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0966__A2
timestamp 1698431365
transform -1 0 19488 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0966__B
timestamp 1698431365
transform -1 0 19936 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0967__A2
timestamp 1698431365
transform 1 0 24192 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0967__B1
timestamp 1698431365
transform 1 0 24640 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0968__A2
timestamp 1698431365
transform 1 0 11760 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0968__B1
timestamp 1698431365
transform 1 0 11312 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0969__A2
timestamp 1698431365
transform 1 0 17472 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0969__B1
timestamp 1698431365
transform 1 0 17024 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0971__A3
timestamp 1698431365
transform 1 0 18480 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0971__A4
timestamp 1698431365
transform 1 0 18704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0972__A2
timestamp 1698431365
transform 1 0 26992 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0973__A2
timestamp 1698431365
transform -1 0 28784 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0974__A1
timestamp 1698431365
transform 1 0 27440 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0976__A2
timestamp 1698431365
transform 1 0 33264 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0976__B1
timestamp 1698431365
transform 1 0 33712 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0977__B1
timestamp 1698431365
transform 1 0 35056 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0978__A2
timestamp 1698431365
transform -1 0 35168 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0978__B1
timestamp 1698431365
transform -1 0 34720 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0979__A1
timestamp 1698431365
transform 1 0 32368 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0979__A3
timestamp 1698431365
transform 1 0 31920 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0980__A1
timestamp 1698431365
transform 1 0 31472 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0980__A3
timestamp 1698431365
transform 1 0 31808 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0984__A2
timestamp 1698431365
transform 1 0 6608 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0984__B1
timestamp 1698431365
transform -1 0 7504 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0985__A2
timestamp 1698431365
transform -1 0 8176 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0985__B1
timestamp 1698431365
transform -1 0 7728 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0986__A2
timestamp 1698431365
transform 1 0 7280 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0986__B1
timestamp 1698431365
transform 1 0 6832 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0987__A2
timestamp 1698431365
transform 1 0 8064 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0987__B1
timestamp 1698431365
transform 1 0 7168 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0988__A2
timestamp 1698431365
transform 1 0 7728 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0989__A2
timestamp 1698431365
transform 1 0 11872 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0990__A1
timestamp 1698431365
transform 1 0 22288 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0990__A3
timestamp 1698431365
transform -1 0 24416 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0990__A4
timestamp 1698431365
transform 1 0 26880 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0993__A1
timestamp 1698431365
transform 1 0 21392 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0993__A3
timestamp 1698431365
transform -1 0 21616 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0995__A1
timestamp 1698431365
transform 1 0 17696 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0995__A2
timestamp 1698431365
transform 1 0 17696 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0995__A4
timestamp 1698431365
transform 1 0 16800 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0996__A2
timestamp 1698431365
transform 1 0 16576 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0998__A2
timestamp 1698431365
transform 1 0 19264 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0998__B
timestamp 1698431365
transform -1 0 19040 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0999__A2
timestamp 1698431365
transform 1 0 27888 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0999__B1
timestamp 1698431365
transform 1 0 27440 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1000__A2
timestamp 1698431365
transform 1 0 11984 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1000__B1
timestamp 1698431365
transform 1 0 11536 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1001__A2
timestamp 1698431365
transform -1 0 18256 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1001__B1
timestamp 1698431365
transform 1 0 18256 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1003__A3
timestamp 1698431365
transform 1 0 19600 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1003__A4
timestamp 1698431365
transform 1 0 19152 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1004__A2
timestamp 1698431365
transform 1 0 26656 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1005__A2
timestamp 1698431365
transform -1 0 28672 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1006__A1
timestamp 1698431365
transform 1 0 27664 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1008__A2
timestamp 1698431365
transform 1 0 34160 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1008__B1
timestamp 1698431365
transform 1 0 34048 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1009__B1
timestamp 1698431365
transform 1 0 35280 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1010__A2
timestamp 1698431365
transform -1 0 34944 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1010__B1
timestamp 1698431365
transform 1 0 36176 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1011__A1
timestamp 1698431365
transform 1 0 31584 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1011__A3
timestamp 1698431365
transform 1 0 31360 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1012__A1
timestamp 1698431365
transform -1 0 31808 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1012__A3
timestamp 1698431365
transform 1 0 32032 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1016__A2
timestamp 1698431365
transform 1 0 11088 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1016__B1
timestamp 1698431365
transform 1 0 10640 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1017__A2
timestamp 1698431365
transform 1 0 7616 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1017__B1
timestamp 1698431365
transform 1 0 7840 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1018__A2
timestamp 1698431365
transform 1 0 9184 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1018__B1
timestamp 1698431365
transform 1 0 10976 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1019__A2
timestamp 1698431365
transform 1 0 11312 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1019__B1
timestamp 1698431365
transform -1 0 11088 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1020__A2
timestamp 1698431365
transform 1 0 8512 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1021__A2
timestamp 1698431365
transform 1 0 9856 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1022__A1
timestamp 1698431365
transform 1 0 22736 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1022__A3
timestamp 1698431365
transform 1 0 24640 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1022__A4
timestamp 1698431365
transform 1 0 23184 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1025__A1
timestamp 1698431365
transform 1 0 21168 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1025__A3
timestamp 1698431365
transform 1 0 20720 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1027__A1
timestamp 1698431365
transform 1 0 18480 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1027__A2
timestamp 1698431365
transform 1 0 17248 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1027__A4
timestamp 1698431365
transform 1 0 16800 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1028__A2
timestamp 1698431365
transform 1 0 18144 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1029__A1
timestamp 1698431365
transform -1 0 18816 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1030__A2
timestamp 1698431365
transform 1 0 21504 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1030__B
timestamp 1698431365
transform 1 0 20720 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1031__A2
timestamp 1698431365
transform 1 0 26320 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1031__B1
timestamp 1698431365
transform 1 0 25872 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1032__A2
timestamp 1698431365
transform 1 0 12880 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1032__B1
timestamp 1698431365
transform 1 0 13776 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1032__B2
timestamp 1698431365
transform 1 0 13328 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1033__A2
timestamp 1698431365
transform 1 0 19712 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1033__B1
timestamp 1698431365
transform 1 0 18256 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1035__A3
timestamp 1698431365
transform 1 0 20832 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1035__A4
timestamp 1698431365
transform -1 0 19376 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1036__A2
timestamp 1698431365
transform 1 0 29232 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1037__A2
timestamp 1698431365
transform -1 0 27776 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1038__A1
timestamp 1698431365
transform 1 0 31584 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1040__A2
timestamp 1698431365
transform 1 0 19936 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1041__A2
timestamp 1698431365
transform 1 0 12320 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1042__A1
timestamp 1698431365
transform 1 0 30576 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1043__A1
timestamp 1698431365
transform 1 0 16352 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1043__A2
timestamp 1698431365
transform 1 0 25088 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1043__A3
timestamp 1698431365
transform 1 0 25760 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1043__A4
timestamp 1698431365
transform 1 0 17248 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1044__A1
timestamp 1698431365
transform -1 0 23520 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1044__A3
timestamp 1698431365
transform 1 0 23744 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1045__A3
timestamp 1698431365
transform -1 0 25760 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1046__A2
timestamp 1698431365
transform 1 0 17024 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1046__B1
timestamp 1698431365
transform 1 0 18480 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1047__A2
timestamp 1698431365
transform 1 0 25872 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1047__B1
timestamp 1698431365
transform 1 0 25424 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1050__A1
timestamp 1698431365
transform 1 0 31248 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1050__A2
timestamp 1698431365
transform 1 0 30128 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1050__A3
timestamp 1698431365
transform 1 0 30800 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1051__A1
timestamp 1698431365
transform 1 0 30128 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1051__A3
timestamp 1698431365
transform 1 0 30912 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1052__A2
timestamp 1698431365
transform 1 0 18928 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1052__B1
timestamp 1698431365
transform 1 0 21392 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1053__C
timestamp 1698431365
transform 1 0 30464 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1055__A1
timestamp 1698431365
transform 1 0 29232 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1055__A2
timestamp 1698431365
transform 1 0 29680 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1055__A3
timestamp 1698431365
transform -1 0 29120 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1056__A1
timestamp 1698431365
transform -1 0 24416 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1056__A3
timestamp 1698431365
transform -1 0 25984 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1057__A2
timestamp 1698431365
transform 1 0 12880 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1057__B1
timestamp 1698431365
transform 1 0 12432 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1061__A2
timestamp 1698431365
transform -1 0 13104 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1062__A2
timestamp 1698431365
transform -1 0 14448 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1062__B1
timestamp 1698431365
transform 1 0 15008 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1063__A2
timestamp 1698431365
transform 1 0 15904 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1064__A1
timestamp 1698431365
transform 1 0 28000 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1065__A1
timestamp 1698431365
transform 1 0 17696 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1065__A3
timestamp 1698431365
transform -1 0 20160 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1067__A1
timestamp 1698431365
transform 1 0 22848 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1067__A2
timestamp 1698431365
transform 1 0 19712 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1067__A4
timestamp 1698431365
transform 1 0 23408 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1068__A1
timestamp 1698431365
transform -1 0 17920 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1068__A3
timestamp 1698431365
transform 1 0 19824 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1069__A1
timestamp 1698431365
transform -1 0 23520 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1069__A2
timestamp 1698431365
transform -1 0 22512 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1070__A1
timestamp 1698431365
transform 1 0 25312 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1070__A2
timestamp 1698431365
transform 1 0 28224 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1071__A2
timestamp 1698431365
transform -1 0 10864 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1071__B1
timestamp 1698431365
transform -1 0 11200 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1073__A1
timestamp 1698431365
transform 1 0 28112 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1073__A2
timestamp 1698431365
transform 1 0 27664 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1073__A3
timestamp 1698431365
transform 1 0 27216 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1074__A1
timestamp 1698431365
transform 1 0 27552 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1075__A2
timestamp 1698431365
transform 1 0 8512 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1075__B1
timestamp 1698431365
transform -1 0 9184 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1076__A2
timestamp 1698431365
transform -1 0 17920 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1078__A2
timestamp 1698431365
transform 1 0 30464 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1078__B1
timestamp 1698431365
transform 1 0 30016 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1082__A2
timestamp 1698431365
transform 1 0 16800 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1082__B1
timestamp 1698431365
transform 1 0 16352 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1083__A2
timestamp 1698431365
transform 1 0 14896 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1083__B1
timestamp 1698431365
transform 1 0 16800 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1085__A1
timestamp 1698431365
transform -1 0 16464 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1085__A2
timestamp 1698431365
transform 1 0 17920 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1086__B1
timestamp 1698431365
transform -1 0 15456 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1087__A2
timestamp 1698431365
transform 1 0 12320 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1087__B1
timestamp 1698431365
transform 1 0 9632 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1090__A1
timestamp 1698431365
transform 1 0 24192 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1090__A3
timestamp 1698431365
transform -1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1091__A2
timestamp 1698431365
transform -1 0 14448 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1091__B1
timestamp 1698431365
transform -1 0 15008 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1092__A2
timestamp 1698431365
transform -1 0 14896 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1092__B
timestamp 1698431365
transform -1 0 15680 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1093__A2
timestamp 1698431365
transform 1 0 20384 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1094__A1
timestamp 1698431365
transform -1 0 27216 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1094__A2
timestamp 1698431365
transform 1 0 23744 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1094__A3
timestamp 1698431365
transform 1 0 26208 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1094__A4
timestamp 1698431365
transform -1 0 25984 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1095__B1
timestamp 1698431365
transform 1 0 17472 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1096__A1
timestamp 1698431365
transform -1 0 14448 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1097__A1
timestamp 1698431365
transform -1 0 16352 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1098__A1
timestamp 1698431365
transform 1 0 22176 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1098__A2
timestamp 1698431365
transform 1 0 23520 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1098__B1
timestamp 1698431365
transform 1 0 23072 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1099__A1
timestamp 1698431365
transform -1 0 20608 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1099__A2
timestamp 1698431365
transform 1 0 23408 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1101__A2
timestamp 1698431365
transform 1 0 20496 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1102__A2
timestamp 1698431365
transform 1 0 12208 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1102__B1
timestamp 1698431365
transform 1 0 12656 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1103__A1
timestamp 1698431365
transform 1 0 28448 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1103__A3
timestamp 1698431365
transform 1 0 22960 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1105__A1
timestamp 1698431365
transform 1 0 29680 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1105__A2
timestamp 1698431365
transform 1 0 28448 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1105__A3
timestamp 1698431365
transform 1 0 29232 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1106__A1
timestamp 1698431365
transform 1 0 24304 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1106__A2
timestamp 1698431365
transform 1 0 25312 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1106__B2
timestamp 1698431365
transform 1 0 25760 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1108__A1
timestamp 1698431365
transform 1 0 29680 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1108__A2
timestamp 1698431365
transform 1 0 27888 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1108__B1
timestamp 1698431365
transform 1 0 29008 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1108__B2
timestamp 1698431365
transform 1 0 28560 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1109__B1
timestamp 1698431365
transform 1 0 32816 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1112__A2
timestamp 1698431365
transform 1 0 28784 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1112__B
timestamp 1698431365
transform 1 0 32256 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1113__A1
timestamp 1698431365
transform -1 0 27440 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1114__A1
timestamp 1698431365
transform -1 0 17808 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1115__A3
timestamp 1698431365
transform 1 0 33152 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1116__A1
timestamp 1698431365
transform 1 0 34160 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1119__A1
timestamp 1698431365
transform 1 0 30576 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1119__A2
timestamp 1698431365
transform 1 0 30016 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1120__A1
timestamp 1698431365
transform -1 0 19824 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1120__A2
timestamp 1698431365
transform 1 0 20048 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1121__A1
timestamp 1698431365
transform -1 0 20720 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1121__A2
timestamp 1698431365
transform 1 0 19824 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1122__A1
timestamp 1698431365
transform 1 0 20048 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1122__A2
timestamp 1698431365
transform 1 0 19600 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1123__A1
timestamp 1698431365
transform -1 0 25200 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1123__A2
timestamp 1698431365
transform -1 0 24864 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1124__A1
timestamp 1698431365
transform -1 0 27104 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1124__A2
timestamp 1698431365
transform 1 0 22064 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1125__A1
timestamp 1698431365
transform -1 0 22288 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1125__A2
timestamp 1698431365
transform -1 0 22736 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1125__A3
timestamp 1698431365
transform -1 0 24304 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1132__A1
timestamp 1698431365
transform 1 0 30576 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1135__A1
timestamp 1698431365
transform 1 0 29792 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1137__A1
timestamp 1698431365
transform 1 0 30240 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1138__A1
timestamp 1698431365
transform 1 0 27328 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1140__A1
timestamp 1698431365
transform -1 0 31360 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1142__A1
timestamp 1698431365
transform 1 0 32368 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1144__A1
timestamp 1698431365
transform 1 0 35616 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1145__A2
timestamp 1698431365
transform -1 0 33376 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1146__A1
timestamp 1698431365
transform 1 0 33264 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1147__A1
timestamp 1698431365
transform 1 0 31920 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1150__A1
timestamp 1698431365
transform 1 0 29456 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1152__A1
timestamp 1698431365
transform 1 0 30464 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1153__A1
timestamp 1698431365
transform 1 0 29232 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1155__A1
timestamp 1698431365
transform 1 0 31360 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1157__A1
timestamp 1698431365
transform 1 0 28224 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1158__A2
timestamp 1698431365
transform 1 0 31584 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1159__A2
timestamp 1698431365
transform 1 0 33600 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1160__A1
timestamp 1698431365
transform 1 0 33152 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1162__A1
timestamp 1698431365
transform 1 0 30912 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1164__A1
timestamp 1698431365
transform 1 0 29232 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1165__A1
timestamp 1698431365
transform 1 0 30688 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1166__A1
timestamp 1698431365
transform 1 0 31024 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1168__A2
timestamp 1698431365
transform -1 0 23632 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1171__A1
timestamp 1698431365
transform 1 0 19152 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1171__A2
timestamp 1698431365
transform 1 0 18704 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1174__A1
timestamp 1698431365
transform 1 0 27888 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1175__A2
timestamp 1698431365
transform -1 0 29120 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1176__A2
timestamp 1698431365
transform 1 0 33712 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1177__A1
timestamp 1698431365
transform 1 0 32144 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1179__A1
timestamp 1698431365
transform 1 0 32368 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1180__A1
timestamp 1698431365
transform 1 0 31472 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1182__A1
timestamp 1698431365
transform 1 0 16800 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1183__A2
timestamp 1698431365
transform -1 0 21840 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1185__A3
timestamp 1698431365
transform 1 0 17584 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1187__I
timestamp 1698431365
transform 1 0 23520 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1188__A1
timestamp 1698431365
transform 1 0 27776 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1189__A2
timestamp 1698431365
transform 1 0 29232 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1190__A2
timestamp 1698431365
transform 1 0 32480 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1191__A1
timestamp 1698431365
transform 1 0 30576 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1192__I0
timestamp 1698431365
transform -1 0 33040 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1193__A1
timestamp 1698431365
transform -1 0 30352 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1195__A1
timestamp 1698431365
transform -1 0 24864 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1196__A2
timestamp 1698431365
transform 1 0 30352 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1199__A1
timestamp 1698431365
transform 1 0 28000 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1202__A1
timestamp 1698431365
transform 1 0 28000 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1203__A2
timestamp 1698431365
transform -1 0 28336 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1204__A2
timestamp 1698431365
transform 1 0 33040 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1205__A1
timestamp 1698431365
transform 1 0 32816 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1205__B1
timestamp 1698431365
transform 1 0 34048 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1207__A1
timestamp 1698431365
transform 1 0 29232 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1209__A1
timestamp 1698431365
transform 1 0 28448 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1210__A2
timestamp 1698431365
transform -1 0 28000 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1213__I
timestamp 1698431365
transform -1 0 27440 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1216__A3
timestamp 1698431365
transform 1 0 31136 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1217__A1
timestamp 1698431365
transform 1 0 29008 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1218__A1
timestamp 1698431365
transform 1 0 31024 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1220__A1
timestamp 1698431365
transform -1 0 30128 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1222__A1
timestamp 1698431365
transform 1 0 29232 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1225__A1
timestamp 1698431365
transform 1 0 26208 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1226__A1
timestamp 1698431365
transform 1 0 28448 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1226__A2
timestamp 1698431365
transform 1 0 29232 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1227__A1
timestamp 1698431365
transform 1 0 21392 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1228__I
timestamp 1698431365
transform 1 0 29680 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1230__A1
timestamp 1698431365
transform 1 0 27104 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1230__C
timestamp 1698431365
transform -1 0 32032 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1231__A2
timestamp 1698431365
transform 1 0 31696 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1235__A1
timestamp 1698431365
transform 1 0 28336 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1236__A2
timestamp 1698431365
transform 1 0 28000 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1237__A1
timestamp 1698431365
transform 1 0 30128 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1238__A1
timestamp 1698431365
transform 1 0 30912 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1238__A2
timestamp 1698431365
transform 1 0 30464 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1239__A1
timestamp 1698431365
transform 1 0 30352 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1239__B1
timestamp 1698431365
transform 1 0 29568 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1239__B2
timestamp 1698431365
transform -1 0 31024 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1240__A1
timestamp 1698431365
transform -1 0 25984 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1242__C
timestamp 1698431365
transform 1 0 31584 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1243__A1
timestamp 1698431365
transform 1 0 22960 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1243__A2
timestamp 1698431365
transform -1 0 26656 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1247__I
timestamp 1698431365
transform -1 0 6944 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1262__A1
timestamp 1698431365
transform 1 0 9744 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1262__A3
timestamp 1698431365
transform -1 0 14112 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1263__A2
timestamp 1698431365
transform 1 0 8960 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1263__B1
timestamp 1698431365
transform 1 0 10640 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1264__A1
timestamp 1698431365
transform 1 0 10640 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1265__A2
timestamp 1698431365
transform -1 0 4704 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1266__B
timestamp 1698431365
transform 1 0 18480 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1267__B
timestamp 1698431365
transform -1 0 5936 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1268__A2
timestamp 1698431365
transform 1 0 5600 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1269__B
timestamp 1698431365
transform 1 0 18592 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1270__B
timestamp 1698431365
transform 1 0 7168 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1271__A2
timestamp 1698431365
transform 1 0 7280 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1272__B
timestamp 1698431365
transform 1 0 23408 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1273__A2
timestamp 1698431365
transform -1 0 8848 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1273__B
timestamp 1698431365
transform 1 0 8400 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1274__A2
timestamp 1698431365
transform 1 0 6160 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1275__B
timestamp 1698431365
transform 1 0 19824 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1276__A2
timestamp 1698431365
transform 1 0 6832 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1276__B
timestamp 1698431365
transform 1 0 7280 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1277__A2
timestamp 1698431365
transform 1 0 9632 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1277__B1
timestamp 1698431365
transform 1 0 11088 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1278__A1
timestamp 1698431365
transform 1 0 8960 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1279__A2
timestamp 1698431365
transform 1 0 8288 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1279__B1
timestamp 1698431365
transform 1 0 10640 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1280__A1
timestamp 1698431365
transform 1 0 11088 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1281__A2
timestamp 1698431365
transform -1 0 9408 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1281__B1
timestamp 1698431365
transform 1 0 11088 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1282__A1
timestamp 1698431365
transform -1 0 8848 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1283__I
timestamp 1698431365
transform 1 0 5264 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1285__A2
timestamp 1698431365
transform 1 0 9296 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1286__A2
timestamp 1698431365
transform 1 0 12544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1288__A1
timestamp 1698431365
transform 1 0 35392 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1290__A1
timestamp 1698431365
transform 1 0 28448 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1290__A2
timestamp 1698431365
transform -1 0 26880 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1291__A2
timestamp 1698431365
transform -1 0 26432 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1292__A2
timestamp 1698431365
transform 1 0 27776 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1293__I
timestamp 1698431365
transform 1 0 10976 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1294__A2
timestamp 1698431365
transform 1 0 30016 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1295__A2
timestamp 1698431365
transform 1 0 27888 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1296__A2
timestamp 1698431365
transform 1 0 26992 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1299__A1
timestamp 1698431365
transform 1 0 12992 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1299__A2
timestamp 1698431365
transform 1 0 11648 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1301__A2
timestamp 1698431365
transform 1 0 12208 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1303__A2
timestamp 1698431365
transform 1 0 15232 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1305__I
timestamp 1698431365
transform 1 0 6944 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1306__A2
timestamp 1698431365
transform 1 0 19488 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1308__A2
timestamp 1698431365
transform -1 0 13328 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1310__A2
timestamp 1698431365
transform 1 0 9856 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1312__A2
timestamp 1698431365
transform 1 0 7504 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1314__A2
timestamp 1698431365
transform 1 0 7168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1316__A2
timestamp 1698431365
transform 1 0 8064 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1318__A1
timestamp 1698431365
transform -1 0 12544 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1318__A2
timestamp 1698431365
transform 1 0 10976 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1320__A2
timestamp 1698431365
transform 1 0 12768 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1322__A2
timestamp 1698431365
transform 1 0 7280 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1324__A2
timestamp 1698431365
transform 1 0 4592 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1326__A2
timestamp 1698431365
transform 1 0 5040 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1328__A2
timestamp 1698431365
transform 1 0 4816 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1330__A2
timestamp 1698431365
transform -1 0 6048 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1332__A2
timestamp 1698431365
transform 1 0 8960 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1334__A1
timestamp 1698431365
transform -1 0 11536 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1334__A2
timestamp 1698431365
transform 1 0 9968 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1336__A2
timestamp 1698431365
transform 1 0 10640 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1338__A2
timestamp 1698431365
transform 1 0 13552 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1340__A2
timestamp 1698431365
transform 1 0 14224 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1342__A2
timestamp 1698431365
transform 1 0 16576 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1344__A2
timestamp 1698431365
transform 1 0 20720 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1346__A1
timestamp 1698431365
transform 1 0 24192 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1346__A2
timestamp 1698431365
transform 1 0 22848 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1348__A2
timestamp 1698431365
transform 1 0 26880 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1350__A2
timestamp 1698431365
transform 1 0 30016 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1352__A2
timestamp 1698431365
transform 1 0 31248 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1354__A2
timestamp 1698431365
transform 1 0 26432 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1356__A2
timestamp 1698431365
transform 1 0 28336 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1358__A1
timestamp 1698431365
transform -1 0 25536 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1358__A2
timestamp 1698431365
transform 1 0 26320 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1360__A2
timestamp 1698431365
transform 1 0 15344 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1361__A2
timestamp 1698431365
transform 1 0 16800 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1362__A2
timestamp 1698431365
transform 1 0 22512 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1363__A2
timestamp 1698431365
transform 1 0 18928 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1364__A2
timestamp 1698431365
transform 1 0 18480 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1366__A2
timestamp 1698431365
transform 1 0 7280 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1368__A2
timestamp 1698431365
transform 1 0 4592 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1370__I
timestamp 1698431365
transform 1 0 5712 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1371__A2
timestamp 1698431365
transform 1 0 4144 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1373__A2
timestamp 1698431365
transform 1 0 5264 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1375__A2
timestamp 1698431365
transform 1 0 7504 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1377__A2
timestamp 1698431365
transform 1 0 8960 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1379__A2
timestamp 1698431365
transform 1 0 8624 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1381__A2
timestamp 1698431365
transform 1 0 4592 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1383__A2
timestamp 1698431365
transform 1 0 4592 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1385__A2
timestamp 1698431365
transform 1 0 5040 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1387__I
timestamp 1698431365
transform 1 0 34832 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1388__A2
timestamp 1698431365
transform 1 0 11312 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1390__A2
timestamp 1698431365
transform 1 0 15008 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1392__A2
timestamp 1698431365
transform -1 0 23408 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1394__A2
timestamp 1698431365
transform 1 0 30912 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1396__A2
timestamp 1698431365
transform -1 0 35504 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1398__A2
timestamp 1698431365
transform 1 0 35728 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1400__A2
timestamp 1698431365
transform 1 0 37072 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1402__A2
timestamp 1698431365
transform 1 0 32704 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1404__A2
timestamp 1698431365
transform 1 0 32256 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1406__A2
timestamp 1698431365
transform 1 0 33152 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1408__A2
timestamp 1698431365
transform 1 0 34944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1410__A2
timestamp 1698431365
transform 1 0 36064 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1412__A2
timestamp 1698431365
transform 1 0 35728 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1414__A2
timestamp 1698431365
transform 1 0 30576 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1415__A2
timestamp 1698431365
transform 1 0 30576 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1417__A2
timestamp 1698431365
transform 1 0 33152 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1419__A2
timestamp 1698431365
transform 1 0 37968 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1421__A2
timestamp 1698431365
transform 1 0 36400 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1423__A2
timestamp 1698431365
transform 1 0 35616 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1425__A2
timestamp 1698431365
transform 1 0 27440 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1427__A2
timestamp 1698431365
transform 1 0 27664 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1429__A2
timestamp 1698431365
transform 1 0 31136 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1431__A2
timestamp 1698431365
transform 1 0 34048 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1433__A2
timestamp 1698431365
transform 1 0 36288 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1435__A2
timestamp 1698431365
transform 1 0 36624 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1437__A1
timestamp 1698431365
transform -1 0 12992 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1437__A2
timestamp 1698431365
transform 1 0 11424 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1439__A2
timestamp 1698431365
transform 1 0 12208 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1441__A2
timestamp 1698431365
transform 1 0 7504 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1443__A2
timestamp 1698431365
transform 1 0 9184 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1445__A2
timestamp 1698431365
transform 1 0 10528 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1447__A2
timestamp 1698431365
transform 1 0 6608 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1449__A2
timestamp 1698431365
transform 1 0 9968 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1451__A2
timestamp 1698431365
transform -1 0 9968 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1453__A2
timestamp 1698431365
transform 1 0 15232 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1454__A2
timestamp 1698431365
transform 1 0 17808 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1455__A2
timestamp 1698431365
transform 1 0 20720 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1456__A2
timestamp 1698431365
transform 1 0 20272 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1457__A1
timestamp 1698431365
transform 1 0 27440 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1457__A2
timestamp 1698431365
transform 1 0 28336 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1459__A2
timestamp 1698431365
transform 1 0 16800 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1461__I
timestamp 1698431365
transform 1 0 30240 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1462__A2
timestamp 1698431365
transform 1 0 13888 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1464__A2
timestamp 1698431365
transform 1 0 15792 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1466__A2
timestamp 1698431365
transform -1 0 17696 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1468__I
timestamp 1698431365
transform 1 0 7392 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1469__A2
timestamp 1698431365
transform 1 0 20944 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1471__A2
timestamp 1698431365
transform 1 0 23184 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1473__A1
timestamp 1698431365
transform 1 0 24528 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1473__A2
timestamp 1698431365
transform 1 0 23184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1475__A2
timestamp 1698431365
transform 1 0 25200 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1477__A2
timestamp 1698431365
transform 1 0 25088 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1479__A2
timestamp 1698431365
transform 1 0 31920 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1481__A2
timestamp 1698431365
transform 1 0 32144 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1483__A2
timestamp 1698431365
transform 1 0 26880 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1485__A1
timestamp 1698431365
transform 1 0 21504 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1485__A2
timestamp 1698431365
transform 1 0 19936 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1487__A2
timestamp 1698431365
transform 1 0 5040 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1489__A2
timestamp 1698431365
transform 1 0 4368 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1491__A2
timestamp 1698431365
transform 1 0 6944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1493__A2
timestamp 1698431365
transform 1 0 10528 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1495__A2
timestamp 1698431365
transform -1 0 12432 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1497__A2
timestamp 1698431365
transform 1 0 12880 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1499__A2
timestamp 1698431365
transform -1 0 13104 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1500__A2
timestamp 1698431365
transform 1 0 12432 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1501__A2
timestamp 1698431365
transform 1 0 15120 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1502__A2
timestamp 1698431365
transform 1 0 14112 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1503__A2
timestamp 1698431365
transform 1 0 12432 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1504__A2
timestamp 1698431365
transform 1 0 13776 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1505__A2
timestamp 1698431365
transform 1 0 15120 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1507__A2
timestamp 1698431365
transform 1 0 15008 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1509__A2
timestamp 1698431365
transform 1 0 15904 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1511__A2
timestamp 1698431365
transform 1 0 18592 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1513__A2
timestamp 1698431365
transform 1 0 15456 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1515__A2
timestamp 1698431365
transform 1 0 10528 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1517__A2
timestamp 1698431365
transform 1 0 6608 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1519__A2
timestamp 1698431365
transform 1 0 5040 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1521__A2
timestamp 1698431365
transform 1 0 7392 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1523__A2
timestamp 1698431365
transform 1 0 10528 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1525__A2
timestamp 1698431365
transform 1 0 12656 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1527__A2
timestamp 1698431365
transform 1 0 19040 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1529__A2
timestamp 1698431365
transform 1 0 27776 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1531__A2
timestamp 1698431365
transform 1 0 31024 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1533__A2
timestamp 1698431365
transform 1 0 31472 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1535__A2
timestamp 1698431365
transform 1 0 29232 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1537__A2
timestamp 1698431365
transform 1 0 25200 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1539__A2
timestamp 1698431365
transform 1 0 26656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1541__A2
timestamp 1698431365
transform 1 0 31360 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1543__A2
timestamp 1698431365
transform 1 0 34608 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1545__A2
timestamp 1698431365
transform 1 0 34272 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1547__A2
timestamp 1698431365
transform 1 0 32704 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1549__A2
timestamp 1698431365
transform 1 0 21504 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1551__A1
timestamp 1698431365
transform -1 0 21616 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1551__A2
timestamp 1698431365
transform 1 0 21056 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1553__A2
timestamp 1698431365
transform 1 0 19712 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1555__A2
timestamp 1698431365
transform 1 0 19712 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1557__A2
timestamp 1698431365
transform -1 0 23184 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1559__I
timestamp 1698431365
transform 1 0 21840 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1560__A2
timestamp 1698431365
transform 1 0 22848 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1562__A2
timestamp 1698431365
transform 1 0 23072 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1564__A2
timestamp 1698431365
transform 1 0 22848 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1566__A2
timestamp 1698431365
transform 1 0 23520 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1568__A2
timestamp 1698431365
transform 1 0 24864 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1570__A2
timestamp 1698431365
transform 1 0 28000 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1572__A2
timestamp 1698431365
transform 1 0 27104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1574__A2
timestamp 1698431365
transform 1 0 26432 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1576__A1
timestamp 1698431365
transform -1 0 28784 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1576__A2
timestamp 1698431365
transform 1 0 28784 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1578__A2
timestamp 1698431365
transform 1 0 30576 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1580__A2
timestamp 1698431365
transform 1 0 34608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1582__A2
timestamp 1698431365
transform 1 0 34944 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1584__A2
timestamp 1698431365
transform 1 0 35168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1586__A1
timestamp 1698431365
transform 1 0 24080 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1586__A2
timestamp 1698431365
transform 1 0 22960 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1588__A1
timestamp 1698431365
transform -1 0 23520 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1588__A2
timestamp 1698431365
transform 1 0 22848 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1590__A2
timestamp 1698431365
transform -1 0 23968 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1592__A2
timestamp 1698431365
transform 1 0 26656 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1594__A2
timestamp 1698431365
transform 1 0 26208 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1596__A2
timestamp 1698431365
transform 1 0 23744 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1598__A2
timestamp 1698431365
transform 1 0 23856 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1599__A2
timestamp 1698431365
transform 1 0 23408 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1602__A2
timestamp 1698431365
transform 1 0 4480 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1604__A2
timestamp 1698431365
transform 1 0 4816 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1606__A2
timestamp 1698431365
transform 1 0 5040 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1608__A2
timestamp 1698431365
transform 1 0 8064 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1610__A2
timestamp 1698431365
transform 1 0 12320 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1612__A2
timestamp 1698431365
transform 1 0 11088 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1614__A2
timestamp 1698431365
transform 1 0 8960 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1616__A2
timestamp 1698431365
transform 1 0 8960 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1618__A2
timestamp 1698431365
transform 1 0 10080 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1620__A2
timestamp 1698431365
transform 1 0 11424 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1622__A2
timestamp 1698431365
transform 1 0 12880 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1624__A2
timestamp 1698431365
transform 1 0 14896 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1626__A2
timestamp 1698431365
transform 1 0 13664 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1628__A2
timestamp 1698431365
transform 1 0 15008 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1630__A2
timestamp 1698431365
transform 1 0 16800 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1632__A2
timestamp 1698431365
transform 1 0 16800 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1634__A2
timestamp 1698431365
transform 1 0 17584 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1636__A2
timestamp 1698431365
transform 1 0 5040 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1638__A2
timestamp 1698431365
transform 1 0 4592 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1640__A2
timestamp 1698431365
transform -1 0 4816 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1642__A2
timestamp 1698431365
transform 1 0 7616 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1644__A2
timestamp 1698431365
transform 1 0 7616 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1646__A2
timestamp 1698431365
transform 1 0 8176 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1648__A2
timestamp 1698431365
transform 1 0 5712 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1650__A2
timestamp 1698431365
transform 1 0 4928 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1652__A2
timestamp 1698431365
transform 1 0 5488 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1654__A2
timestamp 1698431365
transform 1 0 8064 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1656__A2
timestamp 1698431365
transform 1 0 8960 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1658__A2
timestamp 1698431365
transform 1 0 17024 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1660__A2
timestamp 1698431365
transform 1 0 18032 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1663__A1
timestamp 1698431365
transform 1 0 15904 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1663__B
timestamp 1698431365
transform 1 0 15904 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1664__A1
timestamp 1698431365
transform 1 0 15792 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1665__A1
timestamp 1698431365
transform 1 0 15008 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1665__B
timestamp 1698431365
transform -1 0 14448 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1666__A1
timestamp 1698431365
transform 1 0 15344 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1667__A1
timestamp 1698431365
transform 1 0 15008 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1667__B
timestamp 1698431365
transform 1 0 12880 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1668__A1
timestamp 1698431365
transform -1 0 12208 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1669__A1
timestamp 1698431365
transform 1 0 18368 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1669__B
timestamp 1698431365
transform 1 0 18816 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1670__A1
timestamp 1698431365
transform 1 0 15456 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1671__A1
timestamp 1698431365
transform 1 0 21392 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1671__B
timestamp 1698431365
transform 1 0 19488 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1672__A1
timestamp 1698431365
transform -1 0 17808 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1673__B
timestamp 1698431365
transform 1 0 22176 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1674__A1
timestamp 1698431365
transform 1 0 24304 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1675__A2
timestamp 1698431365
transform 1 0 18144 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1676__A1
timestamp 1698431365
transform 1 0 17584 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1677__A1
timestamp 1698431365
transform 1 0 20272 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1677__A2
timestamp 1698431365
transform 1 0 19936 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1678__A1
timestamp 1698431365
transform 1 0 17136 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1678__B
timestamp 1698431365
transform 1 0 17584 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1679__A1
timestamp 1698431365
transform 1 0 14000 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1679__A2
timestamp 1698431365
transform 1 0 14448 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1680__A1
timestamp 1698431365
transform 1 0 11536 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1682__A1
timestamp 1698431365
transform -1 0 13104 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1682__A2
timestamp 1698431365
transform 1 0 15232 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1682__B
timestamp 1698431365
transform 1 0 14784 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1683__B
timestamp 1698431365
transform 1 0 13664 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1684__A1
timestamp 1698431365
transform 1 0 13776 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1685__B
timestamp 1698431365
transform 1 0 12880 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1686__A1
timestamp 1698431365
transform 1 0 16016 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1687__A1
timestamp 1698431365
transform 1 0 13776 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1688__A1
timestamp 1698431365
transform 1 0 15232 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1689__A1
timestamp 1698431365
transform 1 0 18256 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1690__A1
timestamp 1698431365
transform 1 0 15904 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1691__A1
timestamp 1698431365
transform -1 0 27552 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1692__A1
timestamp 1698431365
transform 1 0 24080 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1694__A1
timestamp 1698431365
transform 1 0 29680 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1696__B
timestamp 1698431365
transform 1 0 31248 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1698__B
timestamp 1698431365
transform 1 0 32032 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1699__A1
timestamp 1698431365
transform 1 0 37296 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1700__A1
timestamp 1698431365
transform 1 0 35056 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1701__A1
timestamp 1698431365
transform 1 0 36848 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1703__A1
timestamp 1698431365
transform 1 0 38080 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1705__B
timestamp 1698431365
transform -1 0 34160 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1706__A1
timestamp 1698431365
transform 1 0 33936 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1707__A1
timestamp 1698431365
transform 1 0 36176 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1708__CLK
timestamp 1698431365
transform 1 0 11536 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1709__CLK
timestamp 1698431365
transform 1 0 7056 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1710__CLK
timestamp 1698431365
transform 1 0 6944 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1711__CLK
timestamp 1698431365
transform 1 0 7728 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1712__CLK
timestamp 1698431365
transform 1 0 5264 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1713__CLK
timestamp 1698431365
transform 1 0 10640 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1714__CLK
timestamp 1698431365
transform 1 0 10976 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1715__CLK
timestamp 1698431365
transform -1 0 9856 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1716__CLK
timestamp 1698431365
transform 1 0 8960 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1717__CLK
timestamp 1698431365
transform 1 0 38192 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1718__CLK
timestamp 1698431365
transform 1 0 29232 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1719__CLK
timestamp 1698431365
transform 1 0 30128 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1720__CLK
timestamp 1698431365
transform 1 0 30576 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1721__CLK
timestamp 1698431365
transform 1 0 32256 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1722__CLK
timestamp 1698431365
transform 1 0 30912 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1723__CLK
timestamp 1698431365
transform 1 0 28560 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1724__CLK
timestamp 1698431365
transform 1 0 13552 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1725__CLK
timestamp 1698431365
transform 1 0 15120 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1726__CLK
timestamp 1698431365
transform 1 0 19040 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1727__CLK
timestamp 1698431365
transform 1 0 21728 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1728__CLK
timestamp 1698431365
transform 1 0 14672 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1729__CLK
timestamp 1698431365
transform 1 0 11312 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1730__CLK
timestamp 1698431365
transform 1 0 7952 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1731__CLK
timestamp 1698431365
transform 1 0 8960 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1732__CLK
timestamp 1698431365
transform 1 0 12432 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1733__CLK
timestamp 1698431365
transform 1 0 13552 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1734__CLK
timestamp 1698431365
transform 1 0 11648 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1735__CLK
timestamp 1698431365
transform 1 0 5040 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1736__CLK
timestamp 1698431365
transform 1 0 5040 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1737__CLK
timestamp 1698431365
transform 1 0 5040 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1738__CLK
timestamp 1698431365
transform 1 0 6160 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1739__CLK
timestamp 1698431365
transform 1 0 9632 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1740__CLK
timestamp 1698431365
transform 1 0 11648 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1741__CLK
timestamp 1698431365
transform 1 0 12320 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1742__CLK
timestamp 1698431365
transform 1 0 14000 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1743__CLK
timestamp 1698431365
transform 1 0 16240 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1744__CLK
timestamp 1698431365
transform 1 0 16352 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1745__CLK
timestamp 1698431365
transform 1 0 16800 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1746__CLK
timestamp 1698431365
transform 1 0 24640 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1747__CLK
timestamp 1698431365
transform 1 0 29232 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1748__CLK
timestamp 1698431365
transform 1 0 30688 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1749__CLK
timestamp 1698431365
transform 1 0 32816 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1750__CLK
timestamp 1698431365
transform 1 0 33824 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1751__CLK
timestamp 1698431365
transform 1 0 31808 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1752__CLK
timestamp 1698431365
transform 1 0 27216 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1753__CLK
timestamp 1698431365
transform 1 0 27776 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1754__CLK
timestamp 1698431365
transform 1 0 14448 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1755__CLK
timestamp 1698431365
transform 1 0 15792 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1756__CLK
timestamp 1698431365
transform 1 0 16800 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1757__CLK
timestamp 1698431365
transform 1 0 16800 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1758__CLK
timestamp 1698431365
transform 1 0 15792 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1759__CLK
timestamp 1698431365
transform 1 0 4816 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1760__CLK
timestamp 1698431365
transform 1 0 5040 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1761__CLK
timestamp 1698431365
transform 1 0 5040 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1762__CLK
timestamp 1698431365
transform 1 0 7168 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1763__CLK
timestamp 1698431365
transform -1 0 9856 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1764__CLK
timestamp 1698431365
transform -1 0 9408 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1765__CLK
timestamp 1698431365
transform 1 0 5040 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1766__CLK
timestamp 1698431365
transform 1 0 5040 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1767__CLK
timestamp 1698431365
transform 1 0 5488 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1768__CLK
timestamp 1698431365
transform 1 0 10080 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1769__CLK
timestamp 1698431365
transform 1 0 13552 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1770__CLK
timestamp 1698431365
transform 1 0 17248 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1771__CLK
timestamp 1698431365
transform 1 0 28560 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1772__CLK
timestamp 1698431365
transform 1 0 36400 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1773__CLK
timestamp 1698431365
transform 1 0 38192 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1774__CLK
timestamp 1698431365
transform 1 0 38192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1775__CLK
timestamp 1698431365
transform 1 0 38192 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1776__CLK
timestamp 1698431365
transform 1 0 33152 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1777__CLK
timestamp 1698431365
transform 1 0 33712 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1778__CLK
timestamp 1698431365
transform 1 0 35504 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1779__CLK
timestamp 1698431365
transform 1 0 38192 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1780__CLK
timestamp 1698431365
transform 1 0 38192 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1781__CLK
timestamp 1698431365
transform 1 0 36400 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1782__CLK
timestamp 1698431365
transform 1 0 31024 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1783__CLK
timestamp 1698431365
transform 1 0 30800 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1784__CLK
timestamp 1698431365
transform 1 0 34944 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1785__CLK
timestamp 1698431365
transform 1 0 38192 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1786__CLK
timestamp 1698431365
transform 1 0 38192 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1787__CLK
timestamp 1698431365
transform 1 0 35168 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1788__CLK
timestamp 1698431365
transform 1 0 29680 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1789__CLK
timestamp 1698431365
transform 1 0 30240 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1790__CLK
timestamp 1698431365
transform 1 0 33824 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1791__CLK
timestamp 1698431365
transform 1 0 34944 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1792__CLK
timestamp 1698431365
transform 1 0 38192 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1793__CLK
timestamp 1698431365
transform 1 0 38192 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1794__CLK
timestamp 1698431365
transform 1 0 14224 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1795__CLK
timestamp 1698431365
transform 1 0 12432 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1796__CLK
timestamp 1698431365
transform 1 0 8848 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1797__CLK
timestamp 1698431365
transform 1 0 9520 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1798__CLK
timestamp 1698431365
transform 1 0 7056 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1799__CLK
timestamp 1698431365
transform 1 0 8736 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1800__CLK
timestamp 1698431365
transform -1 0 10080 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1801__CLK
timestamp 1698431365
transform -1 0 14560 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1802__CLK
timestamp 1698431365
transform 1 0 18816 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1803__CLK
timestamp 1698431365
transform -1 0 22400 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1804__CLK
timestamp 1698431365
transform 1 0 23072 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1805__CLK
timestamp 1698431365
transform 1 0 24640 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1806__CLK
timestamp 1698431365
transform -1 0 22848 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1807__CLK
timestamp 1698431365
transform -1 0 16688 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1808__CLK
timestamp 1698431365
transform 1 0 15120 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1809__CLK
timestamp 1698431365
transform 1 0 17472 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1810__CLK
timestamp 1698431365
transform 1 0 16800 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1811__CLK
timestamp 1698431365
transform 1 0 24640 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1812__CLK
timestamp 1698431365
transform 1 0 24640 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1813__CLK
timestamp 1698431365
transform 1 0 26656 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1814__CLK
timestamp 1698431365
transform 1 0 28336 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1815__CLK
timestamp 1698431365
transform 1 0 30352 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1816__CLK
timestamp 1698431365
transform 1 0 32480 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1817__CLK
timestamp 1698431365
transform 1 0 29904 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1818__CLK
timestamp 1698431365
transform 1 0 27104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1819__CLK
timestamp 1698431365
transform 1 0 11424 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1820__CLK
timestamp 1698431365
transform 1 0 6720 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1821__CLK
timestamp 1698431365
transform 1 0 4816 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1822__CLK
timestamp 1698431365
transform 1 0 9856 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1823__CLK
timestamp 1698431365
transform 1 0 12992 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1824__CLK
timestamp 1698431365
transform 1 0 14448 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1825__CLK
timestamp 1698431365
transform 1 0 13552 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1826__CLK
timestamp 1698431365
transform 1 0 14672 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1827__CLK
timestamp 1698431365
transform 1 0 14784 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1828__CLK
timestamp 1698431365
transform 1 0 16800 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1829__CLK
timestamp 1698431365
transform 1 0 15568 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1830__CLK
timestamp 1698431365
transform 1 0 14672 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1831__CLK
timestamp 1698431365
transform 1 0 16800 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1831__D
timestamp 1698431365
transform 1 0 17248 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1832__CLK
timestamp 1698431365
transform 1 0 15456 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1833__CLK
timestamp 1698431365
transform 1 0 16800 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1834__CLK
timestamp 1698431365
transform 1 0 18928 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1835__CLK
timestamp 1698431365
transform 1 0 19040 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1836__CLK
timestamp 1698431365
transform 1 0 16800 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1837__CLK
timestamp 1698431365
transform 1 0 9632 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1838__CLK
timestamp 1698431365
transform 1 0 5040 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1839__CLK
timestamp 1698431365
transform -1 0 6048 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1840__CLK
timestamp 1698431365
transform -1 0 9632 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1841__CLK
timestamp 1698431365
transform 1 0 14000 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1842__CLK
timestamp 1698431365
transform 1 0 16688 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1843__CLK
timestamp 1698431365
transform 1 0 24640 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1844__CLK
timestamp 1698431365
transform 1 0 30128 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1845__CLK
timestamp 1698431365
transform 1 0 33600 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1846__CLK
timestamp 1698431365
transform 1 0 33152 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1847__CLK
timestamp 1698431365
transform 1 0 28560 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1848__CLK
timestamp 1698431365
transform -1 0 27776 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1849__CLK
timestamp 1698431365
transform 1 0 32480 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1850__CLK
timestamp 1698431365
transform 1 0 30016 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1851__CLK
timestamp 1698431365
transform 1 0 32480 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1852__CLK
timestamp 1698431365
transform 1 0 34944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1853__CLK
timestamp 1698431365
transform 1 0 32704 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1854__CLK
timestamp 1698431365
transform 1 0 23856 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1855__CLK
timestamp 1698431365
transform 1 0 20944 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1856__CLK
timestamp 1698431365
transform 1 0 22400 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1857__CLK
timestamp 1698431365
transform 1 0 22288 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1858__CLK
timestamp 1698431365
transform 1 0 23296 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1859__CLK
timestamp 1698431365
transform 1 0 24192 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1860__CLK
timestamp 1698431365
transform 1 0 23072 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1861__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1862__CLK
timestamp 1698431365
transform -1 0 26656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1863__CLK
timestamp 1698431365
transform 1 0 27440 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1864__CLK
timestamp 1698431365
transform 1 0 28672 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1865__CLK
timestamp 1698431365
transform 1 0 30128 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1866__CLK
timestamp 1698431365
transform 1 0 29232 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1867__CLK
timestamp 1698431365
transform 1 0 32256 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1868__CLK
timestamp 1698431365
transform 1 0 31472 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1869__CLK
timestamp 1698431365
transform 1 0 35056 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1870__CLK
timestamp 1698431365
transform 1 0 34496 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1871__CLK
timestamp 1698431365
transform 1 0 34608 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1872__CLK
timestamp 1698431365
transform 1 0 25536 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1873__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1874__CLK
timestamp 1698431365
transform 1 0 25984 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1875__CLK
timestamp 1698431365
transform 1 0 27440 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1876__CLK
timestamp 1698431365
transform 1 0 27776 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1877__CLK
timestamp 1698431365
transform 1 0 28448 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1878__CLK
timestamp 1698431365
transform 1 0 26880 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1879__CLK
timestamp 1698431365
transform 1 0 9184 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1880__CLK
timestamp 1698431365
transform 1 0 4368 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1881__CLK
timestamp 1698431365
transform 1 0 5488 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1882__CLK
timestamp 1698431365
transform 1 0 8624 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1883__CLK
timestamp 1698431365
transform 1 0 12768 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1884__CLK
timestamp 1698431365
transform 1 0 14112 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1885__CLK
timestamp 1698431365
transform 1 0 11648 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1886__CLK
timestamp 1698431365
transform 1 0 10864 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1887__CLK
timestamp 1698431365
transform 1 0 10640 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1888__CLK
timestamp 1698431365
transform -1 0 12880 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1889__CLK
timestamp 1698431365
transform 1 0 14448 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1890__CLK
timestamp 1698431365
transform 1 0 14896 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1891__CLK
timestamp 1698431365
transform 1 0 16464 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1892__CLK
timestamp 1698431365
transform 1 0 16240 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1893__CLK
timestamp 1698431365
transform 1 0 18256 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1894__CLK
timestamp 1698431365
transform -1 0 19152 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1895__CLK
timestamp 1698431365
transform 1 0 20496 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1896__CLK
timestamp 1698431365
transform 1 0 20384 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1897__CLK
timestamp 1698431365
transform 1 0 5712 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1898__CLK
timestamp 1698431365
transform 1 0 4816 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1899__CLK
timestamp 1698431365
transform 1 0 5712 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1900__CLK
timestamp 1698431365
transform 1 0 9632 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1901__CLK
timestamp 1698431365
transform 1 0 9632 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1902__CLK
timestamp 1698431365
transform 1 0 9408 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1903__CLK
timestamp 1698431365
transform 1 0 5264 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1904__CLK
timestamp 1698431365
transform 1 0 5712 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1905__CLK
timestamp 1698431365
transform 1 0 7392 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1906__CLK
timestamp 1698431365
transform 1 0 10528 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1907__CLK
timestamp 1698431365
transform 1 0 13552 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1908__CLK
timestamp 1698431365
transform 1 0 20272 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1909__CLK
timestamp 1698431365
transform 1 0 16800 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1910__CLK
timestamp 1698431365
transform 1 0 16352 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1911__CLK
timestamp 1698431365
transform 1 0 14560 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1912__CLK
timestamp 1698431365
transform 1 0 17472 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1913__CLK
timestamp 1698431365
transform 1 0 20720 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1914__CLK
timestamp 1698431365
transform -1 0 25088 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1915__CLK
timestamp 1698431365
transform 1 0 16352 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1916__CLK
timestamp 1698431365
transform -1 0 17360 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1917__CLK
timestamp 1698431365
transform 1 0 17024 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1918__CLK
timestamp 1698431365
transform 1 0 14112 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1919__CLK
timestamp 1698431365
transform 1 0 15456 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1920__CLK
timestamp 1698431365
transform 1 0 15904 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1921__CLK
timestamp 1698431365
transform -1 0 16576 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1922__CLK
timestamp 1698431365
transform 1 0 19488 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1923__CLK
timestamp 1698431365
transform -1 0 31136 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1924__CLK
timestamp 1698431365
transform 1 0 32480 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1925__CLK
timestamp 1698431365
transform 1 0 32480 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1926__CLK
timestamp 1698431365
transform 1 0 32480 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1927__CLK
timestamp 1698431365
transform 1 0 34496 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1928__CLK
timestamp 1698431365
transform 1 0 33824 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1929__CLK
timestamp 1698431365
transform 1 0 34608 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698431365
transform 1 0 20272 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_0__f_clk_I
timestamp 1698431365
transform 1 0 15456 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_1__f_clk_I
timestamp 1698431365
transform 1 0 20384 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_2__f_clk_I
timestamp 1698431365
transform 1 0 31248 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_3__f_clk_I
timestamp 1698431365
transform 1 0 25312 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_dec1._061__I
timestamp 1698431365
transform 1 0 33600 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_dec1._062__A1
timestamp 1698431365
transform 1 0 37184 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_dec1._101__A1
timestamp 1698431365
transform 1 0 36064 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_dec1._114__A1
timestamp 1698431365
transform 1 0 38192 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_dec1._118__A1
timestamp 1698431365
transform 1 0 36736 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_dec1._122__A1
timestamp 1698431365
transform 1 0 37632 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_dec1._123__B2
timestamp 1698431365
transform 1 0 34048 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout43_I
timestamp 1698431365
transform 1 0 17472 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout44_I
timestamp 1698431365
transform 1 0 20048 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout45_I
timestamp 1698431365
transform 1 0 18256 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout46_I
timestamp 1698431365
transform -1 0 31472 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout47_I
timestamp 1698431365
transform -1 0 35056 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout48_I
timestamp 1698431365
transform 1 0 30800 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout49_I
timestamp 1698431365
transform 1 0 13216 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout50_I
timestamp 1698431365
transform 1 0 15568 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout51_I
timestamp 1698431365
transform 1 0 16576 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout52_I
timestamp 1698431365
transform 1 0 37744 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout53_I
timestamp 1698431365
transform 1 0 37744 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform 1 0 37408 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform 1 0 27776 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform 1 0 27328 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform 1 0 26432 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform -1 0 24864 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform -1 0 24416 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform -1 0 22736 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform 1 0 23632 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform -1 0 20944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform -1 0 19600 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform -1 0 19152 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform 1 0 36512 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698431365
transform -1 0 17360 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698431365
transform 1 0 18368 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698431365
transform 1 0 18144 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698431365
transform 1 0 15456 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698431365
transform 1 0 15008 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1698431365
transform -1 0 13776 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1698431365
transform -1 0 12544 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1698431365
transform 1 0 12096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1698431365
transform 1 0 11424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1698431365
transform -1 0 9856 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1698431365
transform 1 0 36064 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1698431365
transform -1 0 9184 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1698431365
transform 1 0 8512 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1698431365
transform 1 0 35280 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1698431365
transform -1 0 32704 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1698431365
transform -1 0 32032 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1698431365
transform -1 0 30800 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1698431365
transform -1 0 29904 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1698431365
transform -1 0 29008 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1698431365
transform -1 0 28448 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1698431365
transform 1 0 7616 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input34_I
timestamp 1698431365
transform -1 0 5152 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input35_I
timestamp 1698431365
transform -1 0 3920 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input36_I
timestamp 1698431365
transform -1 0 38416 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input37_I
timestamp 1698431365
transform -1 0 38416 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input38_I
timestamp 1698431365
transform -1 0 38416 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input39_I
timestamp 1698431365
transform -1 0 38416 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input40_I
timestamp 1698431365
transform -1 0 38416 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input41_I
timestamp 1698431365
transform -1 0 37744 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input42_I
timestamp 1698431365
transform -1 0 3472 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac._4__I
timestamp 1698431365
transform 1 0 15120 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac._5__A2
timestamp 1698431365
transform 1 0 14224 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[0\].vdac_batch._4__A2
timestamp 1698431365
transform -1 0 24192 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[0\].vdac_batch._5__A1
timestamp 1698431365
transform 1 0 25088 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[0\].vdac_batch._7__I
timestamp 1698431365
transform 1 0 26096 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].vref_I
timestamp 1698431365
transform 1 0 24640 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[1\].vdac_batch._4__A2
timestamp 1698431365
transform 1 0 22288 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[1\].vdac_batch._5__A1
timestamp 1698431365
transform 1 0 20720 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[1\].vdac_batch._7__I
timestamp 1698431365
transform 1 0 23184 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[0\].vref_I
timestamp 1698431365
transform 1 0 20720 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].vref_I
timestamp 1698431365
transform 1 0 20048 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[2\].vdac_batch._4__A2
timestamp 1698431365
transform 1 0 18592 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[2\].vdac_batch._5__A1
timestamp 1698431365
transform 1 0 17248 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[2\].vdac_batch._7__I
timestamp 1698431365
transform 1 0 17696 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].vref_I
timestamp 1698431365
transform 1 0 16128 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref_I
timestamp 1698431365
transform 1 0 15120 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[2\].vref_I
timestamp 1698431365
transform 1 0 16240 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].vref_I
timestamp 1698431365
transform 1 0 15120 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch._4__A2
timestamp 1698431365
transform 1 0 14336 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch._5__A1
timestamp 1698431365
transform 1 0 12880 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch._7__I
timestamp 1698431365
transform 1 0 12096 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[0\].vref_I
timestamp 1698431365
transform 1 0 4704 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref_I
timestamp 1698431365
transform 1 0 4704 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[2\].vref_I
timestamp 1698431365
transform 1 0 7280 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[3\].vref_I
timestamp 1698431365
transform 1 0 5152 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref_I
timestamp 1698431365
transform 1 0 4704 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[5\].vref_I
timestamp 1698431365
transform 1 0 4704 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[6\].vref_I
timestamp 1698431365
transform 1 0 4704 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref_I
timestamp 1698431365
transform 1 0 4704 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch._4__A2
timestamp 1698431365
transform 1 0 24640 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch._5__A1
timestamp 1698431365
transform 1 0 28224 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch._7__I
timestamp 1698431365
transform -1 0 10080 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[0\].vref_I
timestamp 1698431365
transform 1 0 6272 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[1\].vref_I
timestamp 1698431365
transform 1 0 9632 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref_I
timestamp 1698431365
transform 1 0 10080 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[3\].vref_I
timestamp 1698431365
transform 1 0 4816 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[4\].vref_I
timestamp 1698431365
transform 1 0 11984 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[5\].vref_I
timestamp 1698431365
transform 1 0 5712 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[6\].vref_I
timestamp 1698431365
transform 1 0 5600 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].vref_I
timestamp 1698431365
transform 1 0 9632 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].vref_I
timestamp 1698431365
transform 1 0 4592 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[9\].vref_I
timestamp 1698431365
transform 1 0 5712 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[10\].vref_I
timestamp 1698431365
transform 1 0 5712 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[11\].vref_I
timestamp 1698431365
transform 1 0 5712 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref_I
timestamp 1698431365
transform 1 0 8848 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].vref_I
timestamp 1698431365
transform 1 0 5712 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[14\].vref_I
timestamp 1698431365
transform 1 0 9632 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].vref_I
timestamp 1698431365
transform 1 0 9632 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.vdac_single.einvp_batch\[0\].vref_I
timestamp 1698431365
transform 1 0 14672 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dcdc_EN
timestamp 1698431365
transform 1 0 21616 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_wire4_I
timestamp 1698431365
transform 1 0 7616 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_wire5_I
timestamp 1698431365
transform 1 0 11312 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0__0385_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19040 0 -1 83104
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0__0387_
timestamp 1698431365
transform 1 0 18480 0 -1 76832
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0__0737_
timestamp 1698431365
transform 1 0 21952 0 1 79968
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0__0750_
timestamp 1698431365
transform 1 0 23184 0 1 75264
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk
timestamp 1698431365
transform 1 0 21168 0 1 47040
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_net66
timestamp 1698431365
transform 1 0 22512 0 1 84672
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_temp1.i_precharge_n
timestamp 1698431365
transform 1 0 25088 0 -1 89376
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f__0385_
timestamp 1698431365
transform -1 0 24416 0 -1 78400
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f__0387_
timestamp 1698431365
transform -1 0 20944 0 1 76832
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f__0737_
timestamp 1698431365
transform -1 0 26768 0 1 76832
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f__0750_
timestamp 1698431365
transform -1 0 27440 0 1 73696
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_net66
timestamp 1698431365
transform -1 0 26768 0 1 81536
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_temp1.i_precharge_n
timestamp 1698431365
transform -1 0 31136 0 -1 86240
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f__0385_
timestamp 1698431365
transform -1 0 24864 0 -1 86240
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f__0387_
timestamp 1698431365
transform 1 0 19264 0 -1 73696
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f__0737_
timestamp 1698431365
transform 1 0 23184 0 1 83104
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f__0750_
timestamp 1698431365
transform 1 0 25088 0 -1 79968
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_net66
timestamp 1698431365
transform 1 0 25088 0 -1 87808
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_temp1.i_precharge_n
timestamp 1698431365
transform -1 0 28112 0 1 90944
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1698431365
transform -1 0 15232 0 -1 67424
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1698431365
transform -1 0 20160 0 1 72128
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1698431365
transform -1 0 28000 0 1 72128
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1698431365
transform 1 0 26544 0 -1 72128
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  dec1._060_
timestamp 1698431365
transform 1 0 32928 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  dec1._061_
timestamp 1698431365
transform 1 0 33152 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  dec1._062_
timestamp 1698431365
transform -1 0 36624 0 1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  dec1._063_
timestamp 1698431365
transform 1 0 32928 0 -1 59584
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  dec1._064_
timestamp 1698431365
transform 1 0 32256 0 1 61152
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  dec1._065_
timestamp 1698431365
transform -1 0 32704 0 -1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  dec1._066_
timestamp 1698431365
transform 1 0 31248 0 1 61152
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  dec1._067_
timestamp 1698431365
transform -1 0 33712 0 1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  dec1._068_
timestamp 1698431365
transform 1 0 33376 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  dec1._069_
timestamp 1698431365
transform 1 0 32256 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  dec1._070_
timestamp 1698431365
transform -1 0 36400 0 1 58016
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__inv_3  dec1._071_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 37744 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  dec1._072_
timestamp 1698431365
transform -1 0 37632 0 -1 59584
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  dec1._073_
timestamp 1698431365
transform -1 0 38192 0 -1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  dec1._074_
timestamp 1698431365
transform 1 0 32704 0 1 59584
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  dec1._075_
timestamp 1698431365
transform 1 0 36848 0 1 58016
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  dec1._076_
timestamp 1698431365
transform -1 0 32704 0 -1 62720
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  dec1._077_
timestamp 1698431365
transform -1 0 36624 0 1 61152
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  dec1._078_
timestamp 1698431365
transform -1 0 38416 0 1 62720
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  dec1._079_
timestamp 1698431365
transform -1 0 36624 0 1 59584
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  dec1._080_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 32928 0 -1 61152
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  dec1._081_
timestamp 1698431365
transform 1 0 31808 0 1 62720
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  dec1._082_
timestamp 1698431365
transform 1 0 33152 0 -1 58016
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  dec1._083_
timestamp 1698431365
transform -1 0 34272 0 1 64288
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  dec1._084_
timestamp 1698431365
transform -1 0 38416 0 1 59584
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  dec1._085_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 37744 0 -1 62720
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  dec1._086_
timestamp 1698431365
transform 1 0 33040 0 -1 64288
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  dec1._087_
timestamp 1698431365
transform -1 0 38304 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and3_2  dec1._088_
timestamp 1698431365
transform 1 0 36848 0 1 61152
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  dec1._089_
timestamp 1698431365
transform 1 0 34496 0 1 56448
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  dec1._090_
timestamp 1698431365
transform 1 0 35056 0 -1 58016
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  dec1._091_
timestamp 1698431365
transform -1 0 37856 0 1 64288
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  dec1._092_
timestamp 1698431365
transform 1 0 35056 0 1 64288
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  dec1._093_
timestamp 1698431365
transform -1 0 36624 0 1 65856
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  dec1._094_
timestamp 1698431365
transform 1 0 34384 0 -1 61152
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  dec1._095_
timestamp 1698431365
transform 1 0 31808 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  dec1._096_
timestamp 1698431365
transform 1 0 31920 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  dec1._097_
timestamp 1698431365
transform -1 0 37744 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  dec1._098_
timestamp 1698431365
transform 1 0 34832 0 1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  dec1._099_
timestamp 1698431365
transform 1 0 35728 0 -1 64288
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  dec1._100_
timestamp 1698431365
transform 1 0 35392 0 -1 65856
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  dec1._101_
timestamp 1698431365
transform -1 0 35168 0 -1 72128
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  dec1._102_
timestamp 1698431365
transform -1 0 37632 0 -1 70560
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  dec1._103_
timestamp 1698431365
transform -1 0 32704 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  dec1._104_
timestamp 1698431365
transform -1 0 32704 0 -1 65856
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  dec1._105_
timestamp 1698431365
transform -1 0 33376 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  dec1._106_
timestamp 1698431365
transform -1 0 32704 0 -1 68992
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  dec1._107_
timestamp 1698431365
transform -1 0 35056 0 1 67424
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  dec1._108_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 33936 0 -1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  dec1._109_
timestamp 1698431365
transform -1 0 33712 0 -1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  dec1._110_
timestamp 1698431365
transform -1 0 38416 0 1 64288
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  dec1._111_
timestamp 1698431365
transform -1 0 35392 0 -1 65856
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  dec1._112_
timestamp 1698431365
transform 1 0 32480 0 1 68992
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  dec1._113_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 33936 0 -1 67424
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  dec1._114_
timestamp 1698431365
transform 1 0 33936 0 1 68992
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  dec1._115_
timestamp 1698431365
transform -1 0 33712 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  dec1._116_
timestamp 1698431365
transform 1 0 36848 0 1 68992
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  dec1._117_
timestamp 1698431365
transform -1 0 36512 0 1 67424
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  dec1._118_
timestamp 1698431365
transform -1 0 34608 0 -1 72128
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  dec1._119_
timestamp 1698431365
transform -1 0 38416 0 -1 68992
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  dec1._120_
timestamp 1698431365
transform 1 0 34272 0 1 64288
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  dec1._121_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 37968 0 1 67424
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  dec1._122_
timestamp 1698431365
transform -1 0 36512 0 -1 72128
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  dec1._123_
timestamp 1698431365
transform 1 0 32928 0 -1 70560
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout43
timestamp 1698431365
transform 1 0 15456 0 -1 10976
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout44
timestamp 1698431365
transform 1 0 18480 0 1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout45
timestamp 1698431365
transform 1 0 17136 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout46
timestamp 1698431365
transform 1 0 29232 0 1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout47
timestamp 1698431365
transform 1 0 35056 0 1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  fanout48
timestamp 1698431365
transform 1 0 29456 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout49
timestamp 1698431365
transform 1 0 13440 0 -1 40768
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout50
timestamp 1698431365
transform 1 0 14000 0 -1 58016
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  fanout51
timestamp 1698431365
transform -1 0 16576 0 1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout52
timestamp 1698431365
transform -1 0 36624 0 1 37632
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout53
timestamp 1698431365
transform 1 0 36848 0 1 39200
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_2 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 1568
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_10 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2464 0 1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_14 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2912 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_16 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3136 0 1 1568
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_19
timestamp 1698431365
transform 1 0 3472 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_29
timestamp 1698431365
transform 1 0 4592 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_31
timestamp 1698431365
transform 1 0 4816 0 1 1568
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_36
timestamp 1698431365
transform 1 0 5376 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_38
timestamp 1698431365
transform 1 0 5600 0 1 1568
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_45
timestamp 1698431365
transform 1 0 6384 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_53
timestamp 1698431365
transform 1 0 7280 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_61
timestamp 1698431365
transform 1 0 8176 0 1 1568
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 1568
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_77
timestamp 1698431365
transform 1 0 9968 0 1 1568
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_138
timestamp 1698431365
transform 1 0 16800 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_140
timestamp 1698431365
transform 1 0 17024 0 1 1568
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_149
timestamp 1698431365
transform 1 0 18032 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_157
timestamp 1698431365
transform 1 0 18928 0 1 1568
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_172
timestamp 1698431365
transform 1 0 20608 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_174
timestamp 1698431365
transform 1 0 20832 0 1 1568
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_181
timestamp 1698431365
transform 1 0 21616 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_189
timestamp 1698431365
transform 1 0 22512 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_197
timestamp 1698431365
transform 1 0 23408 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_201
timestamp 1698431365
transform 1 0 23856 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_203
timestamp 1698431365
transform 1 0 24080 0 1 1568
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_230
timestamp 1698431365
transform 1 0 27104 0 1 1568
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_237
timestamp 1698431365
transform 1 0 27888 0 1 1568
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_246
timestamp 1698431365
transform 1 0 28896 0 1 1568
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_253
timestamp 1698431365
transform 1 0 29680 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_261
timestamp 1698431365
transform 1 0 30576 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_269
timestamp 1698431365
transform 1 0 31472 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_271
timestamp 1698431365
transform 1 0 31696 0 1 1568
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_286
timestamp 1698431365
transform 1 0 33376 0 1 1568
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_293
timestamp 1698431365
transform 1 0 34160 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_301
timestamp 1698431365
transform 1 0 35056 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_305
timestamp 1698431365
transform 1 0 35504 0 1 1568
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_320
timestamp 1698431365
transform 1 0 37184 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_324
timestamp 1698431365
transform 1 0 37632 0 1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_328
timestamp 1698431365
transform 1 0 38080 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_330
timestamp 1698431365
transform 1 0 38304 0 1 1568
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_2 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_18
timestamp 1698431365
transform 1 0 3360 0 -1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_26
timestamp 1698431365
transform 1 0 4256 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_54
timestamp 1698431365
transform 1 0 7392 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_58
timestamp 1698431365
transform 1 0 7840 0 -1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_62
timestamp 1698431365
transform 1 0 8288 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_66
timestamp 1698431365
transform 1 0 8736 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_94
timestamp 1698431365
transform 1 0 11872 0 -1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_137
timestamp 1698431365
transform 1 0 16688 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_139
timestamp 1698431365
transform 1 0 16912 0 -1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_148
timestamp 1698431365
transform 1 0 17920 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_152
timestamp 1698431365
transform 1 0 18368 0 -1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_156
timestamp 1698431365
transform 1 0 18816 0 -1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_159
timestamp 1698431365
transform 1 0 19152 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_200
timestamp 1698431365
transform 1 0 23744 0 -1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_206
timestamp 1698431365
transform 1 0 24416 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_230
timestamp 1698431365
transform 1 0 27104 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_234
timestamp 1698431365
transform 1 0 27552 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_238
timestamp 1698431365
transform 1 0 28000 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_242
timestamp 1698431365
transform 1 0 28448 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_244
timestamp 1698431365
transform 1 0 28672 0 -1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_247
timestamp 1698431365
transform 1 0 29008 0 -1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_251
timestamp 1698431365
transform 1 0 29456 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_255
timestamp 1698431365
transform 1 0 29904 0 -1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_259
timestamp 1698431365
transform 1 0 30352 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_263
timestamp 1698431365
transform 1 0 30800 0 -1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_271
timestamp 1698431365
transform 1 0 31696 0 -1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_274
timestamp 1698431365
transform 1 0 32032 0 -1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_308
timestamp 1698431365
transform 1 0 35840 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_312
timestamp 1698431365
transform 1 0 36288 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_316
timestamp 1698431365
transform 1 0 36736 0 -1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_324
timestamp 1698431365
transform 1 0 37632 0 -1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_328
timestamp 1698431365
transform 1 0 38080 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_330
timestamp 1698431365
transform 1 0 38304 0 -1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_41
timestamp 1698431365
transform 1 0 5936 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_46
timestamp 1698431365
transform 1 0 6496 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_88
timestamp 1698431365
transform 1 0 11200 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_92
timestamp 1698431365
transform 1 0 11648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_98
timestamp 1698431365
transform 1 0 12320 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_102
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_104
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_117
timestamp 1698431365
transform 1 0 14448 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_167
timestamp 1698431365
transform 1 0 20048 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_171
timestamp 1698431365
transform 1 0 20496 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_185
timestamp 1698431365
transform 1 0 22064 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_191
timestamp 1698431365
transform 1 0 22736 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_222
timestamp 1698431365
transform 1 0 26208 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_226
timestamp 1698431365
transform 1 0 26656 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_247
timestamp 1698431365
transform 1 0 29008 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_263
timestamp 1698431365
transform 1 0 30800 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_301
timestamp 1698431365
transform 1 0 35056 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_309
timestamp 1698431365
transform 1 0 35952 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_313
timestamp 1698431365
transform 1 0 36400 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_317
timestamp 1698431365
transform 1 0 36848 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_325
timestamp 1698431365
transform 1 0 37744 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_329
timestamp 1698431365
transform 1 0 38192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_34
timestamp 1698431365
transform 1 0 5152 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_36
timestamp 1698431365
transform 1 0 5376 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_66
timestamp 1698431365
transform 1 0 8736 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_74
timestamp 1698431365
transform 1 0 9632 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_82
timestamp 1698431365
transform 1 0 10528 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_120
timestamp 1698431365
transform 1 0 14784 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_124
timestamp 1698431365
transform 1 0 15232 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_134
timestamp 1698431365
transform 1 0 16352 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_150
timestamp 1698431365
transform 1 0 18144 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_154
timestamp 1698431365
transform 1 0 18592 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_156
timestamp 1698431365
transform 1 0 18816 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_194
timestamp 1698431365
transform 1 0 23072 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_198
timestamp 1698431365
transform 1 0 23520 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_202
timestamp 1698431365
transform 1 0 23968 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_221
timestamp 1698431365
transform 1 0 26096 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_223
timestamp 1698431365
transform 1 0 26320 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_226
timestamp 1698431365
transform 1 0 26656 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_258
timestamp 1698431365
transform 1 0 30240 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_274
timestamp 1698431365
transform 1 0 32032 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_278
timestamp 1698431365
transform 1 0 32480 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_282
timestamp 1698431365
transform 1 0 32928 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_286
timestamp 1698431365
transform 1 0 33376 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_288
timestamp 1698431365
transform 1 0 33600 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_303
timestamp 1698431365
transform 1 0 35280 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_319
timestamp 1698431365
transform 1 0 37072 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_327
timestamp 1698431365
transform 1 0 37968 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_53
timestamp 1698431365
transform 1 0 7280 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_57
timestamp 1698431365
transform 1 0 7728 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_69
timestamp 1698431365
transform 1 0 9072 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_73
timestamp 1698431365
transform 1 0 9520 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_77
timestamp 1698431365
transform 1 0 9968 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_80
timestamp 1698431365
transform 1 0 10304 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_88
timestamp 1698431365
transform 1 0 11200 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_92
timestamp 1698431365
transform 1 0 11648 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_99
timestamp 1698431365
transform 1 0 12432 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_103
timestamp 1698431365
transform 1 0 12880 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_111
timestamp 1698431365
transform 1 0 13776 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_120
timestamp 1698431365
transform 1 0 14784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_161
timestamp 1698431365
transform 1 0 19376 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_163
timestamp 1698431365
transform 1 0 19600 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_174
timestamp 1698431365
transform 1 0 20832 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_191
timestamp 1698431365
transform 1 0 22736 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_195
timestamp 1698431365
transform 1 0 23184 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_231
timestamp 1698431365
transform 1 0 27216 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_235
timestamp 1698431365
transform 1 0 27664 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_243
timestamp 1698431365
transform 1 0 28560 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698431365
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_317
timestamp 1698431365
transform 1 0 36848 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_325
timestamp 1698431365
transform 1 0 37744 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_329
timestamp 1698431365
transform 1 0 38192 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698431365
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_101
timestamp 1698431365
transform 1 0 12656 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_131
timestamp 1698431365
transform 1 0 16016 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_135
timestamp 1698431365
transform 1 0 16464 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_139
timestamp 1698431365
transform 1 0 16912 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_148
timestamp 1698431365
transform 1 0 17920 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_152
timestamp 1698431365
transform 1 0 18368 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_154
timestamp 1698431365
transform 1 0 18592 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_184
timestamp 1698431365
transform 1 0 21952 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_199
timestamp 1698431365
transform 1 0 23632 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_208
timestamp 1698431365
transform 1 0 24640 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_220
timestamp 1698431365
transform 1 0 25984 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_252
timestamp 1698431365
transform 1 0 29568 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_268
timestamp 1698431365
transform 1 0 31360 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698431365
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_282
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_314
timestamp 1698431365
transform 1 0 36512 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_330
timestamp 1698431365
transform 1 0 38304 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_45
timestamp 1698431365
transform 1 0 6384 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_49
timestamp 1698431365
transform 1 0 6832 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_88
timestamp 1698431365
transform 1 0 11200 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_100
timestamp 1698431365
transform 1 0 12544 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_104
timestamp 1698431365
transform 1 0 12992 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_109
timestamp 1698431365
transform 1 0 13552 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_149
timestamp 1698431365
transform 1 0 18032 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_153
timestamp 1698431365
transform 1 0 18480 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_169
timestamp 1698431365
transform 1 0 20272 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_173
timestamp 1698431365
transform 1 0 20720 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_181
timestamp 1698431365
transform 1 0 21616 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_185
timestamp 1698431365
transform 1 0 22064 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_189
timestamp 1698431365
transform 1 0 22512 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_197
timestamp 1698431365
transform 1 0 23408 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_200
timestamp 1698431365
transform 1 0 23744 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_208
timestamp 1698431365
transform 1 0 24640 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_212
timestamp 1698431365
transform 1 0 25088 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_244
timestamp 1698431365
transform 1 0 28672 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_247
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_255
timestamp 1698431365
transform 1 0 29904 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_261
timestamp 1698431365
transform 1 0 30576 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_293
timestamp 1698431365
transform 1 0 34160 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_309
timestamp 1698431365
transform 1 0 35952 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_313
timestamp 1698431365
transform 1 0 36400 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_317
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_325
timestamp 1698431365
transform 1 0 37744 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_329
timestamp 1698431365
transform 1 0 38192 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_34
timestamp 1698431365
transform 1 0 5152 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_52
timestamp 1698431365
transform 1 0 7168 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_56
timestamp 1698431365
transform 1 0 7616 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_64
timestamp 1698431365
transform 1 0 8512 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_68
timestamp 1698431365
transform 1 0 8960 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_74
timestamp 1698431365
transform 1 0 9632 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_81
timestamp 1698431365
transform 1 0 10416 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_85
timestamp 1698431365
transform 1 0 10864 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_115
timestamp 1698431365
transform 1 0 14224 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_119
timestamp 1698431365
transform 1 0 14672 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_135
timestamp 1698431365
transform 1 0 16464 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_139
timestamp 1698431365
transform 1 0 16912 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_150
timestamp 1698431365
transform 1 0 18144 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_154
timestamp 1698431365
transform 1 0 18592 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_156
timestamp 1698431365
transform 1 0 18816 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_186
timestamp 1698431365
transform 1 0 22176 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_190
timestamp 1698431365
transform 1 0 22624 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698431365
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_220
timestamp 1698431365
transform 1 0 25984 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_265
timestamp 1698431365
transform 1 0 31024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_269
timestamp 1698431365
transform 1 0 31472 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_277
timestamp 1698431365
transform 1 0 32368 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_279
timestamp 1698431365
transform 1 0 32592 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_282
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_314
timestamp 1698431365
transform 1 0 36512 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_330
timestamp 1698431365
transform 1 0 38304 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_53
timestamp 1698431365
transform 1 0 7280 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_61
timestamp 1698431365
transform 1 0 8176 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_69
timestamp 1698431365
transform 1 0 9072 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698431365
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_123
timestamp 1698431365
transform 1 0 15120 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_127
timestamp 1698431365
transform 1 0 15568 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_129
timestamp 1698431365
transform 1 0 15792 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_132
timestamp 1698431365
transform 1 0 16128 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_164
timestamp 1698431365
transform 1 0 19712 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_172
timestamp 1698431365
transform 1 0 20608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_174
timestamp 1698431365
transform 1 0 20832 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_209
timestamp 1698431365
transform 1 0 24752 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_211
timestamp 1698431365
transform 1 0 24976 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_236
timestamp 1698431365
transform 1 0 27776 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_240
timestamp 1698431365
transform 1 0 28224 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_244
timestamp 1698431365
transform 1 0 28672 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_247
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_271
timestamp 1698431365
transform 1 0 31696 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_275
timestamp 1698431365
transform 1 0 32144 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_307
timestamp 1698431365
transform 1 0 35728 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_317
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_325
timestamp 1698431365
transform 1 0 37744 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_34
timestamp 1698431365
transform 1 0 5152 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_37
timestamp 1698431365
transform 1 0 5488 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_53
timestamp 1698431365
transform 1 0 7280 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_61
timestamp 1698431365
transform 1 0 8176 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_65
timestamp 1698431365
transform 1 0 8624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_67
timestamp 1698431365
transform 1 0 8848 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_80
timestamp 1698431365
transform 1 0 10304 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_112
timestamp 1698431365
transform 1 0 13888 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_120
timestamp 1698431365
transform 1 0 14784 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_130
timestamp 1698431365
transform 1 0 15904 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_146
timestamp 1698431365
transform 1 0 17696 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_148
timestamp 1698431365
transform 1 0 17920 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_151
timestamp 1698431365
transform 1 0 18256 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_159
timestamp 1698431365
transform 1 0 19152 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_163
timestamp 1698431365
transform 1 0 19600 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_166
timestamp 1698431365
transform 1 0 19936 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_173
timestamp 1698431365
transform 1 0 20720 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_205
timestamp 1698431365
transform 1 0 24304 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_209
timestamp 1698431365
transform 1 0 24752 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_242
timestamp 1698431365
transform 1 0 28448 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_246
timestamp 1698431365
transform 1 0 28896 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_276
timestamp 1698431365
transform 1 0 32256 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_282
timestamp 1698431365
transform 1 0 32928 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_314
timestamp 1698431365
transform 1 0 36512 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_316
timestamp 1698431365
transform 1 0 36736 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_18
timestamp 1698431365
transform 1 0 3360 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_26
timestamp 1698431365
transform 1 0 4256 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_28
timestamp 1698431365
transform 1 0 4480 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_63
timestamp 1698431365
transform 1 0 8400 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_79
timestamp 1698431365
transform 1 0 10192 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_89
timestamp 1698431365
transform 1 0 11312 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_93
timestamp 1698431365
transform 1 0 11760 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_97
timestamp 1698431365
transform 1 0 12208 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_136
timestamp 1698431365
transform 1 0 16576 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_149
timestamp 1698431365
transform 1 0 18032 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_153
timestamp 1698431365
transform 1 0 18480 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_155
timestamp 1698431365
transform 1 0 18704 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_158
timestamp 1698431365
transform 1 0 19040 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_162
timestamp 1698431365
transform 1 0 19488 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_174
timestamp 1698431365
transform 1 0 20832 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_177
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_231
timestamp 1698431365
transform 1 0 27216 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_235
timestamp 1698431365
transform 1 0 27664 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_239
timestamp 1698431365
transform 1 0 28112 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_243
timestamp 1698431365
transform 1 0 28560 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_247
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_261
timestamp 1698431365
transform 1 0 30576 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_273
timestamp 1698431365
transform 1 0 31920 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_277
timestamp 1698431365
transform 1 0 32368 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_309
timestamp 1698431365
transform 1 0 35952 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_313
timestamp 1698431365
transform 1 0 36400 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_317
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_325
timestamp 1698431365
transform 1 0 37744 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_329
timestamp 1698431365
transform 1 0 38192 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_18
timestamp 1698431365
transform 1 0 3360 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_22
timestamp 1698431365
transform 1 0 3808 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_66
timestamp 1698431365
transform 1 0 8736 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_87
timestamp 1698431365
transform 1 0 11088 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_91
timestamp 1698431365
transform 1 0 11536 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_124
timestamp 1698431365
transform 1 0 15232 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_146
timestamp 1698431365
transform 1 0 17696 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_158
timestamp 1698431365
transform 1 0 19040 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_178
timestamp 1698431365
transform 1 0 21280 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_190
timestamp 1698431365
transform 1 0 22624 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_194
timestamp 1698431365
transform 1 0 23072 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_202
timestamp 1698431365
transform 1 0 23968 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_206
timestamp 1698431365
transform 1 0 24416 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_221
timestamp 1698431365
transform 1 0 26096 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_240
timestamp 1698431365
transform 1 0 28224 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_256
timestamp 1698431365
transform 1 0 30016 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_270
timestamp 1698431365
transform 1 0 31584 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_278
timestamp 1698431365
transform 1 0 32480 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_282
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_314
timestamp 1698431365
transform 1 0 36512 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_330
timestamp 1698431365
transform 1 0 38304 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_63
timestamp 1698431365
transform 1 0 8400 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_67
timestamp 1698431365
transform 1 0 8848 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_97
timestamp 1698431365
transform 1 0 12208 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_101
timestamp 1698431365
transform 1 0 12656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_111
timestamp 1698431365
transform 1 0 13776 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_113
timestamp 1698431365
transform 1 0 14000 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_157
timestamp 1698431365
transform 1 0 18928 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_170
timestamp 1698431365
transform 1 0 20384 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_172
timestamp 1698431365
transform 1 0 20608 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_191
timestamp 1698431365
transform 1 0 22736 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_199
timestamp 1698431365
transform 1 0 23632 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_201
timestamp 1698431365
transform 1 0 23856 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_208
timestamp 1698431365
transform 1 0 24640 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_216
timestamp 1698431365
transform 1 0 25536 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_218
timestamp 1698431365
transform 1 0 25760 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_221
timestamp 1698431365
transform 1 0 26096 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_225
timestamp 1698431365
transform 1 0 26544 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_229
timestamp 1698431365
transform 1 0 26992 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_232
timestamp 1698431365
transform 1 0 27328 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_240
timestamp 1698431365
transform 1 0 28224 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_244
timestamp 1698431365
transform 1 0 28672 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_247
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_286
timestamp 1698431365
transform 1 0 33376 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_302
timestamp 1698431365
transform 1 0 35168 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_310
timestamp 1698431365
transform 1 0 36064 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_314
timestamp 1698431365
transform 1 0 36512 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_317
timestamp 1698431365
transform 1 0 36848 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_325
timestamp 1698431365
transform 1 0 37744 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_329
timestamp 1698431365
transform 1 0 38192 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_2
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_34
timestamp 1698431365
transform 1 0 5152 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_38
timestamp 1698431365
transform 1 0 5600 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_54
timestamp 1698431365
transform 1 0 7392 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_58
timestamp 1698431365
transform 1 0 7840 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_80
timestamp 1698431365
transform 1 0 10304 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_88
timestamp 1698431365
transform 1 0 11200 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_92
timestamp 1698431365
transform 1 0 11648 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_103
timestamp 1698431365
transform 1 0 12880 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_109
timestamp 1698431365
transform 1 0 13552 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_113
timestamp 1698431365
transform 1 0 14000 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_121
timestamp 1698431365
transform 1 0 14896 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_124
timestamp 1698431365
transform 1 0 15232 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_128
timestamp 1698431365
transform 1 0 15680 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_138
timestamp 1698431365
transform 1 0 16800 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_162
timestamp 1698431365
transform 1 0 19488 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_166
timestamp 1698431365
transform 1 0 19936 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_170
timestamp 1698431365
transform 1 0 20384 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_172
timestamp 1698431365
transform 1 0 20608 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_202
timestamp 1698431365
transform 1 0 23968 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_206
timestamp 1698431365
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_212
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_220
timestamp 1698431365
transform 1 0 25984 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_224
timestamp 1698431365
transform 1 0 26432 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_255
timestamp 1698431365
transform 1 0 29904 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_259
timestamp 1698431365
transform 1 0 30352 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_275
timestamp 1698431365
transform 1 0 32144 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_279
timestamp 1698431365
transform 1 0 32592 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_282
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_314
timestamp 1698431365
transform 1 0 36512 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_330
timestamp 1698431365
transform 1 0 38304 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_45
timestamp 1698431365
transform 1 0 6384 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_49
timestamp 1698431365
transform 1 0 6832 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_51
timestamp 1698431365
transform 1 0 7056 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_83
timestamp 1698431365
transform 1 0 10640 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_87
timestamp 1698431365
transform 1 0 11088 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_103
timestamp 1698431365
transform 1 0 12880 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_113
timestamp 1698431365
transform 1 0 14000 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_129
timestamp 1698431365
transform 1 0 15792 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_137
timestamp 1698431365
transform 1 0 16688 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_139
timestamp 1698431365
transform 1 0 16912 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_142
timestamp 1698431365
transform 1 0 17248 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_146
timestamp 1698431365
transform 1 0 17696 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_150
timestamp 1698431365
transform 1 0 18144 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_153
timestamp 1698431365
transform 1 0 18480 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_159
timestamp 1698431365
transform 1 0 19152 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_193
timestamp 1698431365
transform 1 0 22960 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_201
timestamp 1698431365
transform 1 0 23856 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_211
timestamp 1698431365
transform 1 0 24976 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_215
timestamp 1698431365
transform 1 0 25424 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_231
timestamp 1698431365
transform 1 0 27216 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_239
timestamp 1698431365
transform 1 0 28112 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_243
timestamp 1698431365
transform 1 0 28560 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_247
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_255
timestamp 1698431365
transform 1 0 29904 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_257
timestamp 1698431365
transform 1 0 30128 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_274
timestamp 1698431365
transform 1 0 32032 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_306
timestamp 1698431365
transform 1 0 35616 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_314
timestamp 1698431365
transform 1 0 36512 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_317
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_325
timestamp 1698431365
transform 1 0 37744 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_329
timestamp 1698431365
transform 1 0 38192 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_2
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_18
timestamp 1698431365
transform 1 0 3360 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_26
timestamp 1698431365
transform 1 0 4256 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_57
timestamp 1698431365
transform 1 0 7728 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_61
timestamp 1698431365
transform 1 0 8176 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_69
timestamp 1698431365
transform 1 0 9072 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_78
timestamp 1698431365
transform 1 0 10080 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_110
timestamp 1698431365
transform 1 0 13664 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_126
timestamp 1698431365
transform 1 0 15456 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_134
timestamp 1698431365
transform 1 0 16352 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_138
timestamp 1698431365
transform 1 0 16800 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_152
timestamp 1698431365
transform 1 0 18368 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_156
timestamp 1698431365
transform 1 0 18816 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_188
timestamp 1698431365
transform 1 0 22400 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_204
timestamp 1698431365
transform 1 0 24192 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_208
timestamp 1698431365
transform 1 0 24640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_212
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_216
timestamp 1698431365
transform 1 0 25536 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_248
timestamp 1698431365
transform 1 0 29120 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_264
timestamp 1698431365
transform 1 0 30912 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_268
timestamp 1698431365
transform 1 0 31360 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_271
timestamp 1698431365
transform 1 0 31696 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_279
timestamp 1698431365
transform 1 0 32592 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_288
timestamp 1698431365
transform 1 0 33600 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_320
timestamp 1698431365
transform 1 0 37184 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_328
timestamp 1698431365
transform 1 0 38080 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_330
timestamp 1698431365
transform 1 0 38304 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698431365
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_39
timestamp 1698431365
transform 1 0 5712 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_46
timestamp 1698431365
transform 1 0 6496 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_78
timestamp 1698431365
transform 1 0 10080 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_94
timestamp 1698431365
transform 1 0 11872 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_102
timestamp 1698431365
transform 1 0 12768 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_104
timestamp 1698431365
transform 1 0 12992 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_111
timestamp 1698431365
transform 1 0 13776 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_121
timestamp 1698431365
transform 1 0 14896 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_125
timestamp 1698431365
transform 1 0 15344 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_141
timestamp 1698431365
transform 1 0 17136 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_148
timestamp 1698431365
transform 1 0 17920 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_156
timestamp 1698431365
transform 1 0 18816 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_159
timestamp 1698431365
transform 1 0 19152 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_177
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_210
timestamp 1698431365
transform 1 0 24864 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_214
timestamp 1698431365
transform 1 0 25312 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_217
timestamp 1698431365
transform 1 0 25648 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_221
timestamp 1698431365
transform 1 0 26096 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_223
timestamp 1698431365
transform 1 0 26320 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_234
timestamp 1698431365
transform 1 0 27552 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_242
timestamp 1698431365
transform 1 0 28448 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_244
timestamp 1698431365
transform 1 0 28672 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_247
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_254
timestamp 1698431365
transform 1 0 29792 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_258
timestamp 1698431365
transform 1 0 30240 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_260
timestamp 1698431365
transform 1 0 30464 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_300
timestamp 1698431365
transform 1 0 34944 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_308
timestamp 1698431365
transform 1 0 35840 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_312
timestamp 1698431365
transform 1 0 36288 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_314
timestamp 1698431365
transform 1 0 36512 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_317
timestamp 1698431365
transform 1 0 36848 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_325
timestamp 1698431365
transform 1 0 37744 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_329
timestamp 1698431365
transform 1 0 38192 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_2
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_34
timestamp 1698431365
transform 1 0 5152 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_42
timestamp 1698431365
transform 1 0 6048 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_44
timestamp 1698431365
transform 1 0 6272 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_53
timestamp 1698431365
transform 1 0 7280 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_57
timestamp 1698431365
transform 1 0 7728 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_65
timestamp 1698431365
transform 1 0 8624 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_67
timestamp 1698431365
transform 1 0 8848 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_72
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_74
timestamp 1698431365
transform 1 0 9632 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_83
timestamp 1698431365
transform 1 0 10640 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_91
timestamp 1698431365
transform 1 0 11536 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_94
timestamp 1698431365
transform 1 0 11872 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_98
timestamp 1698431365
transform 1 0 12320 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_100
timestamp 1698431365
transform 1 0 12544 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_103
timestamp 1698431365
transform 1 0 12880 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_133
timestamp 1698431365
transform 1 0 16240 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_137
timestamp 1698431365
transform 1 0 16688 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_139
timestamp 1698431365
transform 1 0 16912 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_153
timestamp 1698431365
transform 1 0 18480 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_167
timestamp 1698431365
transform 1 0 20048 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_171
timestamp 1698431365
transform 1 0 20496 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_175
timestamp 1698431365
transform 1 0 20944 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_185
timestamp 1698431365
transform 1 0 22064 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_192
timestamp 1698431365
transform 1 0 22848 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_196
timestamp 1698431365
transform 1 0 23296 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_198
timestamp 1698431365
transform 1 0 23520 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_208
timestamp 1698431365
transform 1 0 24640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_212
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_216
timestamp 1698431365
transform 1 0 25536 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_218
timestamp 1698431365
transform 1 0 25760 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_234
timestamp 1698431365
transform 1 0 27552 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_242
timestamp 1698431365
transform 1 0 28448 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_274
timestamp 1698431365
transform 1 0 32032 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_278
timestamp 1698431365
transform 1 0 32480 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_282
timestamp 1698431365
transform 1 0 32928 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_314
timestamp 1698431365
transform 1 0 36512 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_330
timestamp 1698431365
transform 1 0 38304 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698431365
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_53
timestamp 1698431365
transform 1 0 7280 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_61
timestamp 1698431365
transform 1 0 8176 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_101
timestamp 1698431365
transform 1 0 12656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_115
timestamp 1698431365
transform 1 0 14224 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_119
timestamp 1698431365
transform 1 0 14672 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_123
timestamp 1698431365
transform 1 0 15120 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_127
timestamp 1698431365
transform 1 0 15568 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_158
timestamp 1698431365
transform 1 0 19040 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_177
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_181
timestamp 1698431365
transform 1 0 21616 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_190
timestamp 1698431365
transform 1 0 22624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_194
timestamp 1698431365
transform 1 0 23072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_196
timestamp 1698431365
transform 1 0 23296 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_199
timestamp 1698431365
transform 1 0 23632 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_215
timestamp 1698431365
transform 1 0 25424 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_255
timestamp 1698431365
transform 1 0 29904 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_287
timestamp 1698431365
transform 1 0 33488 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_295
timestamp 1698431365
transform 1 0 34384 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_307
timestamp 1698431365
transform 1 0 35728 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_317
timestamp 1698431365
transform 1 0 36848 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_325
timestamp 1698431365
transform 1 0 37744 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_329
timestamp 1698431365
transform 1 0 38192 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_2
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_63
timestamp 1698431365
transform 1 0 8400 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_67
timestamp 1698431365
transform 1 0 8848 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_69
timestamp 1698431365
transform 1 0 9072 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_88
timestamp 1698431365
transform 1 0 11200 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_129
timestamp 1698431365
transform 1 0 15792 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_139
timestamp 1698431365
transform 1 0 16912 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_146
timestamp 1698431365
transform 1 0 17696 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_150
timestamp 1698431365
transform 1 0 18144 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_160
timestamp 1698431365
transform 1 0 19264 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_162
timestamp 1698431365
transform 1 0 19488 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_192
timestamp 1698431365
transform 1 0 22848 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_196
timestamp 1698431365
transform 1 0 23296 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_204
timestamp 1698431365
transform 1 0 24192 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_208
timestamp 1698431365
transform 1 0 24640 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_212
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_216
timestamp 1698431365
transform 1 0 25536 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_226
timestamp 1698431365
transform 1 0 26656 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_230
timestamp 1698431365
transform 1 0 27104 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_238
timestamp 1698431365
transform 1 0 28000 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_242
timestamp 1698431365
transform 1 0 28448 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_244
timestamp 1698431365
transform 1 0 28672 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_247
timestamp 1698431365
transform 1 0 29008 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_251
timestamp 1698431365
transform 1 0 29456 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_267
timestamp 1698431365
transform 1 0 31248 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_275
timestamp 1698431365
transform 1 0 32144 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_277
timestamp 1698431365
transform 1 0 32368 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_317
timestamp 1698431365
transform 1 0 36848 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_325
timestamp 1698431365
transform 1 0 37744 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_329
timestamp 1698431365
transform 1 0 38192 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_2
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_10
timestamp 1698431365
transform 1 0 2464 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_14
timestamp 1698431365
transform 1 0 2912 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_22
timestamp 1698431365
transform 1 0 3808 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_30
timestamp 1698431365
transform 1 0 4704 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_32
timestamp 1698431365
transform 1 0 4928 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_51
timestamp 1698431365
transform 1 0 7056 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_55
timestamp 1698431365
transform 1 0 7504 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_57
timestamp 1698431365
transform 1 0 7728 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_87
timestamp 1698431365
transform 1 0 11088 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_91
timestamp 1698431365
transform 1 0 11536 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_99
timestamp 1698431365
transform 1 0 12432 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_103
timestamp 1698431365
transform 1 0 12880 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_119
timestamp 1698431365
transform 1 0 14672 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_123
timestamp 1698431365
transform 1 0 15120 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_139
timestamp 1698431365
transform 1 0 16912 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_143
timestamp 1698431365
transform 1 0 17360 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_145
timestamp 1698431365
transform 1 0 17584 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_183
timestamp 1698431365
transform 1 0 21840 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_187
timestamp 1698431365
transform 1 0 22288 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_224
timestamp 1698431365
transform 1 0 26432 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_228
timestamp 1698431365
transform 1 0 26880 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_244
timestamp 1698431365
transform 1 0 28672 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_247
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_255
timestamp 1698431365
transform 1 0 29904 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_295
timestamp 1698431365
transform 1 0 34384 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_299
timestamp 1698431365
transform 1 0 34832 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_303
timestamp 1698431365
transform 1 0 35280 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698431365
transform 1 0 36176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_317
timestamp 1698431365
transform 1 0 36848 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_325
timestamp 1698431365
transform 1 0 37744 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_329
timestamp 1698431365
transform 1 0 38192 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_35
timestamp 1698431365
transform 1 0 5264 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_39
timestamp 1698431365
transform 1 0 5712 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_55
timestamp 1698431365
transform 1 0 7504 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_63
timestamp 1698431365
transform 1 0 8400 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_67
timestamp 1698431365
transform 1 0 8848 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_69
timestamp 1698431365
transform 1 0 9072 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_78
timestamp 1698431365
transform 1 0 10080 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_85
timestamp 1698431365
transform 1 0 10864 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_117
timestamp 1698431365
transform 1 0 14448 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_133
timestamp 1698431365
transform 1 0 16240 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_137
timestamp 1698431365
transform 1 0 16688 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_142
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_144
timestamp 1698431365
transform 1 0 17472 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_153
timestamp 1698431365
transform 1 0 18480 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_161
timestamp 1698431365
transform 1 0 19376 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_168
timestamp 1698431365
transform 1 0 20160 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_172
timestamp 1698431365
transform 1 0 20608 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_174
timestamp 1698431365
transform 1 0 20832 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_177
timestamp 1698431365
transform 1 0 21168 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_209
timestamp 1698431365
transform 1 0 24752 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_212
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_228
timestamp 1698431365
transform 1 0 26880 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_232
timestamp 1698431365
transform 1 0 27328 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_276
timestamp 1698431365
transform 1 0 32256 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_282
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_284
timestamp 1698431365
transform 1 0 33152 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_291
timestamp 1698431365
transform 1 0 33936 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_293
timestamp 1698431365
transform 1 0 34160 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_296
timestamp 1698431365
transform 1 0 34496 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_2
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_18
timestamp 1698431365
transform 1 0 3360 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_20
timestamp 1698431365
transform 1 0 3584 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_29
timestamp 1698431365
transform 1 0 4592 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_33
timestamp 1698431365
transform 1 0 5040 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698431365
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_136
timestamp 1698431365
transform 1 0 16576 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_140
timestamp 1698431365
transform 1 0 17024 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_144
timestamp 1698431365
transform 1 0 17472 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_160
timestamp 1698431365
transform 1 0 19264 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_168
timestamp 1698431365
transform 1 0 20160 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_172
timestamp 1698431365
transform 1 0 20608 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_174
timestamp 1698431365
transform 1 0 20832 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_177
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_228
timestamp 1698431365
transform 1 0 26880 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_232
timestamp 1698431365
transform 1 0 27328 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_240
timestamp 1698431365
transform 1 0 28224 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_244
timestamp 1698431365
transform 1 0 28672 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_247
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_251
timestamp 1698431365
transform 1 0 29456 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_255
timestamp 1698431365
transform 1 0 29904 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_266
timestamp 1698431365
transform 1 0 31136 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_270
timestamp 1698431365
transform 1 0 31584 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_274
timestamp 1698431365
transform 1 0 32032 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_276
timestamp 1698431365
transform 1 0 32256 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_279
timestamp 1698431365
transform 1 0 32592 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_283
timestamp 1698431365
transform 1 0 33040 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_294
timestamp 1698431365
transform 1 0 34272 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_312
timestamp 1698431365
transform 1 0 36288 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_314
timestamp 1698431365
transform 1 0 36512 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_323
timestamp 1698431365
transform 1 0 37520 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_6
timestamp 1698431365
transform 1 0 2016 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_8
timestamp 1698431365
transform 1 0 2240 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_38
timestamp 1698431365
transform 1 0 5600 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_42
timestamp 1698431365
transform 1 0 6048 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_58
timestamp 1698431365
transform 1 0 7840 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698431365
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_80
timestamp 1698431365
transform 1 0 10304 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_84
timestamp 1698431365
transform 1 0 10752 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_86
timestamp 1698431365
transform 1 0 10976 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_97
timestamp 1698431365
transform 1 0 12208 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_129
timestamp 1698431365
transform 1 0 15792 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_137
timestamp 1698431365
transform 1 0 16688 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_139
timestamp 1698431365
transform 1 0 16912 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_142
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_152
timestamp 1698431365
transform 1 0 18368 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_168
timestamp 1698431365
transform 1 0 20160 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_170
timestamp 1698431365
transform 1 0 20384 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_177
timestamp 1698431365
transform 1 0 21168 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_193
timestamp 1698431365
transform 1 0 22960 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_205
timestamp 1698431365
transform 1 0 24304 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_209
timestamp 1698431365
transform 1 0 24752 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_212
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_228
timestamp 1698431365
transform 1 0 26880 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_232
timestamp 1698431365
transform 1 0 27328 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_234
timestamp 1698431365
transform 1 0 27552 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_241
timestamp 1698431365
transform 1 0 28336 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_273
timestamp 1698431365
transform 1 0 31920 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_277
timestamp 1698431365
transform 1 0 32368 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1698431365
transform 1 0 32592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_282
timestamp 1698431365
transform 1 0 32928 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_284
timestamp 1698431365
transform 1 0 33152 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_287
timestamp 1698431365
transform 1 0 33488 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_291
timestamp 1698431365
transform 1 0 33936 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_18
timestamp 1698431365
transform 1 0 3360 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_20
timestamp 1698431365
transform 1 0 3584 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_27
timestamp 1698431365
transform 1 0 4368 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_31
timestamp 1698431365
transform 1 0 4816 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_52
timestamp 1698431365
transform 1 0 7168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_56
timestamp 1698431365
transform 1 0 7616 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_70
timestamp 1698431365
transform 1 0 9184 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_74
timestamp 1698431365
transform 1 0 9632 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_90
timestamp 1698431365
transform 1 0 11424 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_98
timestamp 1698431365
transform 1 0 12320 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_102
timestamp 1698431365
transform 1 0 12768 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_104
timestamp 1698431365
transform 1 0 12992 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_107
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_123
timestamp 1698431365
transform 1 0 15120 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_131
timestamp 1698431365
transform 1 0 16016 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_133
timestamp 1698431365
transform 1 0 16240 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_136
timestamp 1698431365
transform 1 0 16576 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_140
timestamp 1698431365
transform 1 0 17024 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_149
timestamp 1698431365
transform 1 0 18032 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_153
timestamp 1698431365
transform 1 0 18480 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_169
timestamp 1698431365
transform 1 0 20272 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_173
timestamp 1698431365
transform 1 0 20720 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_177
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_181
timestamp 1698431365
transform 1 0 21616 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_213
timestamp 1698431365
transform 1 0 25200 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_221
timestamp 1698431365
transform 1 0 26096 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_225
timestamp 1698431365
transform 1 0 26544 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_236
timestamp 1698431365
transform 1 0 27776 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_244
timestamp 1698431365
transform 1 0 28672 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_247
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_263
timestamp 1698431365
transform 1 0 30800 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_267
timestamp 1698431365
transform 1 0 31248 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_274
timestamp 1698431365
transform 1 0 32032 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_278
timestamp 1698431365
transform 1 0 32480 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_282
timestamp 1698431365
transform 1 0 32928 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_298
timestamp 1698431365
transform 1 0 34720 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_302
timestamp 1698431365
transform 1 0 35168 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_312
timestamp 1698431365
transform 1 0 36288 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_314
timestamp 1698431365
transform 1 0 36512 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_317
timestamp 1698431365
transform 1 0 36848 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_325
timestamp 1698431365
transform 1 0 37744 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_329
timestamp 1698431365
transform 1 0 38192 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_2
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_18
timestamp 1698431365
transform 1 0 3360 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_26
timestamp 1698431365
transform 1 0 4256 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_37
timestamp 1698431365
transform 1 0 5488 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_39
timestamp 1698431365
transform 1 0 5712 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_69
timestamp 1698431365
transform 1 0 9072 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_78
timestamp 1698431365
transform 1 0 10080 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_82
timestamp 1698431365
transform 1 0 10528 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_112
timestamp 1698431365
transform 1 0 13888 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_116
timestamp 1698431365
transform 1 0 14336 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_124
timestamp 1698431365
transform 1 0 15232 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_126
timestamp 1698431365
transform 1 0 15456 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_136
timestamp 1698431365
transform 1 0 16576 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_171
timestamp 1698431365
transform 1 0 20496 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_175
timestamp 1698431365
transform 1 0 20944 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_186
timestamp 1698431365
transform 1 0 22176 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_202
timestamp 1698431365
transform 1 0 23968 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_212
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_244
timestamp 1698431365
transform 1 0 28672 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_248
timestamp 1698431365
transform 1 0 29120 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_250
timestamp 1698431365
transform 1 0 29344 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_290
timestamp 1698431365
transform 1 0 33824 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_294
timestamp 1698431365
transform 1 0 34272 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_327
timestamp 1698431365
transform 1 0 37968 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_31
timestamp 1698431365
transform 1 0 4816 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_37
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_47
timestamp 1698431365
transform 1 0 6608 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_51
timestamp 1698431365
transform 1 0 7056 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_55
timestamp 1698431365
transform 1 0 7504 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_100
timestamp 1698431365
transform 1 0 12544 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_104
timestamp 1698431365
transform 1 0 12992 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_107
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_115
timestamp 1698431365
transform 1 0 14224 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_119
timestamp 1698431365
transform 1 0 14672 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_132
timestamp 1698431365
transform 1 0 16128 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_168
timestamp 1698431365
transform 1 0 20160 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_172
timestamp 1698431365
transform 1 0 20608 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_174
timestamp 1698431365
transform 1 0 20832 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_177
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_179
timestamp 1698431365
transform 1 0 21392 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_190
timestamp 1698431365
transform 1 0 22624 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_198
timestamp 1698431365
transform 1 0 23520 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_202
timestamp 1698431365
transform 1 0 23968 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_232
timestamp 1698431365
transform 1 0 27328 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_236
timestamp 1698431365
transform 1 0 27776 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698431365
transform 1 0 28672 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_247
timestamp 1698431365
transform 1 0 29008 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_251
timestamp 1698431365
transform 1 0 29456 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_267
timestamp 1698431365
transform 1 0 31248 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_275
timestamp 1698431365
transform 1 0 32144 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_279
timestamp 1698431365
transform 1 0 32592 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_282
timestamp 1698431365
transform 1 0 32928 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_290
timestamp 1698431365
transform 1 0 33824 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_292
timestamp 1698431365
transform 1 0 34048 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_295
timestamp 1698431365
transform 1 0 34384 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_299
timestamp 1698431365
transform 1 0 34832 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_301
timestamp 1698431365
transform 1 0 35056 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_304
timestamp 1698431365
transform 1 0 35392 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_312
timestamp 1698431365
transform 1 0 36288 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_314
timestamp 1698431365
transform 1 0 36512 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_317
timestamp 1698431365
transform 1 0 36848 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_325
timestamp 1698431365
transform 1 0 37744 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_329
timestamp 1698431365
transform 1 0 38192 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_2
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_32
timestamp 1698431365
transform 1 0 4928 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_42
timestamp 1698431365
transform 1 0 6048 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_46
timestamp 1698431365
transform 1 0 6496 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_50
timestamp 1698431365
transform 1 0 6944 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_58
timestamp 1698431365
transform 1 0 7840 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_60
timestamp 1698431365
transform 1 0 8064 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_80
timestamp 1698431365
transform 1 0 10304 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_84
timestamp 1698431365
transform 1 0 10752 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_88
timestamp 1698431365
transform 1 0 11200 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_96
timestamp 1698431365
transform 1 0 12096 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_100
timestamp 1698431365
transform 1 0 12544 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_104
timestamp 1698431365
transform 1 0 12992 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_135
timestamp 1698431365
transform 1 0 16464 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_139
timestamp 1698431365
transform 1 0 16912 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_142
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_144
timestamp 1698431365
transform 1 0 17472 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_155
timestamp 1698431365
transform 1 0 18704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_157
timestamp 1698431365
transform 1 0 18928 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_160
timestamp 1698431365
transform 1 0 19264 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_164
timestamp 1698431365
transform 1 0 19712 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_168
timestamp 1698431365
transform 1 0 20160 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_199
timestamp 1698431365
transform 1 0 23632 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_203
timestamp 1698431365
transform 1 0 24080 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_241
timestamp 1698431365
transform 1 0 28336 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_245
timestamp 1698431365
transform 1 0 28784 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_247
timestamp 1698431365
transform 1 0 29008 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_256
timestamp 1698431365
transform 1 0 30016 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_272
timestamp 1698431365
transform 1 0 31808 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_282
timestamp 1698431365
transform 1 0 32928 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_286
timestamp 1698431365
transform 1 0 33376 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_290
timestamp 1698431365
transform 1 0 33824 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_294
timestamp 1698431365
transform 1 0 34272 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_312
timestamp 1698431365
transform 1 0 36288 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_328
timestamp 1698431365
transform 1 0 38080 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_330
timestamp 1698431365
transform 1 0 38304 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_2
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_18
timestamp 1698431365
transform 1 0 3360 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_26
timestamp 1698431365
transform 1 0 4256 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_30
timestamp 1698431365
transform 1 0 4704 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_32
timestamp 1698431365
transform 1 0 4928 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_45
timestamp 1698431365
transform 1 0 6384 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_61
timestamp 1698431365
transform 1 0 8176 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_69
timestamp 1698431365
transform 1 0 9072 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_72
timestamp 1698431365
transform 1 0 9408 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_79
timestamp 1698431365
transform 1 0 10192 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_95
timestamp 1698431365
transform 1 0 11984 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_97
timestamp 1698431365
transform 1 0 12208 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_107
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_114
timestamp 1698431365
transform 1 0 14112 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_130
timestamp 1698431365
transform 1 0 15904 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_141
timestamp 1698431365
transform 1 0 17136 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_149
timestamp 1698431365
transform 1 0 18032 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_158
timestamp 1698431365
transform 1 0 19040 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_160
timestamp 1698431365
transform 1 0 19264 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_166
timestamp 1698431365
transform 1 0 19936 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_168
timestamp 1698431365
transform 1 0 20160 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_177
timestamp 1698431365
transform 1 0 21168 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_187
timestamp 1698431365
transform 1 0 22288 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_203
timestamp 1698431365
transform 1 0 24080 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_211
timestamp 1698431365
transform 1 0 24976 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_223
timestamp 1698431365
transform 1 0 26320 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_231
timestamp 1698431365
transform 1 0 27216 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_239
timestamp 1698431365
transform 1 0 28112 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_243
timestamp 1698431365
transform 1 0 28560 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_247
timestamp 1698431365
transform 1 0 29008 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_251
timestamp 1698431365
transform 1 0 29456 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_310
timestamp 1698431365
transform 1 0 36064 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_314
timestamp 1698431365
transform 1 0 36512 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_317
timestamp 1698431365
transform 1 0 36848 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_325
timestamp 1698431365
transform 1 0 37744 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_2
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_10
timestamp 1698431365
transform 1 0 2464 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_14
timestamp 1698431365
transform 1 0 2912 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_28
timestamp 1698431365
transform 1 0 4480 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_60
timestamp 1698431365
transform 1 0 8064 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_68
timestamp 1698431365
transform 1 0 8960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_101
timestamp 1698431365
transform 1 0 12656 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_111
timestamp 1698431365
transform 1 0 13776 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_115
timestamp 1698431365
transform 1 0 14224 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_131
timestamp 1698431365
transform 1 0 16016 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_139
timestamp 1698431365
transform 1 0 16912 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_142
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_174
timestamp 1698431365
transform 1 0 20832 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_176
timestamp 1698431365
transform 1 0 21056 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_206
timestamp 1698431365
transform 1 0 24416 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_212
timestamp 1698431365
transform 1 0 25088 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_218
timestamp 1698431365
transform 1 0 25760 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_226
timestamp 1698431365
transform 1 0 26656 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_279
timestamp 1698431365
transform 1 0 32592 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_288
timestamp 1698431365
transform 1 0 33600 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_296
timestamp 1698431365
transform 1 0 34496 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_328
timestamp 1698431365
transform 1 0 38080 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_330
timestamp 1698431365
transform 1 0 38304 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_2
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_18
timestamp 1698431365
transform 1 0 3360 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_26
timestamp 1698431365
transform 1 0 4256 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698431365
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_45
timestamp 1698431365
transform 1 0 6384 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_49
timestamp 1698431365
transform 1 0 6832 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_81
timestamp 1698431365
transform 1 0 10416 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_97
timestamp 1698431365
transform 1 0 12208 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_103
timestamp 1698431365
transform 1 0 12880 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_107
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_139
timestamp 1698431365
transform 1 0 16912 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_142
timestamp 1698431365
transform 1 0 17248 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_174
timestamp 1698431365
transform 1 0 20832 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_177
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_181
timestamp 1698431365
transform 1 0 21616 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_183
timestamp 1698431365
transform 1 0 21840 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_216
timestamp 1698431365
transform 1 0 25536 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_234
timestamp 1698431365
transform 1 0 27552 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_238
timestamp 1698431365
transform 1 0 28000 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_242
timestamp 1698431365
transform 1 0 28448 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698431365
transform 1 0 28672 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_247
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_255
timestamp 1698431365
transform 1 0 29904 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_259
timestamp 1698431365
transform 1 0 30352 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_263
timestamp 1698431365
transform 1 0 30800 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_267
timestamp 1698431365
transform 1 0 31248 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_271
timestamp 1698431365
transform 1 0 31696 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_303
timestamp 1698431365
transform 1 0 35280 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_312
timestamp 1698431365
transform 1 0 36288 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_314
timestamp 1698431365
transform 1 0 36512 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_2
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_18
timestamp 1698431365
transform 1 0 3360 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_26
timestamp 1698431365
transform 1 0 4256 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_38
timestamp 1698431365
transform 1 0 5600 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_54
timestamp 1698431365
transform 1 0 7392 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_64
timestamp 1698431365
transform 1 0 8512 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_68
timestamp 1698431365
transform 1 0 8960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_72
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_104
timestamp 1698431365
transform 1 0 12992 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_112
timestamp 1698431365
transform 1 0 13888 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_116
timestamp 1698431365
transform 1 0 14336 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_124
timestamp 1698431365
transform 1 0 15232 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_136
timestamp 1698431365
transform 1 0 16576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_150
timestamp 1698431365
transform 1 0 18144 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_166
timestamp 1698431365
transform 1 0 19936 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_174
timestamp 1698431365
transform 1 0 20832 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_178
timestamp 1698431365
transform 1 0 21280 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_180
timestamp 1698431365
transform 1 0 21504 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_194
timestamp 1698431365
transform 1 0 23072 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_198
timestamp 1698431365
transform 1 0 23520 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_202
timestamp 1698431365
transform 1 0 23968 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_206
timestamp 1698431365
transform 1 0 24416 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_212
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_221
timestamp 1698431365
transform 1 0 26096 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_225
timestamp 1698431365
transform 1 0 26544 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_257
timestamp 1698431365
transform 1 0 30128 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_265
timestamp 1698431365
transform 1 0 31024 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_269
timestamp 1698431365
transform 1 0 31472 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_272
timestamp 1698431365
transform 1 0 31808 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698431365
transform 1 0 32256 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_282
timestamp 1698431365
transform 1 0 32928 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_298
timestamp 1698431365
transform 1 0 34720 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_2
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_32
timestamp 1698431365
transform 1 0 4928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698431365
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_37
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_41
timestamp 1698431365
transform 1 0 5936 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_72
timestamp 1698431365
transform 1 0 9408 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_76
timestamp 1698431365
transform 1 0 9856 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_92
timestamp 1698431365
transform 1 0 11648 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_100
timestamp 1698431365
transform 1 0 12544 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_104
timestamp 1698431365
transform 1 0 12992 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_136
timestamp 1698431365
transform 1 0 16576 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_167
timestamp 1698431365
transform 1 0 20048 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698431365
transform 1 0 20496 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_177
timestamp 1698431365
transform 1 0 21168 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_193
timestamp 1698431365
transform 1 0 22960 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_201
timestamp 1698431365
transform 1 0 23856 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_203
timestamp 1698431365
transform 1 0 24080 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_206
timestamp 1698431365
transform 1 0 24416 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_210
timestamp 1698431365
transform 1 0 24864 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_212
timestamp 1698431365
transform 1 0 25088 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_226
timestamp 1698431365
transform 1 0 26656 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_230
timestamp 1698431365
transform 1 0 27104 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_238
timestamp 1698431365
transform 1 0 28000 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_242
timestamp 1698431365
transform 1 0 28448 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_244
timestamp 1698431365
transform 1 0 28672 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_247
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_257
timestamp 1698431365
transform 1 0 30128 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_261
timestamp 1698431365
transform 1 0 30576 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_270
timestamp 1698431365
transform 1 0 31584 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_281
timestamp 1698431365
transform 1 0 32816 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_297
timestamp 1698431365
transform 1 0 34608 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_323
timestamp 1698431365
transform 1 0 37520 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_327
timestamp 1698431365
transform 1 0 37968 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_2
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_18
timestamp 1698431365
transform 1 0 3360 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_26
timestamp 1698431365
transform 1 0 4256 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_28
timestamp 1698431365
transform 1 0 4480 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_31
timestamp 1698431365
transform 1 0 4816 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_39
timestamp 1698431365
transform 1 0 5712 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_80
timestamp 1698431365
transform 1 0 10304 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_84
timestamp 1698431365
transform 1 0 10752 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_100
timestamp 1698431365
transform 1 0 12544 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_104
timestamp 1698431365
transform 1 0 12992 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_107
timestamp 1698431365
transform 1 0 13328 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_111
timestamp 1698431365
transform 1 0 13776 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_127
timestamp 1698431365
transform 1 0 15568 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_131
timestamp 1698431365
transform 1 0 16016 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_133
timestamp 1698431365
transform 1 0 16240 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_151
timestamp 1698431365
transform 1 0 18256 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_155
timestamp 1698431365
transform 1 0 18704 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_163
timestamp 1698431365
transform 1 0 19600 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_169
timestamp 1698431365
transform 1 0 20272 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_173
timestamp 1698431365
transform 1 0 20720 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_177
timestamp 1698431365
transform 1 0 21168 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_208
timestamp 1698431365
transform 1 0 24640 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_212
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_219
timestamp 1698431365
transform 1 0 25872 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_221
timestamp 1698431365
transform 1 0 26096 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_229
timestamp 1698431365
transform 1 0 26992 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_260
timestamp 1698431365
transform 1 0 30464 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_264
timestamp 1698431365
transform 1 0 30912 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_268
timestamp 1698431365
transform 1 0 31360 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_271
timestamp 1698431365
transform 1 0 31696 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_282
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_314
timestamp 1698431365
transform 1 0 36512 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_320
timestamp 1698431365
transform 1 0 37184 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_328
timestamp 1698431365
transform 1 0 38080 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_330
timestamp 1698431365
transform 1 0 38304 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_2
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_10
timestamp 1698431365
transform 1 0 2464 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_20
timestamp 1698431365
transform 1 0 3584 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_29
timestamp 1698431365
transform 1 0 4592 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_33
timestamp 1698431365
transform 1 0 5040 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_37
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_41
timestamp 1698431365
transform 1 0 5936 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_51
timestamp 1698431365
transform 1 0 7056 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_55
timestamp 1698431365
transform 1 0 7504 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_57
timestamp 1698431365
transform 1 0 7728 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_64
timestamp 1698431365
transform 1 0 8512 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_68
timestamp 1698431365
transform 1 0 8960 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_72
timestamp 1698431365
transform 1 0 9408 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_115
timestamp 1698431365
transform 1 0 14224 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_131
timestamp 1698431365
transform 1 0 16016 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_139
timestamp 1698431365
transform 1 0 16912 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_142
timestamp 1698431365
transform 1 0 17248 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_150
timestamp 1698431365
transform 1 0 18144 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_152
timestamp 1698431365
transform 1 0 18368 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_172
timestamp 1698431365
transform 1 0 20608 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_174
timestamp 1698431365
transform 1 0 20832 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_177
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_193
timestamp 1698431365
transform 1 0 22960 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_244
timestamp 1698431365
transform 1 0 28672 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_247
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_251
timestamp 1698431365
transform 1 0 29456 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_255
timestamp 1698431365
transform 1 0 29904 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_266
timestamp 1698431365
transform 1 0 31136 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_270
timestamp 1698431365
transform 1 0 31584 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_279
timestamp 1698431365
transform 1 0 32592 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_283
timestamp 1698431365
transform 1 0 33040 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_317
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_325
timestamp 1698431365
transform 1 0 37744 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_39
timestamp 1698431365
transform 1 0 5712 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_47
timestamp 1698431365
transform 1 0 6608 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_53
timestamp 1698431365
transform 1 0 7280 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_69
timestamp 1698431365
transform 1 0 9072 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_72
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_86
timestamp 1698431365
transform 1 0 10976 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_117
timestamp 1698431365
transform 1 0 14448 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_121
timestamp 1698431365
transform 1 0 14896 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_123
timestamp 1698431365
transform 1 0 15120 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_142
timestamp 1698431365
transform 1 0 17248 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_146
timestamp 1698431365
transform 1 0 17696 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_150
timestamp 1698431365
transform 1 0 18144 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_180
timestamp 1698431365
transform 1 0 21504 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_184
timestamp 1698431365
transform 1 0 21952 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_186
timestamp 1698431365
transform 1 0 22176 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_193
timestamp 1698431365
transform 1 0 22960 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_207
timestamp 1698431365
transform 1 0 24528 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_209
timestamp 1698431365
transform 1 0 24752 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_212
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_216
timestamp 1698431365
transform 1 0 25536 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_220
timestamp 1698431365
transform 1 0 25984 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_224
timestamp 1698431365
transform 1 0 26432 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_241
timestamp 1698431365
transform 1 0 28336 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_249
timestamp 1698431365
transform 1 0 29232 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_290
timestamp 1698431365
transform 1 0 33824 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_298
timestamp 1698431365
transform 1 0 34720 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_2
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_24
timestamp 1698431365
transform 1 0 4032 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_28
timestamp 1698431365
transform 1 0 4480 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_31
timestamp 1698431365
transform 1 0 4816 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_37
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_69
timestamp 1698431365
transform 1 0 9072 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_77
timestamp 1698431365
transform 1 0 9968 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_81
timestamp 1698431365
transform 1 0 10416 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_88
timestamp 1698431365
transform 1 0 11200 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_96
timestamp 1698431365
transform 1 0 12096 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_98
timestamp 1698431365
transform 1 0 12320 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_107
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_123
timestamp 1698431365
transform 1 0 15120 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_127
timestamp 1698431365
transform 1 0 15568 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_172
timestamp 1698431365
transform 1 0 20608 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_174
timestamp 1698431365
transform 1 0 20832 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_177
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_193
timestamp 1698431365
transform 1 0 22960 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_197
timestamp 1698431365
transform 1 0 23408 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_201
timestamp 1698431365
transform 1 0 23856 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_208
timestamp 1698431365
transform 1 0 24640 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_224
timestamp 1698431365
transform 1 0 26432 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_230
timestamp 1698431365
transform 1 0 27104 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_238
timestamp 1698431365
transform 1 0 28000 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_242
timestamp 1698431365
transform 1 0 28448 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_244
timestamp 1698431365
transform 1 0 28672 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_247
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_251
timestamp 1698431365
transform 1 0 29456 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_253
timestamp 1698431365
transform 1 0 29680 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_284
timestamp 1698431365
transform 1 0 33152 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_300
timestamp 1698431365
transform 1 0 34944 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_308
timestamp 1698431365
transform 1 0 35840 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_312
timestamp 1698431365
transform 1 0 36288 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_314
timestamp 1698431365
transform 1 0 36512 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_317
timestamp 1698431365
transform 1 0 36848 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_325
timestamp 1698431365
transform 1 0 37744 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_329
timestamp 1698431365
transform 1 0 38192 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_2
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_6
timestamp 1698431365
transform 1 0 2016 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_37
timestamp 1698431365
transform 1 0 5488 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_41
timestamp 1698431365
transform 1 0 5936 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_49
timestamp 1698431365
transform 1 0 6832 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_53
timestamp 1698431365
transform 1 0 7280 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_61
timestamp 1698431365
transform 1 0 8176 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_65
timestamp 1698431365
transform 1 0 8624 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_67
timestamp 1698431365
transform 1 0 8848 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_72
timestamp 1698431365
transform 1 0 9408 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_74
timestamp 1698431365
transform 1 0 9632 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_83
timestamp 1698431365
transform 1 0 10640 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_115
timestamp 1698431365
transform 1 0 14224 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_131
timestamp 1698431365
transform 1 0 16016 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_138
timestamp 1698431365
transform 1 0 16800 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_142
timestamp 1698431365
transform 1 0 17248 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_160
timestamp 1698431365
transform 1 0 19264 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_169
timestamp 1698431365
transform 1 0 20272 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_185
timestamp 1698431365
transform 1 0 22064 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_189
timestamp 1698431365
transform 1 0 22512 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_191
timestamp 1698431365
transform 1 0 22736 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_202
timestamp 1698431365
transform 1 0 23968 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698431365
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_212
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_244
timestamp 1698431365
transform 1 0 28672 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_262
timestamp 1698431365
transform 1 0 30688 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_266
timestamp 1698431365
transform 1 0 31136 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_269
timestamp 1698431365
transform 1 0 31472 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_275
timestamp 1698431365
transform 1 0 32144 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_279
timestamp 1698431365
transform 1 0 32592 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_311
timestamp 1698431365
transform 1 0 36176 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_315
timestamp 1698431365
transform 1 0 36624 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698431365
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_37
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_45
timestamp 1698431365
transform 1 0 6384 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_49
timestamp 1698431365
transform 1 0 6832 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_80
timestamp 1698431365
transform 1 0 10304 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_84
timestamp 1698431365
transform 1 0 10752 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_100
timestamp 1698431365
transform 1 0 12544 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_104
timestamp 1698431365
transform 1 0 12992 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_107
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_123
timestamp 1698431365
transform 1 0 15120 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_134
timestamp 1698431365
transform 1 0 16352 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_142
timestamp 1698431365
transform 1 0 17248 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_146
timestamp 1698431365
transform 1 0 17696 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_162
timestamp 1698431365
transform 1 0 19488 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_170
timestamp 1698431365
transform 1 0 20384 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_174
timestamp 1698431365
transform 1 0 20832 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_206
timestamp 1698431365
transform 1 0 24416 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_210
timestamp 1698431365
transform 1 0 24864 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_214
timestamp 1698431365
transform 1 0 25312 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_247
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_251
timestamp 1698431365
transform 1 0 29456 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_283
timestamp 1698431365
transform 1 0 33040 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_299
timestamp 1698431365
transform 1 0 34832 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_313
timestamp 1698431365
transform 1 0 36400 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_323
timestamp 1698431365
transform 1 0 37520 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_327
timestamp 1698431365
transform 1 0 37968 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_2
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_18
timestamp 1698431365
transform 1 0 3360 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_20
timestamp 1698431365
transform 1 0 3584 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_58
timestamp 1698431365
transform 1 0 7840 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_62
timestamp 1698431365
transform 1 0 8288 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_72
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_88
timestamp 1698431365
transform 1 0 11200 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_121
timestamp 1698431365
transform 1 0 14896 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_125
timestamp 1698431365
transform 1 0 15344 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_133
timestamp 1698431365
transform 1 0 16240 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_137
timestamp 1698431365
transform 1 0 16688 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_142
timestamp 1698431365
transform 1 0 17248 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_154
timestamp 1698431365
transform 1 0 18592 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_170
timestamp 1698431365
transform 1 0 20384 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_174
timestamp 1698431365
transform 1 0 20832 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_181
timestamp 1698431365
transform 1 0 21616 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_197
timestamp 1698431365
transform 1 0 23408 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_205
timestamp 1698431365
transform 1 0 24304 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_209
timestamp 1698431365
transform 1 0 24752 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_212
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_220
timestamp 1698431365
transform 1 0 25984 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_224
timestamp 1698431365
transform 1 0 26432 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_255
timestamp 1698431365
transform 1 0 29904 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_259
timestamp 1698431365
transform 1 0 30352 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_275
timestamp 1698431365
transform 1 0 32144 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_279
timestamp 1698431365
transform 1 0 32592 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_288
timestamp 1698431365
transform 1 0 33600 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_296
timestamp 1698431365
transform 1 0 34496 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_300
timestamp 1698431365
transform 1 0 34944 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_2
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_18
timestamp 1698431365
transform 1 0 3360 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_26
timestamp 1698431365
transform 1 0 4256 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_30
timestamp 1698431365
transform 1 0 4704 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_33
timestamp 1698431365
transform 1 0 5040 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_37
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_39
timestamp 1698431365
transform 1 0 5712 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_48
timestamp 1698431365
transform 1 0 6720 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_52
timestamp 1698431365
transform 1 0 7168 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_56
timestamp 1698431365
transform 1 0 7616 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_88
timestamp 1698431365
transform 1 0 11200 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_96
timestamp 1698431365
transform 1 0 12096 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_104
timestamp 1698431365
transform 1 0 12992 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_107
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_115
timestamp 1698431365
transform 1 0 14224 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_145
timestamp 1698431365
transform 1 0 17584 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_185
timestamp 1698431365
transform 1 0 22064 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_201
timestamp 1698431365
transform 1 0 23856 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_205
timestamp 1698431365
transform 1 0 24304 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_221
timestamp 1698431365
transform 1 0 26096 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_224
timestamp 1698431365
transform 1 0 26432 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_240
timestamp 1698431365
transform 1 0 28224 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_244
timestamp 1698431365
transform 1 0 28672 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_251
timestamp 1698431365
transform 1 0 29456 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_259
timestamp 1698431365
transform 1 0 30352 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_263
timestamp 1698431365
transform 1 0 30800 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_280
timestamp 1698431365
transform 1 0 32704 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_282
timestamp 1698431365
transform 1 0 32928 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_294
timestamp 1698431365
transform 1 0 34272 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_298
timestamp 1698431365
transform 1 0 34720 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_310
timestamp 1698431365
transform 1 0 36064 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_314
timestamp 1698431365
transform 1 0 36512 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_323
timestamp 1698431365
transform 1 0 37520 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_37
timestamp 1698431365
transform 1 0 5488 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_39
timestamp 1698431365
transform 1 0 5712 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_51
timestamp 1698431365
transform 1 0 7056 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_55
timestamp 1698431365
transform 1 0 7504 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_59
timestamp 1698431365
transform 1 0 7952 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_67
timestamp 1698431365
transform 1 0 8848 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_69
timestamp 1698431365
transform 1 0 9072 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_72
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_78
timestamp 1698431365
transform 1 0 10080 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_94
timestamp 1698431365
transform 1 0 11872 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_96
timestamp 1698431365
transform 1 0 12096 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_107
timestamp 1698431365
transform 1 0 13328 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_115
timestamp 1698431365
transform 1 0 14224 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_119
timestamp 1698431365
transform 1 0 14672 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_127
timestamp 1698431365
transform 1 0 15568 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_135
timestamp 1698431365
transform 1 0 16464 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_139
timestamp 1698431365
transform 1 0 16912 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_151
timestamp 1698431365
transform 1 0 18256 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_168
timestamp 1698431365
transform 1 0 20160 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_172
timestamp 1698431365
transform 1 0 20608 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_174
timestamp 1698431365
transform 1 0 20832 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_177
timestamp 1698431365
transform 1 0 21168 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_209
timestamp 1698431365
transform 1 0 24752 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_212
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_228
timestamp 1698431365
transform 1 0 26880 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_274
timestamp 1698431365
transform 1 0 32032 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_278
timestamp 1698431365
transform 1 0 32480 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_282
timestamp 1698431365
transform 1 0 32928 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_284
timestamp 1698431365
transform 1 0 33152 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_307
timestamp 1698431365
transform 1 0 35728 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_323
timestamp 1698431365
transform 1 0 37520 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_2
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_10
timestamp 1698431365
transform 1 0 2464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_12
timestamp 1698431365
transform 1 0 2688 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_19
timestamp 1698431365
transform 1 0 3472 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_29
timestamp 1698431365
transform 1 0 4592 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_33
timestamp 1698431365
transform 1 0 5040 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_37
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_107
timestamp 1698431365
transform 1 0 13328 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_111
timestamp 1698431365
transform 1 0 13776 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_127
timestamp 1698431365
transform 1 0 15568 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_131
timestamp 1698431365
transform 1 0 16016 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_139
timestamp 1698431365
transform 1 0 16912 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_143
timestamp 1698431365
transform 1 0 17360 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_145
timestamp 1698431365
transform 1 0 17584 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_157
timestamp 1698431365
transform 1 0 18928 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_161
timestamp 1698431365
transform 1 0 19376 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_165
timestamp 1698431365
transform 1 0 19824 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_173
timestamp 1698431365
transform 1 0 20720 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_177
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_214
timestamp 1698431365
transform 1 0 25312 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_218
timestamp 1698431365
transform 1 0 25760 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_234
timestamp 1698431365
transform 1 0 27552 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_238
timestamp 1698431365
transform 1 0 28000 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_240
timestamp 1698431365
transform 1 0 28224 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_247
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_255
timestamp 1698431365
transform 1 0 29904 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_257
timestamp 1698431365
transform 1 0 30128 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_260
timestamp 1698431365
transform 1 0 30464 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_264
timestamp 1698431365
transform 1 0 30912 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_301
timestamp 1698431365
transform 1 0 35056 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_312
timestamp 1698431365
transform 1 0 36288 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_314
timestamp 1698431365
transform 1 0 36512 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_317
timestamp 1698431365
transform 1 0 36848 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_325
timestamp 1698431365
transform 1 0 37744 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_329
timestamp 1698431365
transform 1 0 38192 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_2
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_18
timestamp 1698431365
transform 1 0 3360 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_35
timestamp 1698431365
transform 1 0 5264 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_39
timestamp 1698431365
transform 1 0 5712 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_55
timestamp 1698431365
transform 1 0 7504 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_63
timestamp 1698431365
transform 1 0 8400 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_67
timestamp 1698431365
transform 1 0 8848 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_69
timestamp 1698431365
transform 1 0 9072 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_81
timestamp 1698431365
transform 1 0 10416 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_85
timestamp 1698431365
transform 1 0 10864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_89
timestamp 1698431365
transform 1 0 11312 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_93
timestamp 1698431365
transform 1 0 11760 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_123
timestamp 1698431365
transform 1 0 15120 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_134
timestamp 1698431365
transform 1 0 16352 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_138
timestamp 1698431365
transform 1 0 16800 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_153
timestamp 1698431365
transform 1 0 18480 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_157
timestamp 1698431365
transform 1 0 18928 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_172
timestamp 1698431365
transform 1 0 20608 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_176
timestamp 1698431365
transform 1 0 21056 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_192
timestamp 1698431365
transform 1 0 22848 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_194
timestamp 1698431365
transform 1 0 23072 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_197
timestamp 1698431365
transform 1 0 23408 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_205
timestamp 1698431365
transform 1 0 24304 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698431365
transform 1 0 24752 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_212
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_220
timestamp 1698431365
transform 1 0 25984 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_224
timestamp 1698431365
transform 1 0 26432 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_269
timestamp 1698431365
transform 1 0 31472 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_279
timestamp 1698431365
transform 1 0 32592 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_282
timestamp 1698431365
transform 1 0 32928 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_286
timestamp 1698431365
transform 1 0 33376 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_294
timestamp 1698431365
transform 1 0 34272 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_298
timestamp 1698431365
transform 1 0 34720 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_300
timestamp 1698431365
transform 1 0 34944 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_303
timestamp 1698431365
transform 1 0 35280 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_307
timestamp 1698431365
transform 1 0 35728 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_309
timestamp 1698431365
transform 1 0 35952 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_320
timestamp 1698431365
transform 1 0 37184 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_328
timestamp 1698431365
transform 1 0 38080 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_330
timestamp 1698431365
transform 1 0 38304 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_2
timestamp 1698431365
transform 1 0 1568 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_18
timestamp 1698431365
transform 1 0 3360 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_26
timestamp 1698431365
transform 1 0 4256 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_30
timestamp 1698431365
transform 1 0 4704 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_32
timestamp 1698431365
transform 1 0 4928 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_46
timestamp 1698431365
transform 1 0 6496 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_50
timestamp 1698431365
transform 1 0 6944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_54
timestamp 1698431365
transform 1 0 7392 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_62
timestamp 1698431365
transform 1 0 8288 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_77
timestamp 1698431365
transform 1 0 9968 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_85
timestamp 1698431365
transform 1 0 10864 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_95
timestamp 1698431365
transform 1 0 11984 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_103
timestamp 1698431365
transform 1 0 12880 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_107
timestamp 1698431365
transform 1 0 13328 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_125
timestamp 1698431365
transform 1 0 15344 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_133
timestamp 1698431365
transform 1 0 16240 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_137
timestamp 1698431365
transform 1 0 16688 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_141
timestamp 1698431365
transform 1 0 17136 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_144
timestamp 1698431365
transform 1 0 17472 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_152
timestamp 1698431365
transform 1 0 18368 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_155
timestamp 1698431365
transform 1 0 18704 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_171
timestamp 1698431365
transform 1 0 20496 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_177
timestamp 1698431365
transform 1 0 21168 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_179
timestamp 1698431365
transform 1 0 21392 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_182
timestamp 1698431365
transform 1 0 21728 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_188
timestamp 1698431365
transform 1 0 22400 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_192
timestamp 1698431365
transform 1 0 22848 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_196
timestamp 1698431365
transform 1 0 23296 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_200
timestamp 1698431365
transform 1 0 23744 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_207
timestamp 1698431365
transform 1 0 24528 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_211
timestamp 1698431365
transform 1 0 24976 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_241
timestamp 1698431365
transform 1 0 28336 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_279
timestamp 1698431365
transform 1 0 32592 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_283
timestamp 1698431365
transform 1 0 33040 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_299
timestamp 1698431365
transform 1 0 34832 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_325
timestamp 1698431365
transform 1 0 37744 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_31
timestamp 1698431365
transform 1 0 4816 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_46
timestamp 1698431365
transform 1 0 6496 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_50
timestamp 1698431365
transform 1 0 6944 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_66
timestamp 1698431365
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_80
timestamp 1698431365
transform 1 0 10304 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_84
timestamp 1698431365
transform 1 0 10752 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_102
timestamp 1698431365
transform 1 0 12768 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_106
timestamp 1698431365
transform 1 0 13216 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_113
timestamp 1698431365
transform 1 0 14000 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_121
timestamp 1698431365
transform 1 0 14896 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_133
timestamp 1698431365
transform 1 0 16240 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_135
timestamp 1698431365
transform 1 0 16464 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_138
timestamp 1698431365
transform 1 0 16800 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_142
timestamp 1698431365
transform 1 0 17248 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_148
timestamp 1698431365
transform 1 0 17920 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_152
timestamp 1698431365
transform 1 0 18368 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_160
timestamp 1698431365
transform 1 0 19264 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_164
timestamp 1698431365
transform 1 0 19712 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_168
timestamp 1698431365
transform 1 0 20160 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_180
timestamp 1698431365
transform 1 0 21504 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_184
timestamp 1698431365
transform 1 0 21952 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_186
timestamp 1698431365
transform 1 0 22176 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_195
timestamp 1698431365
transform 1 0 23184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_199
timestamp 1698431365
transform 1 0 23632 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_203
timestamp 1698431365
transform 1 0 24080 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_207
timestamp 1698431365
transform 1 0 24528 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_209
timestamp 1698431365
transform 1 0 24752 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_212
timestamp 1698431365
transform 1 0 25088 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_216
timestamp 1698431365
transform 1 0 25536 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_220
timestamp 1698431365
transform 1 0 25984 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_244
timestamp 1698431365
transform 1 0 28672 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_248
timestamp 1698431365
transform 1 0 29120 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_264
timestamp 1698431365
transform 1 0 30912 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_268
timestamp 1698431365
transform 1 0 31360 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_272
timestamp 1698431365
transform 1 0 31808 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_282
timestamp 1698431365
transform 1 0 32928 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_298
timestamp 1698431365
transform 1 0 34720 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_2
timestamp 1698431365
transform 1 0 1568 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_10
timestamp 1698431365
transform 1 0 2464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_12
timestamp 1698431365
transform 1 0 2688 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_19
timestamp 1698431365
transform 1 0 3472 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_23
timestamp 1698431365
transform 1 0 3920 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_33
timestamp 1698431365
transform 1 0 5040 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_37
timestamp 1698431365
transform 1 0 5488 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_41
timestamp 1698431365
transform 1 0 5936 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_49
timestamp 1698431365
transform 1 0 6832 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_88
timestamp 1698431365
transform 1 0 11200 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_92
timestamp 1698431365
transform 1 0 11648 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_100
timestamp 1698431365
transform 1 0 12544 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_104
timestamp 1698431365
transform 1 0 12992 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_107
timestamp 1698431365
transform 1 0 13328 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_111
timestamp 1698431365
transform 1 0 13776 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_122
timestamp 1698431365
transform 1 0 15008 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_173
timestamp 1698431365
transform 1 0 20720 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_177
timestamp 1698431365
transform 1 0 21168 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_179
timestamp 1698431365
transform 1 0 21392 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_189
timestamp 1698431365
transform 1 0 22512 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_222
timestamp 1698431365
transform 1 0 26208 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_226
timestamp 1698431365
transform 1 0 26656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_230
timestamp 1698431365
transform 1 0 27104 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_238
timestamp 1698431365
transform 1 0 28000 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_242
timestamp 1698431365
transform 1 0 28448 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_244
timestamp 1698431365
transform 1 0 28672 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_247
timestamp 1698431365
transform 1 0 29008 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_255
timestamp 1698431365
transform 1 0 29904 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_288
timestamp 1698431365
transform 1 0 33600 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_292
timestamp 1698431365
transform 1 0 34048 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_300
timestamp 1698431365
transform 1 0 34944 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_323
timestamp 1698431365
transform 1 0 37520 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_327
timestamp 1698431365
transform 1 0 37968 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_31
timestamp 1698431365
transform 1 0 4816 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_35
timestamp 1698431365
transform 1 0 5264 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_50
timestamp 1698431365
transform 1 0 6944 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_66
timestamp 1698431365
transform 1 0 8736 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_72
timestamp 1698431365
transform 1 0 9408 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_76
timestamp 1698431365
transform 1 0 9856 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_83
timestamp 1698431365
transform 1 0 10640 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_99
timestamp 1698431365
transform 1 0 12432 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_103
timestamp 1698431365
transform 1 0 12880 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_135
timestamp 1698431365
transform 1 0 16464 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_137
timestamp 1698431365
transform 1 0 16688 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_148
timestamp 1698431365
transform 1 0 17920 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_150
timestamp 1698431365
transform 1 0 18144 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_190
timestamp 1698431365
transform 1 0 22624 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_194
timestamp 1698431365
transform 1 0 23072 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_198
timestamp 1698431365
transform 1 0 23520 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_209
timestamp 1698431365
transform 1 0 24752 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_259
timestamp 1698431365
transform 1 0 30352 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_263
timestamp 1698431365
transform 1 0 30800 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_267
timestamp 1698431365
transform 1 0 31248 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_270
timestamp 1698431365
transform 1 0 31584 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_279
timestamp 1698431365
transform 1 0 32592 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_290
timestamp 1698431365
transform 1 0 33824 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_298
timestamp 1698431365
transform 1 0 34720 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_2
timestamp 1698431365
transform 1 0 1568 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_10
timestamp 1698431365
transform 1 0 2464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_12
timestamp 1698431365
transform 1 0 2688 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_19
timestamp 1698431365
transform 1 0 3472 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_23
timestamp 1698431365
transform 1 0 3920 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_25
timestamp 1698431365
transform 1 0 4144 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_46
timestamp 1698431365
transform 1 0 6496 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_50
timestamp 1698431365
transform 1 0 6944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_54
timestamp 1698431365
transform 1 0 7392 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_86
timestamp 1698431365
transform 1 0 10976 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_94
timestamp 1698431365
transform 1 0 11872 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_98
timestamp 1698431365
transform 1 0 12320 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_101
timestamp 1698431365
transform 1 0 12656 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_107
timestamp 1698431365
transform 1 0 13328 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_109
timestamp 1698431365
transform 1 0 13552 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_162
timestamp 1698431365
transform 1 0 19488 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_164
timestamp 1698431365
transform 1 0 19712 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_167
timestamp 1698431365
transform 1 0 20048 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_171
timestamp 1698431365
transform 1 0 20496 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_177
timestamp 1698431365
transform 1 0 21168 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_179
timestamp 1698431365
transform 1 0 21392 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_194
timestamp 1698431365
transform 1 0 23072 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_247
timestamp 1698431365
transform 1 0 29008 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_251
timestamp 1698431365
transform 1 0 29456 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_257
timestamp 1698431365
transform 1 0 30128 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_287
timestamp 1698431365
transform 1 0 33488 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_291
timestamp 1698431365
transform 1 0 33936 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_293
timestamp 1698431365
transform 1 0 34160 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_314
timestamp 1698431365
transform 1 0 36512 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_2
timestamp 1698431365
transform 1 0 1568 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_18
timestamp 1698431365
transform 1 0 3360 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_30
timestamp 1698431365
transform 1 0 4704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_34
timestamp 1698431365
transform 1 0 5152 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_44
timestamp 1698431365
transform 1 0 6272 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_48
timestamp 1698431365
transform 1 0 6720 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_52
timestamp 1698431365
transform 1 0 7168 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_68
timestamp 1698431365
transform 1 0 8960 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_72
timestamp 1698431365
transform 1 0 9408 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_74
timestamp 1698431365
transform 1 0 9632 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_104
timestamp 1698431365
transform 1 0 12992 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_130
timestamp 1698431365
transform 1 0 15904 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_136
timestamp 1698431365
transform 1 0 16576 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_168
timestamp 1698431365
transform 1 0 20160 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_172
timestamp 1698431365
transform 1 0 20608 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_179
timestamp 1698431365
transform 1 0 21392 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_183
timestamp 1698431365
transform 1 0 21840 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_186
timestamp 1698431365
transform 1 0 22176 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_190
timestamp 1698431365
transform 1 0 22624 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_194
timestamp 1698431365
transform 1 0 23072 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_198
timestamp 1698431365
transform 1 0 23520 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_202
timestamp 1698431365
transform 1 0 23968 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_206
timestamp 1698431365
transform 1 0 24416 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_212
timestamp 1698431365
transform 1 0 25088 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_216
timestamp 1698431365
transform 1 0 25536 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_220
timestamp 1698431365
transform 1 0 25984 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_232
timestamp 1698431365
transform 1 0 27328 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_236
timestamp 1698431365
transform 1 0 27776 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_240
timestamp 1698431365
transform 1 0 28224 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_244
timestamp 1698431365
transform 1 0 28672 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_246
timestamp 1698431365
transform 1 0 28896 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_263
timestamp 1698431365
transform 1 0 30800 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_279
timestamp 1698431365
transform 1 0 32592 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_282
timestamp 1698431365
transform 1 0 32928 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_298
timestamp 1698431365
transform 1 0 34720 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_302
timestamp 1698431365
transform 1 0 35168 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_305
timestamp 1698431365
transform 1 0 35504 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_309
timestamp 1698431365
transform 1 0 35952 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_327
timestamp 1698431365
transform 1 0 37968 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_2
timestamp 1698431365
transform 1 0 1568 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_34
timestamp 1698431365
transform 1 0 5152 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_37
timestamp 1698431365
transform 1 0 5488 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_41
timestamp 1698431365
transform 1 0 5936 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_43
timestamp 1698431365
transform 1 0 6160 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_50
timestamp 1698431365
transform 1 0 6944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_54
timestamp 1698431365
transform 1 0 7392 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_70
timestamp 1698431365
transform 1 0 9184 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_74
timestamp 1698431365
transform 1 0 9632 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_107
timestamp 1698431365
transform 1 0 13328 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_111
timestamp 1698431365
transform 1 0 13776 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_194
timestamp 1698431365
transform 1 0 23072 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_198
timestamp 1698431365
transform 1 0 23520 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_202
timestamp 1698431365
transform 1 0 23968 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_204
timestamp 1698431365
transform 1 0 24192 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_223
timestamp 1698431365
transform 1 0 26320 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_227
timestamp 1698431365
transform 1 0 26768 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_231
timestamp 1698431365
transform 1 0 27216 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_235
timestamp 1698431365
transform 1 0 27664 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_239
timestamp 1698431365
transform 1 0 28112 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_243
timestamp 1698431365
transform 1 0 28560 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_247
timestamp 1698431365
transform 1 0 29008 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_251
timestamp 1698431365
transform 1 0 29456 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_255
timestamp 1698431365
transform 1 0 29904 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_259
timestamp 1698431365
transform 1 0 30352 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_263
timestamp 1698431365
transform 1 0 30800 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_273
timestamp 1698431365
transform 1 0 31920 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_289
timestamp 1698431365
transform 1 0 33712 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_297
timestamp 1698431365
transform 1 0 34608 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_317
timestamp 1698431365
transform 1 0 36848 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_51_2
timestamp 1698431365
transform 1 0 1568 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_34
timestamp 1698431365
transform 1 0 5152 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_36
timestamp 1698431365
transform 1 0 5376 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_54
timestamp 1698431365
transform 1 0 7392 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_58
timestamp 1698431365
transform 1 0 7840 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_62
timestamp 1698431365
transform 1 0 8288 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_80
timestamp 1698431365
transform 1 0 10304 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_87
timestamp 1698431365
transform 1 0 11088 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_91
timestamp 1698431365
transform 1 0 11536 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_95
timestamp 1698431365
transform 1 0 11984 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_107
timestamp 1698431365
transform 1 0 13328 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_115
timestamp 1698431365
transform 1 0 14224 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_119
timestamp 1698431365
transform 1 0 14672 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_121
timestamp 1698431365
transform 1 0 14896 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_124
timestamp 1698431365
transform 1 0 15232 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_128
timestamp 1698431365
transform 1 0 15680 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_132
timestamp 1698431365
transform 1 0 16128 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_136
timestamp 1698431365
transform 1 0 16576 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_142
timestamp 1698431365
transform 1 0 17248 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_191
timestamp 1698431365
transform 1 0 22736 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_204
timestamp 1698431365
transform 1 0 24192 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_208
timestamp 1698431365
transform 1 0 24640 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_219
timestamp 1698431365
transform 1 0 25872 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_234
timestamp 1698431365
transform 1 0 27552 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_238
timestamp 1698431365
transform 1 0 28000 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_242
timestamp 1698431365
transform 1 0 28448 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_244
timestamp 1698431365
transform 1 0 28672 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_258
timestamp 1698431365
transform 1 0 30240 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_262
timestamp 1698431365
transform 1 0 30688 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_274
timestamp 1698431365
transform 1 0 32032 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_278
timestamp 1698431365
transform 1 0 32480 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_282
timestamp 1698431365
transform 1 0 32928 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_290
timestamp 1698431365
transform 1 0 33824 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_294
timestamp 1698431365
transform 1 0 34272 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_301
timestamp 1698431365
transform 1 0 35056 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_2
timestamp 1698431365
transform 1 0 1568 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_18
timestamp 1698431365
transform 1 0 3360 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_26
timestamp 1698431365
transform 1 0 4256 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_30
timestamp 1698431365
transform 1 0 4704 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_32
timestamp 1698431365
transform 1 0 4928 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_83
timestamp 1698431365
transform 1 0 10640 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_87
timestamp 1698431365
transform 1 0 11088 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_91
timestamp 1698431365
transform 1 0 11536 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_95
timestamp 1698431365
transform 1 0 11984 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_103
timestamp 1698431365
transform 1 0 12880 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_107
timestamp 1698431365
transform 1 0 13328 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_117
timestamp 1698431365
transform 1 0 14448 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_171
timestamp 1698431365
transform 1 0 20496 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_243
timestamp 1698431365
transform 1 0 28560 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_247
timestamp 1698431365
transform 1 0 29008 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_249
timestamp 1698431365
transform 1 0 29232 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_266
timestamp 1698431365
transform 1 0 31136 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_270
timestamp 1698431365
transform 1 0 31584 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_274
timestamp 1698431365
transform 1 0 32032 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_278
timestamp 1698431365
transform 1 0 32480 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_311
timestamp 1698431365
transform 1 0 36176 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_323
timestamp 1698431365
transform 1 0 37520 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_327
timestamp 1698431365
transform 1 0 37968 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_2
timestamp 1698431365
transform 1 0 1568 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_35
timestamp 1698431365
transform 1 0 5264 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_39
timestamp 1698431365
transform 1 0 5712 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_72
timestamp 1698431365
transform 1 0 9408 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_76
timestamp 1698431365
transform 1 0 9856 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_80
timestamp 1698431365
transform 1 0 10304 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_117
timestamp 1698431365
transform 1 0 14448 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_142
timestamp 1698431365
transform 1 0 17248 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_206
timestamp 1698431365
transform 1 0 24416 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_212
timestamp 1698431365
transform 1 0 25088 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_214
timestamp 1698431365
transform 1 0 25312 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_244
timestamp 1698431365
transform 1 0 28672 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_248
timestamp 1698431365
transform 1 0 29120 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_250
timestamp 1698431365
transform 1 0 29344 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_282
timestamp 1698431365
transform 1 0 32928 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_286
timestamp 1698431365
transform 1 0 33376 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_294
timestamp 1698431365
transform 1 0 34272 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_53_299
timestamp 1698431365
transform 1 0 34832 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_2
timestamp 1698431365
transform 1 0 1568 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_6
timestamp 1698431365
transform 1 0 2016 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_27
timestamp 1698431365
transform 1 0 4368 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_31
timestamp 1698431365
transform 1 0 4816 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_37
timestamp 1698431365
transform 1 0 5488 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_45
timestamp 1698431365
transform 1 0 6384 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_52
timestamp 1698431365
transform 1 0 7168 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_84
timestamp 1698431365
transform 1 0 10752 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_100
timestamp 1698431365
transform 1 0 12544 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_104
timestamp 1698431365
transform 1 0 12992 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_107
timestamp 1698431365
transform 1 0 13328 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_115
timestamp 1698431365
transform 1 0 14224 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_119
timestamp 1698431365
transform 1 0 14672 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_125
timestamp 1698431365
transform 1 0 15344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_166
timestamp 1698431365
transform 1 0 19936 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_168
timestamp 1698431365
transform 1 0 20160 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_171
timestamp 1698431365
transform 1 0 20496 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_190
timestamp 1698431365
transform 1 0 22624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_240
timestamp 1698431365
transform 1 0 28224 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_244
timestamp 1698431365
transform 1 0 28672 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_247
timestamp 1698431365
transform 1 0 29008 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_251
timestamp 1698431365
transform 1 0 29456 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_255
timestamp 1698431365
transform 1 0 29904 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_271
timestamp 1698431365
transform 1 0 31696 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_275
timestamp 1698431365
transform 1 0 32144 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_279
timestamp 1698431365
transform 1 0 32592 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_283
timestamp 1698431365
transform 1 0 33040 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_317
timestamp 1698431365
transform 1 0 36848 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_325
timestamp 1698431365
transform 1 0 37744 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_329
timestamp 1698431365
transform 1 0 38192 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_31
timestamp 1698431365
transform 1 0 4816 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_35
timestamp 1698431365
transform 1 0 5264 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_51
timestamp 1698431365
transform 1 0 7056 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_55
timestamp 1698431365
transform 1 0 7504 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_66
timestamp 1698431365
transform 1 0 8736 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_72
timestamp 1698431365
transform 1 0 9408 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_80
timestamp 1698431365
transform 1 0 10304 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_84
timestamp 1698431365
transform 1 0 10752 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_96
timestamp 1698431365
transform 1 0 12096 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_100
timestamp 1698431365
transform 1 0 12544 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_108
timestamp 1698431365
transform 1 0 13440 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_114
timestamp 1698431365
transform 1 0 14112 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_118
timestamp 1698431365
transform 1 0 14560 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_207
timestamp 1698431365
transform 1 0 24528 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_209
timestamp 1698431365
transform 1 0 24752 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_261
timestamp 1698431365
transform 1 0 30576 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_265
timestamp 1698431365
transform 1 0 31024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_269
timestamp 1698431365
transform 1 0 31472 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_273
timestamp 1698431365
transform 1 0 31920 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_277
timestamp 1698431365
transform 1 0 32368 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_279
timestamp 1698431365
transform 1 0 32592 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_55_282
timestamp 1698431365
transform 1 0 32928 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_314
timestamp 1698431365
transform 1 0 36512 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_330
timestamp 1698431365
transform 1 0 38304 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_2
timestamp 1698431365
transform 1 0 1568 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_18
timestamp 1698431365
transform 1 0 3360 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_27
timestamp 1698431365
transform 1 0 4368 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_31
timestamp 1698431365
transform 1 0 4816 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_37
timestamp 1698431365
transform 1 0 5488 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_101
timestamp 1698431365
transform 1 0 12656 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_115
timestamp 1698431365
transform 1 0 14224 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_121
timestamp 1698431365
transform 1 0 14896 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_173
timestamp 1698431365
transform 1 0 20720 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_195
timestamp 1698431365
transform 1 0 23184 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_244
timestamp 1698431365
transform 1 0 28672 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_247
timestamp 1698431365
transform 1 0 29008 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_251
timestamp 1698431365
transform 1 0 29456 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_255
timestamp 1698431365
transform 1 0 29904 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_259
timestamp 1698431365
transform 1 0 30352 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_263
timestamp 1698431365
transform 1 0 30800 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_267
timestamp 1698431365
transform 1 0 31248 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_299
timestamp 1698431365
transform 1 0 34832 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_302
timestamp 1698431365
transform 1 0 35168 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_310
timestamp 1698431365
transform 1 0 36064 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_312
timestamp 1698431365
transform 1 0 36288 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_325
timestamp 1698431365
transform 1 0 37744 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_57_2
timestamp 1698431365
transform 1 0 1568 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_34
timestamp 1698431365
transform 1 0 5152 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_37
timestamp 1698431365
transform 1 0 5488 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_59
timestamp 1698431365
transform 1 0 7952 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_67
timestamp 1698431365
transform 1 0 8848 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_69
timestamp 1698431365
transform 1 0 9072 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_72
timestamp 1698431365
transform 1 0 9408 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_76
timestamp 1698431365
transform 1 0 9856 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_84
timestamp 1698431365
transform 1 0 10752 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_86
timestamp 1698431365
transform 1 0 10976 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_93
timestamp 1698431365
transform 1 0 11760 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_109
timestamp 1698431365
transform 1 0 13552 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_118
timestamp 1698431365
transform 1 0 14560 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_124
timestamp 1698431365
transform 1 0 15232 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_128
timestamp 1698431365
transform 1 0 15680 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_132
timestamp 1698431365
transform 1 0 16128 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_136
timestamp 1698431365
transform 1 0 16576 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_142
timestamp 1698431365
transform 1 0 17248 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_202
timestamp 1698431365
transform 1 0 23968 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_206
timestamp 1698431365
transform 1 0 24416 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_229
timestamp 1698431365
transform 1 0 26992 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_233
timestamp 1698431365
transform 1 0 27440 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_237
timestamp 1698431365
transform 1 0 27888 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_241
timestamp 1698431365
transform 1 0 28336 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_245
timestamp 1698431365
transform 1 0 28784 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_249
timestamp 1698431365
transform 1 0 29232 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_259
timestamp 1698431365
transform 1 0 30352 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_263
timestamp 1698431365
transform 1 0 30800 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_279
timestamp 1698431365
transform 1 0 32592 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_282
timestamp 1698431365
transform 1 0 32928 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_284
timestamp 1698431365
transform 1 0 33152 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_287
timestamp 1698431365
transform 1 0 33488 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_295
timestamp 1698431365
transform 1 0 34384 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_298
timestamp 1698431365
transform 1 0 34720 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_2
timestamp 1698431365
transform 1 0 1568 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_37
timestamp 1698431365
transform 1 0 5488 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_70
timestamp 1698431365
transform 1 0 9184 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_74
timestamp 1698431365
transform 1 0 9632 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_107
timestamp 1698431365
transform 1 0 13328 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_111
timestamp 1698431365
transform 1 0 13776 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_117
timestamp 1698431365
transform 1 0 14448 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_130
timestamp 1698431365
transform 1 0 15904 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_171
timestamp 1698431365
transform 1 0 20496 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_227
timestamp 1698431365
transform 1 0 26768 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_231
timestamp 1698431365
transform 1 0 27216 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_235
timestamp 1698431365
transform 1 0 27664 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_239
timestamp 1698431365
transform 1 0 28112 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_243
timestamp 1698431365
transform 1 0 28560 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_247
timestamp 1698431365
transform 1 0 29008 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_249
timestamp 1698431365
transform 1 0 29232 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_256
timestamp 1698431365
transform 1 0 30016 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_260
timestamp 1698431365
transform 1 0 30464 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_262
timestamp 1698431365
transform 1 0 30688 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_325
timestamp 1698431365
transform 1 0 37744 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_329
timestamp 1698431365
transform 1 0 38192 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_2
timestamp 1698431365
transform 1 0 1568 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_18
timestamp 1698431365
transform 1 0 3360 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_26
timestamp 1698431365
transform 1 0 4256 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_28
timestamp 1698431365
transform 1 0 4480 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_37
timestamp 1698431365
transform 1 0 5488 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_39
timestamp 1698431365
transform 1 0 5712 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_69
timestamp 1698431365
transform 1 0 9072 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_72
timestamp 1698431365
transform 1 0 9408 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_85
timestamp 1698431365
transform 1 0 10864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_87
timestamp 1698431365
transform 1 0 11088 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_96
timestamp 1698431365
transform 1 0 12096 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_100
timestamp 1698431365
transform 1 0 12544 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_104
timestamp 1698431365
transform 1 0 12992 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_108
timestamp 1698431365
transform 1 0 13440 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_110
timestamp 1698431365
transform 1 0 13664 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_113
timestamp 1698431365
transform 1 0 14000 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_121
timestamp 1698431365
transform 1 0 14896 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_206
timestamp 1698431365
transform 1 0 24416 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_212
timestamp 1698431365
transform 1 0 25088 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_219
timestamp 1698431365
transform 1 0 25872 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_223
timestamp 1698431365
transform 1 0 26320 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_225
timestamp 1698431365
transform 1 0 26544 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_232
timestamp 1698431365
transform 1 0 27328 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_236
timestamp 1698431365
transform 1 0 27776 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_240
timestamp 1698431365
transform 1 0 28224 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_278
timestamp 1698431365
transform 1 0 32480 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_282
timestamp 1698431365
transform 1 0 32928 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_286
timestamp 1698431365
transform 1 0 33376 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_296
timestamp 1698431365
transform 1 0 34496 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_300
timestamp 1698431365
transform 1 0 34944 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_60_2
timestamp 1698431365
transform 1 0 1568 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_34
timestamp 1698431365
transform 1 0 5152 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_37
timestamp 1698431365
transform 1 0 5488 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_45
timestamp 1698431365
transform 1 0 6384 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_90
timestamp 1698431365
transform 1 0 11424 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_94
timestamp 1698431365
transform 1 0 11872 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_98
timestamp 1698431365
transform 1 0 12320 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_101
timestamp 1698431365
transform 1 0 12656 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_118
timestamp 1698431365
transform 1 0 14560 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_122
timestamp 1698431365
transform 1 0 15008 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_135
timestamp 1698431365
transform 1 0 16464 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_137
timestamp 1698431365
transform 1 0 16688 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_238
timestamp 1698431365
transform 1 0 28000 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_242
timestamp 1698431365
transform 1 0 28448 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_244
timestamp 1698431365
transform 1 0 28672 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_247
timestamp 1698431365
transform 1 0 29008 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_251
timestamp 1698431365
transform 1 0 29456 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_264
timestamp 1698431365
transform 1 0 30912 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_268
timestamp 1698431365
transform 1 0 31360 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_299
timestamp 1698431365
transform 1 0 34832 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_309
timestamp 1698431365
transform 1 0 35952 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_313
timestamp 1698431365
transform 1 0 36400 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_323
timestamp 1698431365
transform 1 0 37520 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_327
timestamp 1698431365
transform 1 0 37968 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_31
timestamp 1698431365
transform 1 0 4816 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_35
timestamp 1698431365
transform 1 0 5264 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_51
timestamp 1698431365
transform 1 0 7056 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_59
timestamp 1698431365
transform 1 0 7952 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_63
timestamp 1698431365
transform 1 0 8400 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_67
timestamp 1698431365
transform 1 0 8848 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_69
timestamp 1698431365
transform 1 0 9072 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_72
timestamp 1698431365
transform 1 0 9408 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_76
timestamp 1698431365
transform 1 0 9856 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_84
timestamp 1698431365
transform 1 0 10752 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_88
timestamp 1698431365
transform 1 0 11200 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_137
timestamp 1698431365
transform 1 0 16688 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_139
timestamp 1698431365
transform 1 0 16912 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_142
timestamp 1698431365
transform 1 0 17248 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_159
timestamp 1698431365
transform 1 0 19152 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_163
timestamp 1698431365
transform 1 0 19600 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_209
timestamp 1698431365
transform 1 0 24752 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_226
timestamp 1698431365
transform 1 0 26656 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_256
timestamp 1698431365
transform 1 0 30016 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_260
timestamp 1698431365
transform 1 0 30464 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_264
timestamp 1698431365
transform 1 0 30912 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_282
timestamp 1698431365
transform 1 0 32928 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_286
timestamp 1698431365
transform 1 0 33376 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_293
timestamp 1698431365
transform 1 0 34160 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_295
timestamp 1698431365
transform 1 0 34384 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_304
timestamp 1698431365
transform 1 0 35392 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_308
timestamp 1698431365
transform 1 0 35840 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_324
timestamp 1698431365
transform 1 0 37632 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_328
timestamp 1698431365
transform 1 0 38080 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_330
timestamp 1698431365
transform 1 0 38304 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_62_2
timestamp 1698431365
transform 1 0 1568 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_34
timestamp 1698431365
transform 1 0 5152 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_37
timestamp 1698431365
transform 1 0 5488 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_41
timestamp 1698431365
transform 1 0 5936 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_51
timestamp 1698431365
transform 1 0 7056 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_55
timestamp 1698431365
transform 1 0 7504 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_63
timestamp 1698431365
transform 1 0 8400 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_87
timestamp 1698431365
transform 1 0 11088 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_91
timestamp 1698431365
transform 1 0 11536 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_99
timestamp 1698431365
transform 1 0 12432 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_103
timestamp 1698431365
transform 1 0 12880 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_107
timestamp 1698431365
transform 1 0 13328 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_115
timestamp 1698431365
transform 1 0 14224 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_121
timestamp 1698431365
transform 1 0 14896 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_123
timestamp 1698431365
transform 1 0 15120 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_131
timestamp 1698431365
transform 1 0 16016 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_135
timestamp 1698431365
transform 1 0 16464 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_195
timestamp 1698431365
transform 1 0 23184 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_199
timestamp 1698431365
transform 1 0 23632 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_229
timestamp 1698431365
transform 1 0 26992 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_233
timestamp 1698431365
transform 1 0 27440 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_237
timestamp 1698431365
transform 1 0 27888 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_62_247
timestamp 1698431365
transform 1 0 29008 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_279
timestamp 1698431365
transform 1 0 32592 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_295
timestamp 1698431365
transform 1 0 34384 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_297
timestamp 1698431365
transform 1 0 34608 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_300
timestamp 1698431365
transform 1 0 34944 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_304
timestamp 1698431365
transform 1 0 35392 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_312
timestamp 1698431365
transform 1 0 36288 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_314
timestamp 1698431365
transform 1 0 36512 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_317
timestamp 1698431365
transform 1 0 36848 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_325
timestamp 1698431365
transform 1 0 37744 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_329
timestamp 1698431365
transform 1 0 38192 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_2
timestamp 1698431365
transform 1 0 1568 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_10
timestamp 1698431365
transform 1 0 2464 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_14
timestamp 1698431365
transform 1 0 2912 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_27
timestamp 1698431365
transform 1 0 4368 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_31
timestamp 1698431365
transform 1 0 4816 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_63_35
timestamp 1698431365
transform 1 0 5264 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_67
timestamp 1698431365
transform 1 0 8848 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_69
timestamp 1698431365
transform 1 0 9072 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_72
timestamp 1698431365
transform 1 0 9408 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_80
timestamp 1698431365
transform 1 0 10304 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_82
timestamp 1698431365
transform 1 0 10528 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_63_85
timestamp 1698431365
transform 1 0 10864 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_117
timestamp 1698431365
transform 1 0 14448 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_125
timestamp 1698431365
transform 1 0 15344 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_129
timestamp 1698431365
transform 1 0 15792 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_132
timestamp 1698431365
transform 1 0 16128 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_136
timestamp 1698431365
transform 1 0 16576 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_142
timestamp 1698431365
transform 1 0 17248 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_212
timestamp 1698431365
transform 1 0 25088 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_216
timestamp 1698431365
transform 1 0 25536 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_63_220
timestamp 1698431365
transform 1 0 25984 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_252
timestamp 1698431365
transform 1 0 29568 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_264
timestamp 1698431365
transform 1 0 30912 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_268
timestamp 1698431365
transform 1 0 31360 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_276
timestamp 1698431365
transform 1 0 32256 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_63_282
timestamp 1698431365
transform 1 0 32928 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_314
timestamp 1698431365
transform 1 0 36512 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_317
timestamp 1698431365
transform 1 0 36848 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_325
timestamp 1698431365
transform 1 0 37744 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_329
timestamp 1698431365
transform 1 0 38192 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_2
timestamp 1698431365
transform 1 0 1568 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_33
timestamp 1698431365
transform 1 0 5040 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_37
timestamp 1698431365
transform 1 0 5488 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_41
timestamp 1698431365
transform 1 0 5936 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_44
timestamp 1698431365
transform 1 0 6272 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_76
timestamp 1698431365
transform 1 0 9856 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_92
timestamp 1698431365
transform 1 0 11648 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_100
timestamp 1698431365
transform 1 0 12544 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_104
timestamp 1698431365
transform 1 0 12992 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_107
timestamp 1698431365
transform 1 0 13328 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_115
timestamp 1698431365
transform 1 0 14224 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_121
timestamp 1698431365
transform 1 0 14896 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_123
timestamp 1698431365
transform 1 0 15120 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_135
timestamp 1698431365
transform 1 0 16464 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_137
timestamp 1698431365
transform 1 0 16688 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_140
timestamp 1698431365
transform 1 0 17024 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_144
timestamp 1698431365
transform 1 0 17472 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_164
timestamp 1698431365
transform 1 0 19712 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_206
timestamp 1698431365
transform 1 0 24416 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_210
timestamp 1698431365
transform 1 0 24864 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_214
timestamp 1698431365
transform 1 0 25312 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_230
timestamp 1698431365
transform 1 0 27104 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_238
timestamp 1698431365
transform 1 0 28000 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_242
timestamp 1698431365
transform 1 0 28448 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_244
timestamp 1698431365
transform 1 0 28672 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_247
timestamp 1698431365
transform 1 0 29008 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_254
timestamp 1698431365
transform 1 0 29792 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_258
timestamp 1698431365
transform 1 0 30240 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_288
timestamp 1698431365
transform 1 0 33600 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_292
timestamp 1698431365
transform 1 0 34048 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_300
timestamp 1698431365
transform 1 0 34944 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_310
timestamp 1698431365
transform 1 0 36064 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_314
timestamp 1698431365
transform 1 0 36512 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_325
timestamp 1698431365
transform 1 0 37744 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_40
timestamp 1698431365
transform 1 0 5824 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_42
timestamp 1698431365
transform 1 0 6048 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_51
timestamp 1698431365
transform 1 0 7056 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_63
timestamp 1698431365
transform 1 0 8400 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_67
timestamp 1698431365
transform 1 0 8848 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_69
timestamp 1698431365
transform 1 0 9072 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_72
timestamp 1698431365
transform 1 0 9408 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_88
timestamp 1698431365
transform 1 0 11200 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_100
timestamp 1698431365
transform 1 0 12544 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_102
timestamp 1698431365
transform 1 0 12768 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_138
timestamp 1698431365
transform 1 0 16800 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_148
timestamp 1698431365
transform 1 0 17920 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_152
timestamp 1698431365
transform 1 0 18368 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_163
timestamp 1698431365
transform 1 0 19600 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_165
timestamp 1698431365
transform 1 0 19824 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_195
timestamp 1698431365
transform 1 0 23184 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_199
timestamp 1698431365
transform 1 0 23632 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_203
timestamp 1698431365
transform 1 0 24080 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_207
timestamp 1698431365
transform 1 0 24528 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_209
timestamp 1698431365
transform 1 0 24752 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_241
timestamp 1698431365
transform 1 0 28336 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_245
timestamp 1698431365
transform 1 0 28784 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_261
timestamp 1698431365
transform 1 0 30576 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_268
timestamp 1698431365
transform 1 0 31360 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_278
timestamp 1698431365
transform 1 0 32480 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_290
timestamp 1698431365
transform 1 0 33824 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_294
timestamp 1698431365
transform 1 0 34272 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_298
timestamp 1698431365
transform 1 0 34720 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_2
timestamp 1698431365
transform 1 0 1568 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_10
timestamp 1698431365
transform 1 0 2464 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_14
timestamp 1698431365
transform 1 0 2912 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_16
timestamp 1698431365
transform 1 0 3136 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_23
timestamp 1698431365
transform 1 0 3920 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_33
timestamp 1698431365
transform 1 0 5040 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_37
timestamp 1698431365
transform 1 0 5488 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_39
timestamp 1698431365
transform 1 0 5712 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_42
timestamp 1698431365
transform 1 0 6048 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_66
timestamp 1698431365
transform 1 0 8736 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_70
timestamp 1698431365
transform 1 0 9184 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_74
timestamp 1698431365
transform 1 0 9632 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_113
timestamp 1698431365
transform 1 0 14000 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_117
timestamp 1698431365
transform 1 0 14448 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_125
timestamp 1698431365
transform 1 0 15344 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_131
timestamp 1698431365
transform 1 0 16016 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_172
timestamp 1698431365
transform 1 0 20608 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_174
timestamp 1698431365
transform 1 0 20832 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_190
timestamp 1698431365
transform 1 0 22624 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_194
timestamp 1698431365
transform 1 0 23072 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_198
timestamp 1698431365
transform 1 0 23520 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_214
timestamp 1698431365
transform 1 0 25312 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_222
timestamp 1698431365
transform 1 0 26208 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_224
timestamp 1698431365
transform 1 0 26432 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_231
timestamp 1698431365
transform 1 0 27216 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_239
timestamp 1698431365
transform 1 0 28112 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_243
timestamp 1698431365
transform 1 0 28560 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_305
timestamp 1698431365
transform 1 0 35504 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_307
timestamp 1698431365
transform 1 0 35728 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_314
timestamp 1698431365
transform 1 0 36512 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_323
timestamp 1698431365
transform 1 0 37520 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_327
timestamp 1698431365
transform 1 0 37968 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_2
timestamp 1698431365
transform 1 0 1568 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_18
timestamp 1698431365
transform 1 0 3360 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_27
timestamp 1698431365
transform 1 0 4368 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_31
timestamp 1698431365
transform 1 0 4816 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_39
timestamp 1698431365
transform 1 0 5712 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_78
timestamp 1698431365
transform 1 0 10080 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_95
timestamp 1698431365
transform 1 0 11984 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_125
timestamp 1698431365
transform 1 0 15344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_129
timestamp 1698431365
transform 1 0 15792 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_137
timestamp 1698431365
transform 1 0 16688 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_171
timestamp 1698431365
transform 1 0 20496 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_181
timestamp 1698431365
transform 1 0 21616 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_185
timestamp 1698431365
transform 1 0 22064 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_189
timestamp 1698431365
transform 1 0 22512 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_191
timestamp 1698431365
transform 1 0 22736 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_194
timestamp 1698431365
transform 1 0 23072 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_198
timestamp 1698431365
transform 1 0 23520 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_208
timestamp 1698431365
transform 1 0 24640 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_212
timestamp 1698431365
transform 1 0 25088 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_228
timestamp 1698431365
transform 1 0 26880 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_239
timestamp 1698431365
transform 1 0 28112 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_243
timestamp 1698431365
transform 1 0 28560 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_247
timestamp 1698431365
transform 1 0 29008 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_259
timestamp 1698431365
transform 1 0 30352 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_275
timestamp 1698431365
transform 1 0 32144 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_279
timestamp 1698431365
transform 1 0 32592 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_282
timestamp 1698431365
transform 1 0 32928 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_289
timestamp 1698431365
transform 1 0 33712 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_297
timestamp 1698431365
transform 1 0 34608 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_301
timestamp 1698431365
transform 1 0 35056 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_68_2
timestamp 1698431365
transform 1 0 1568 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_18
timestamp 1698431365
transform 1 0 3360 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_27
timestamp 1698431365
transform 1 0 4368 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_31
timestamp 1698431365
transform 1 0 4816 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_37
timestamp 1698431365
transform 1 0 5488 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_67
timestamp 1698431365
transform 1 0 8848 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_69
timestamp 1698431365
transform 1 0 9072 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_72
timestamp 1698431365
transform 1 0 9408 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_68_76
timestamp 1698431365
transform 1 0 9856 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_92
timestamp 1698431365
transform 1 0 11648 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_96
timestamp 1698431365
transform 1 0 12096 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_99
timestamp 1698431365
transform 1 0 12432 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_103
timestamp 1698431365
transform 1 0 12880 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_68_107
timestamp 1698431365
transform 1 0 13328 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_68_139
timestamp 1698431365
transform 1 0 16912 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_147
timestamp 1698431365
transform 1 0 17808 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_150
timestamp 1698431365
transform 1 0 18144 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_152
timestamp 1698431365
transform 1 0 18368 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_68_155
timestamp 1698431365
transform 1 0 18704 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_163
timestamp 1698431365
transform 1 0 19600 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_166
timestamp 1698431365
transform 1 0 19936 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_170
timestamp 1698431365
transform 1 0 20384 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_174
timestamp 1698431365
transform 1 0 20832 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_177
timestamp 1698431365
transform 1 0 21168 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_181
timestamp 1698431365
transform 1 0 21616 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_187
timestamp 1698431365
transform 1 0 22288 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_191
timestamp 1698431365
transform 1 0 22736 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_211
timestamp 1698431365
transform 1 0 24976 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_68_219
timestamp 1698431365
transform 1 0 25872 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_235
timestamp 1698431365
transform 1 0 27664 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_244
timestamp 1698431365
transform 1 0 28672 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_274
timestamp 1698431365
transform 1 0 32032 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_68_278
timestamp 1698431365
transform 1 0 32480 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_294
timestamp 1698431365
transform 1 0 34272 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_298
timestamp 1698431365
transform 1 0 34720 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_68_317
timestamp 1698431365
transform 1 0 36848 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_325
timestamp 1698431365
transform 1 0 37744 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_329
timestamp 1698431365
transform 1 0 38192 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_69_2
timestamp 1698431365
transform 1 0 1568 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_10
timestamp 1698431365
transform 1 0 2464 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_69_18
timestamp 1698431365
transform 1 0 3360 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_69_50
timestamp 1698431365
transform 1 0 6944 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_66
timestamp 1698431365
transform 1 0 8736 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_69_72
timestamp 1698431365
transform 1 0 9408 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_80
timestamp 1698431365
transform 1 0 10304 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_84
timestamp 1698431365
transform 1 0 10752 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_86
timestamp 1698431365
transform 1 0 10976 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_95
timestamp 1698431365
transform 1 0 11984 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_69_99
timestamp 1698431365
transform 1 0 12432 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_69_131
timestamp 1698431365
transform 1 0 16016 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_139
timestamp 1698431365
transform 1 0 16912 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_142
timestamp 1698431365
transform 1 0 17248 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_149
timestamp 1698431365
transform 1 0 18032 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_69_155
timestamp 1698431365
transform 1 0 18704 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_69_187
timestamp 1698431365
transform 1 0 22288 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_195
timestamp 1698431365
transform 1 0 23184 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_203
timestamp 1698431365
transform 1 0 24080 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_207
timestamp 1698431365
transform 1 0 24528 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_209
timestamp 1698431365
transform 1 0 24752 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_212
timestamp 1698431365
transform 1 0 25088 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_69_216
timestamp 1698431365
transform 1 0 25536 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_224
timestamp 1698431365
transform 1 0 26432 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_254
timestamp 1698431365
transform 1 0 29792 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_258
timestamp 1698431365
transform 1 0 30240 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_262
timestamp 1698431365
transform 1 0 30688 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_69_266
timestamp 1698431365
transform 1 0 31136 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_274
timestamp 1698431365
transform 1 0 32032 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_278
timestamp 1698431365
transform 1 0 32480 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_69_282
timestamp 1698431365
transform 1 0 32928 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_69_314
timestamp 1698431365
transform 1 0 36512 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_330
timestamp 1698431365
transform 1 0 38304 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70_2
timestamp 1698431365
transform 1 0 1568 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_10
timestamp 1698431365
transform 1 0 2464 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_70_18
timestamp 1698431365
transform 1 0 3360 0 1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_34
timestamp 1698431365
transform 1 0 5152 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70_37
timestamp 1698431365
transform 1 0 5488 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_45
timestamp 1698431365
transform 1 0 6384 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_70_52
timestamp 1698431365
transform 1 0 7168 0 1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_70_84
timestamp 1698431365
transform 1 0 10752 0 1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_100
timestamp 1698431365
transform 1 0 12544 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_104
timestamp 1698431365
transform 1 0 12992 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_107
timestamp 1698431365
transform 1 0 13328 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_111
timestamp 1698431365
transform 1 0 13776 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_113
timestamp 1698431365
transform 1 0 14000 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_121
timestamp 1698431365
transform 1 0 14896 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_125
timestamp 1698431365
transform 1 0 15344 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_129
timestamp 1698431365
transform 1 0 15792 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_133
timestamp 1698431365
transform 1 0 16240 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_135
timestamp 1698431365
transform 1 0 16464 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_146
timestamp 1698431365
transform 1 0 17696 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_158
timestamp 1698431365
transform 1 0 19040 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70_162
timestamp 1698431365
transform 1 0 19488 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_170
timestamp 1698431365
transform 1 0 20384 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_174
timestamp 1698431365
transform 1 0 20832 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_177
timestamp 1698431365
transform 1 0 21168 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_181
timestamp 1698431365
transform 1 0 21616 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_183
timestamp 1698431365
transform 1 0 21840 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_242
timestamp 1698431365
transform 1 0 28448 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_244
timestamp 1698431365
transform 1 0 28672 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_270
timestamp 1698431365
transform 1 0 31584 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70_274
timestamp 1698431365
transform 1 0 32032 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_282
timestamp 1698431365
transform 1 0 32928 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_292
timestamp 1698431365
transform 1 0 34048 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_308
timestamp 1698431365
transform 1 0 35840 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_312
timestamp 1698431365
transform 1 0 36288 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_314
timestamp 1698431365
transform 1 0 36512 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70_317
timestamp 1698431365
transform 1 0 36848 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_325
timestamp 1698431365
transform 1 0 37744 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_31
timestamp 1698431365
transform 1 0 4816 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_71_35
timestamp 1698431365
transform 1 0 5264 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_43
timestamp 1698431365
transform 1 0 6160 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_53
timestamp 1698431365
transform 1 0 7280 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_71_57
timestamp 1698431365
transform 1 0 7728 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_65
timestamp 1698431365
transform 1 0 8624 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_69
timestamp 1698431365
transform 1 0 9072 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_71_72
timestamp 1698431365
transform 1 0 9408 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_80
timestamp 1698431365
transform 1 0 10304 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_71_87
timestamp 1698431365
transform 1 0 11088 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_71_101
timestamp 1698431365
transform 1 0 12656 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_109
timestamp 1698431365
transform 1 0 13552 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_127
timestamp 1698431365
transform 1 0 15568 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_129
timestamp 1698431365
transform 1 0 15792 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_134
timestamp 1698431365
transform 1 0 16352 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_151
timestamp 1698431365
transform 1 0 18256 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_185
timestamp 1698431365
transform 1 0 22064 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_189
timestamp 1698431365
transform 1 0 22512 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_193
timestamp 1698431365
transform 1 0 22960 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_197
timestamp 1698431365
transform 1 0 23408 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_201
timestamp 1698431365
transform 1 0 23856 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_209
timestamp 1698431365
transform 1 0 24752 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_71_212
timestamp 1698431365
transform 1 0 25088 0 -1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_228
timestamp 1698431365
transform 1 0 26880 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_268
timestamp 1698431365
transform 1 0 31360 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_272
timestamp 1698431365
transform 1 0 31808 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_282
timestamp 1698431365
transform 1 0 32928 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_296
timestamp 1698431365
transform 1 0 34496 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_300
timestamp 1698431365
transform 1 0 34944 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_316
timestamp 1698431365
transform 1 0 36736 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_72_2
timestamp 1698431365
transform 1 0 1568 0 1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_72_18
timestamp 1698431365
transform 1 0 3360 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_37
timestamp 1698431365
transform 1 0 5488 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_41
timestamp 1698431365
transform 1 0 5936 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_45
timestamp 1698431365
transform 1 0 6384 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_56
timestamp 1698431365
transform 1 0 7616 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_60
timestamp 1698431365
transform 1 0 8064 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_90
timestamp 1698431365
transform 1 0 11424 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_72_94
timestamp 1698431365
transform 1 0 11872 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_102
timestamp 1698431365
transform 1 0 12768 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_104
timestamp 1698431365
transform 1 0 12992 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_107
timestamp 1698431365
transform 1 0 13328 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_140
timestamp 1698431365
transform 1 0 17024 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_144
timestamp 1698431365
transform 1 0 17472 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_206
timestamp 1698431365
transform 1 0 24416 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_72_210
timestamp 1698431365
transform 1 0 24864 0 1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_72_226
timestamp 1698431365
transform 1 0 26656 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_236
timestamp 1698431365
transform 1 0 27776 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_240
timestamp 1698431365
transform 1 0 28224 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_244
timestamp 1698431365
transform 1 0 28672 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_247
timestamp 1698431365
transform 1 0 29008 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_313
timestamp 1698431365
transform 1 0 36400 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_326
timestamp 1698431365
transform 1 0 37856 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_330
timestamp 1698431365
transform 1 0 38304 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_73_2
timestamp 1698431365
transform 1 0 1568 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_18
timestamp 1698431365
transform 1 0 3360 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_20
timestamp 1698431365
transform 1 0 3584 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_50
timestamp 1698431365
transform 1 0 6944 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_54
timestamp 1698431365
transform 1 0 7392 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_58
timestamp 1698431365
transform 1 0 7840 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_62
timestamp 1698431365
transform 1 0 8288 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_66
timestamp 1698431365
transform 1 0 8736 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_80
timestamp 1698431365
transform 1 0 10304 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_113
timestamp 1698431365
transform 1 0 14000 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_131
timestamp 1698431365
transform 1 0 16016 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_133
timestamp 1698431365
transform 1 0 16240 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_136
timestamp 1698431365
transform 1 0 16576 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_150
timestamp 1698431365
transform 1 0 18144 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_193
timestamp 1698431365
transform 1 0 22960 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_197
timestamp 1698431365
transform 1 0 23408 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_199
timestamp 1698431365
transform 1 0 23632 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_212
timestamp 1698431365
transform 1 0 25088 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_73_216
timestamp 1698431365
transform 1 0 25536 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_224
timestamp 1698431365
transform 1 0 26432 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_228
timestamp 1698431365
transform 1 0 26880 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_230
timestamp 1698431365
transform 1 0 27104 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_275
timestamp 1698431365
transform 1 0 32144 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_329
timestamp 1698431365
transform 1 0 38192 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_31
timestamp 1698431365
transform 1 0 4816 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_43
timestamp 1698431365
transform 1 0 6160 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_47
timestamp 1698431365
transform 1 0 6608 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_49
timestamp 1698431365
transform 1 0 6832 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_97
timestamp 1698431365
transform 1 0 12208 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_101
timestamp 1698431365
transform 1 0 12656 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_136
timestamp 1698431365
transform 1 0 16576 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_74_140
timestamp 1698431365
transform 1 0 17024 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_148
timestamp 1698431365
transform 1 0 17920 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_193
timestamp 1698431365
transform 1 0 22960 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_206
timestamp 1698431365
transform 1 0 24416 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_210
timestamp 1698431365
transform 1 0 24864 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_212
timestamp 1698431365
transform 1 0 25088 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_221
timestamp 1698431365
transform 1 0 26096 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_74_225
timestamp 1698431365
transform 1 0 26544 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_233
timestamp 1698431365
transform 1 0 27440 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_237
timestamp 1698431365
transform 1 0 27888 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_241
timestamp 1698431365
transform 1 0 28336 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_247
timestamp 1698431365
transform 1 0 29008 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_278
timestamp 1698431365
transform 1 0 32480 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_317
timestamp 1698431365
transform 1 0 36848 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_75_2
timestamp 1698431365
transform 1 0 1568 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_10
timestamp 1698431365
transform 1 0 2464 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_14
timestamp 1698431365
transform 1 0 2912 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_16
timestamp 1698431365
transform 1 0 3136 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_33
timestamp 1698431365
transform 1 0 5040 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_67
timestamp 1698431365
transform 1 0 8848 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_69
timestamp 1698431365
transform 1 0 9072 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_78
timestamp 1698431365
transform 1 0 10080 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_87
timestamp 1698431365
transform 1 0 11088 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_75_91
timestamp 1698431365
transform 1 0 11536 0 -1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_75_123
timestamp 1698431365
transform 1 0 15120 0 -1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_139
timestamp 1698431365
transform 1 0 16912 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_75_142
timestamp 1698431365
transform 1 0 17248 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_150
timestamp 1698431365
transform 1 0 18144 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_154
timestamp 1698431365
transform 1 0 18592 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_156
timestamp 1698431365
transform 1 0 18816 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_164
timestamp 1698431365
transform 1 0 19712 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_168
timestamp 1698431365
transform 1 0 20160 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_171
timestamp 1698431365
transform 1 0 20496 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_175
timestamp 1698431365
transform 1 0 20944 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_179
timestamp 1698431365
transform 1 0 21392 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_75_183
timestamp 1698431365
transform 1 0 21840 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_193
timestamp 1698431365
transform 1 0 22960 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_197
timestamp 1698431365
transform 1 0 23408 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_75_201
timestamp 1698431365
transform 1 0 23856 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_209
timestamp 1698431365
transform 1 0 24752 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_212
timestamp 1698431365
transform 1 0 25088 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_75_219
timestamp 1698431365
transform 1 0 25872 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_227
timestamp 1698431365
transform 1 0 26768 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_231
timestamp 1698431365
transform 1 0 27216 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_235
timestamp 1698431365
transform 1 0 27664 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_76_2
timestamp 1698431365
transform 1 0 1568 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_10
timestamp 1698431365
transform 1 0 2464 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_18
timestamp 1698431365
transform 1 0 3360 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_22
timestamp 1698431365
transform 1 0 3808 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_24
timestamp 1698431365
transform 1 0 4032 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_76_27
timestamp 1698431365
transform 1 0 4368 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_37
timestamp 1698431365
transform 1 0 5488 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_39
timestamp 1698431365
transform 1 0 5712 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_50
timestamp 1698431365
transform 1 0 6944 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_54
timestamp 1698431365
transform 1 0 7392 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_57
timestamp 1698431365
transform 1 0 7728 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_61
timestamp 1698431365
transform 1 0 8176 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_65
timestamp 1698431365
transform 1 0 8624 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_67
timestamp 1698431365
transform 1 0 8848 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_70
timestamp 1698431365
transform 1 0 9184 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_74
timestamp 1698431365
transform 1 0 9632 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_76
timestamp 1698431365
transform 1 0 9856 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_76_79
timestamp 1698431365
transform 1 0 10192 0 1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_76_95
timestamp 1698431365
transform 1 0 11984 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_103
timestamp 1698431365
transform 1 0 12880 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_107
timestamp 1698431365
transform 1 0 13328 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_115
timestamp 1698431365
transform 1 0 14224 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_121
timestamp 1698431365
transform 1 0 14896 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_125
timestamp 1698431365
transform 1 0 15344 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_129
timestamp 1698431365
transform 1 0 15792 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_131
timestamp 1698431365
transform 1 0 16016 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_134
timestamp 1698431365
transform 1 0 16352 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_138
timestamp 1698431365
transform 1 0 16800 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_142
timestamp 1698431365
transform 1 0 17248 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_76_148
timestamp 1698431365
transform 1 0 17920 0 1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_164
timestamp 1698431365
transform 1 0 19712 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_170
timestamp 1698431365
transform 1 0 20384 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_172
timestamp 1698431365
transform 1 0 20608 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_177
timestamp 1698431365
transform 1 0 21168 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_199
timestamp 1698431365
transform 1 0 23632 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_203
timestamp 1698431365
transform 1 0 24080 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_234
timestamp 1698431365
transform 1 0 27552 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_238
timestamp 1698431365
transform 1 0 28000 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_244
timestamp 1698431365
transform 1 0 28672 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_247
timestamp 1698431365
transform 1 0 29008 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_266
timestamp 1698431365
transform 1 0 31136 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_328
timestamp 1698431365
transform 1 0 38080 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_330
timestamp 1698431365
transform 1 0 38304 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_31
timestamp 1698431365
transform 1 0 4816 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_35
timestamp 1698431365
transform 1 0 5264 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_37
timestamp 1698431365
transform 1 0 5488 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_67
timestamp 1698431365
transform 1 0 8848 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_69
timestamp 1698431365
transform 1 0 9072 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_72
timestamp 1698431365
transform 1 0 9408 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_77_82
timestamp 1698431365
transform 1 0 10528 0 -1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_114
timestamp 1698431365
transform 1 0 14112 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_117
timestamp 1698431365
transform 1 0 14448 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_136
timestamp 1698431365
transform 1 0 16576 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_142
timestamp 1698431365
transform 1 0 17248 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_148
timestamp 1698431365
transform 1 0 17920 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_152
timestamp 1698431365
transform 1 0 18368 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_156
timestamp 1698431365
transform 1 0 18816 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_212
timestamp 1698431365
transform 1 0 25088 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_214
timestamp 1698431365
transform 1 0 25312 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_77_221
timestamp 1698431365
transform 1 0 26096 0 -1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_77_237
timestamp 1698431365
transform 1 0 27888 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_245
timestamp 1698431365
transform 1 0 28784 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_256
timestamp 1698431365
transform 1 0 30016 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_258
timestamp 1698431365
transform 1 0 30240 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_325
timestamp 1698431365
transform 1 0 37744 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_330
timestamp 1698431365
transform 1 0 38304 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_78_2
timestamp 1698431365
transform 1 0 1568 0 1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_34
timestamp 1698431365
transform 1 0 5152 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_37
timestamp 1698431365
transform 1 0 5488 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_41
timestamp 1698431365
transform 1 0 5936 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_43
timestamp 1698431365
transform 1 0 6160 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_78_50
timestamp 1698431365
transform 1 0 6944 0 1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_66
timestamp 1698431365
transform 1 0 8736 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_96
timestamp 1698431365
transform 1 0 12096 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_100
timestamp 1698431365
transform 1 0 12544 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_104
timestamp 1698431365
transform 1 0 12992 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_115
timestamp 1698431365
transform 1 0 14224 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_144
timestamp 1698431365
transform 1 0 17472 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_203
timestamp 1698431365
transform 1 0 24080 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_234
timestamp 1698431365
transform 1 0 27552 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_238
timestamp 1698431365
transform 1 0 28000 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_242
timestamp 1698431365
transform 1 0 28448 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_244
timestamp 1698431365
transform 1 0 28672 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_247
timestamp 1698431365
transform 1 0 29008 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_269
timestamp 1698431365
transform 1 0 31472 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_271
timestamp 1698431365
transform 1 0 31696 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_317
timestamp 1698431365
transform 1 0 36848 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_79_2
timestamp 1698431365
transform 1 0 1568 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_66
timestamp 1698431365
transform 1 0 8736 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_79_72
timestamp 1698431365
transform 1 0 9408 0 -1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_136
timestamp 1698431365
transform 1 0 16576 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_179
timestamp 1698431365
transform 1 0 21392 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_209
timestamp 1698431365
transform 1 0 24752 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_212
timestamp 1698431365
transform 1 0 25088 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_216
timestamp 1698431365
transform 1 0 25536 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_220
timestamp 1698431365
transform 1 0 25984 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_224
timestamp 1698431365
transform 1 0 26432 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_228
timestamp 1698431365
transform 1 0 26880 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_232
timestamp 1698431365
transform 1 0 27328 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_238
timestamp 1698431365
transform 1 0 28000 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_270
timestamp 1698431365
transform 1 0 31584 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_282
timestamp 1698431365
transform 1 0 32928 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_80_2
timestamp 1698431365
transform 1 0 1568 0 1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_18
timestamp 1698431365
transform 1 0 3360 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_20
timestamp 1698431365
transform 1 0 3584 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_29
timestamp 1698431365
transform 1 0 4592 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_33
timestamp 1698431365
transform 1 0 5040 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_80_37
timestamp 1698431365
transform 1 0 5488 0 1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_53
timestamp 1698431365
transform 1 0 7280 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_80_65
timestamp 1698431365
transform 1 0 8624 0 1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_97
timestamp 1698431365
transform 1 0 12208 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_101
timestamp 1698431365
transform 1 0 12656 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_118
timestamp 1698431365
transform 1 0 14560 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_135
timestamp 1698431365
transform 1 0 16464 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_137
timestamp 1698431365
transform 1 0 16688 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_183
timestamp 1698431365
transform 1 0 21840 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_187
timestamp 1698431365
transform 1 0 22288 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_191
timestamp 1698431365
transform 1 0 22736 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_200
timestamp 1698431365
transform 1 0 23744 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_202
timestamp 1698431365
transform 1 0 23968 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_226
timestamp 1698431365
transform 1 0 26656 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_230
timestamp 1698431365
transform 1 0 27104 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_234
timestamp 1698431365
transform 1 0 27552 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_247
timestamp 1698431365
transform 1 0 29008 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_272
timestamp 1698431365
transform 1 0 31808 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_81_2
timestamp 1698431365
transform 1 0 1568 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_10
timestamp 1698431365
transform 1 0 2464 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_41
timestamp 1698431365
transform 1 0 5936 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_45
timestamp 1698431365
transform 1 0 6384 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_49
timestamp 1698431365
transform 1 0 6832 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_81_56
timestamp 1698431365
transform 1 0 7616 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_64
timestamp 1698431365
transform 1 0 8512 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_66
timestamp 1698431365
transform 1 0 8736 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_69
timestamp 1698431365
transform 1 0 9072 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_72
timestamp 1698431365
transform 1 0 9408 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_78
timestamp 1698431365
transform 1 0 10080 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_82
timestamp 1698431365
transform 1 0 10528 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_86
timestamp 1698431365
transform 1 0 10976 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_90
timestamp 1698431365
transform 1 0 11424 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_135
timestamp 1698431365
transform 1 0 16464 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_139
timestamp 1698431365
transform 1 0 16912 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_179
timestamp 1698431365
transform 1 0 21392 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_185
timestamp 1698431365
transform 1 0 22064 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_206
timestamp 1698431365
transform 1 0 24416 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_220
timestamp 1698431365
transform 1 0 25984 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_224
timestamp 1698431365
transform 1 0 26432 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_81_228
timestamp 1698431365
transform 1 0 26880 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_236
timestamp 1698431365
transform 1 0 27776 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_240
timestamp 1698431365
transform 1 0 28224 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_268
timestamp 1698431365
transform 1 0 31360 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_272
timestamp 1698431365
transform 1 0 31808 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_274
timestamp 1698431365
transform 1 0 32032 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_282
timestamp 1698431365
transform 1 0 32928 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_82_2
timestamp 1698431365
transform 1 0 1568 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_10
timestamp 1698431365
transform 1 0 2464 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_14
timestamp 1698431365
transform 1 0 2912 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_16
timestamp 1698431365
transform 1 0 3136 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_31
timestamp 1698431365
transform 1 0 4816 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_37
timestamp 1698431365
transform 1 0 5488 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_67
timestamp 1698431365
transform 1 0 8848 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_92
timestamp 1698431365
transform 1 0 11648 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_82_96
timestamp 1698431365
transform 1 0 12096 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_104
timestamp 1698431365
transform 1 0 12992 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_107
timestamp 1698431365
transform 1 0 13328 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_111
timestamp 1698431365
transform 1 0 13776 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_117
timestamp 1698431365
transform 1 0 14448 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_119
timestamp 1698431365
transform 1 0 14672 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_122
timestamp 1698431365
transform 1 0 15008 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_126
timestamp 1698431365
transform 1 0 15456 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_177
timestamp 1698431365
transform 1 0 21168 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_181
timestamp 1698431365
transform 1 0 21616 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_218
timestamp 1698431365
transform 1 0 25760 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_82_222
timestamp 1698431365
transform 1 0 26208 0 1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_238
timestamp 1698431365
transform 1 0 28000 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_242
timestamp 1698431365
transform 1 0 28448 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_244
timestamp 1698431365
transform 1 0 28672 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_264
timestamp 1698431365
transform 1 0 30912 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_268
timestamp 1698431365
transform 1 0 31360 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_274
timestamp 1698431365
transform 1 0 32032 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_278
timestamp 1698431365
transform 1 0 32480 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_280
timestamp 1698431365
transform 1 0 32704 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_325
timestamp 1698431365
transform 1 0 37744 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_329
timestamp 1698431365
transform 1 0 38192 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_31
timestamp 1698431365
transform 1 0 4816 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_83_35
timestamp 1698431365
transform 1 0 5264 0 -1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_83_51
timestamp 1698431365
transform 1 0 7056 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_59
timestamp 1698431365
transform 1 0 7952 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_83_61
timestamp 1698431365
transform 1 0 8176 0 -1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_72
timestamp 1698431365
transform 1 0 9408 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_124
timestamp 1698431365
transform 1 0 15232 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_128
timestamp 1698431365
transform 1 0 15680 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_132
timestamp 1698431365
transform 1 0 16128 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_136
timestamp 1698431365
transform 1 0 16576 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_194
timestamp 1698431365
transform 1 0 23072 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_198
timestamp 1698431365
transform 1 0 23520 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_202
timestamp 1698431365
transform 1 0 23968 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_206
timestamp 1698431365
transform 1 0 24416 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_83_212
timestamp 1698431365
transform 1 0 25088 0 -1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_244
timestamp 1698431365
transform 1 0 28672 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_83_246
timestamp 1698431365
transform 1 0 28896 0 -1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_253
timestamp 1698431365
transform 1 0 29680 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_83_255
timestamp 1698431365
transform 1 0 29904 0 -1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_258
timestamp 1698431365
transform 1 0 30240 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_262
timestamp 1698431365
transform 1 0 30688 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_266
timestamp 1698431365
transform 1 0 31136 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_83_270
timestamp 1698431365
transform 1 0 31584 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_278
timestamp 1698431365
transform 1 0 32480 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_282
timestamp 1698431365
transform 1 0 32928 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_83_284
timestamp 1698431365
transform 1 0 33152 0 -1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_84_2
timestamp 1698431365
transform 1 0 1568 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_10
timestamp 1698431365
transform 1 0 2464 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_84_18
timestamp 1698431365
transform 1 0 3360 0 1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_34
timestamp 1698431365
transform 1 0 5152 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_37
timestamp 1698431365
transform 1 0 5488 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_84_41
timestamp 1698431365
transform 1 0 5936 0 1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_63
timestamp 1698431365
transform 1 0 8400 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_67
timestamp 1698431365
transform 1 0 8848 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_69
timestamp 1698431365
transform 1 0 9072 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_84_72
timestamp 1698431365
transform 1 0 9408 0 1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_104
timestamp 1698431365
transform 1 0 12992 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_84_107
timestamp 1698431365
transform 1 0 13328 0 1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_84_123
timestamp 1698431365
transform 1 0 15120 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_131
timestamp 1698431365
transform 1 0 16016 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_135
timestamp 1698431365
transform 1 0 16464 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_137
timestamp 1698431365
transform 1 0 16688 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_140
timestamp 1698431365
transform 1 0 17024 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_150
timestamp 1698431365
transform 1 0 18144 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_156
timestamp 1698431365
transform 1 0 18816 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_166
timestamp 1698431365
transform 1 0 19936 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_177
timestamp 1698431365
transform 1 0 21168 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_84_181
timestamp 1698431365
transform 1 0 21616 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_189
timestamp 1698431365
transform 1 0 22512 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_193
timestamp 1698431365
transform 1 0 22960 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_196
timestamp 1698431365
transform 1 0 23296 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_200
timestamp 1698431365
transform 1 0 23744 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_231
timestamp 1698431365
transform 1 0 27216 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_84_235
timestamp 1698431365
transform 1 0 27664 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_243
timestamp 1698431365
transform 1 0 28560 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_247
timestamp 1698431365
transform 1 0 29008 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_251
timestamp 1698431365
transform 1 0 29456 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_254
timestamp 1698431365
transform 1 0 29792 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_264
timestamp 1698431365
transform 1 0 30912 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_268
timestamp 1698431365
transform 1 0 31360 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_275
timestamp 1698431365
transform 1 0 32144 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_279
timestamp 1698431365
transform 1 0 32592 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_281
timestamp 1698431365
transform 1 0 32816 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_314
timestamp 1698431365
transform 1 0 36512 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_327
timestamp 1698431365
transform 1 0 37968 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_85_2
timestamp 1698431365
transform 1 0 1568 0 -1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_85_24
timestamp 1698431365
transform 1 0 4032 0 -1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_39
timestamp 1698431365
transform 1 0 5712 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_80
timestamp 1698431365
transform 1 0 10304 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_85_84
timestamp 1698431365
transform 1 0 10752 0 -1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_85_116
timestamp 1698431365
transform 1 0 14336 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_85_124
timestamp 1698431365
transform 1 0 15232 0 -1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_127
timestamp 1698431365
transform 1 0 15568 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_137
timestamp 1698431365
transform 1 0 16688 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_85_139
timestamp 1698431365
transform 1 0 16912 0 -1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_171
timestamp 1698431365
transform 1 0 20496 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_85_179
timestamp 1698431365
transform 1 0 21392 0 -1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_85_195
timestamp 1698431365
transform 1 0 23184 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_203
timestamp 1698431365
transform 1 0 24080 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_207
timestamp 1698431365
transform 1 0 24528 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_85_209
timestamp 1698431365
transform 1 0 24752 0 -1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_85_212
timestamp 1698431365
transform 1 0 25088 0 -1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_85_228
timestamp 1698431365
transform 1 0 26880 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_236
timestamp 1698431365
transform 1 0 27776 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_245
timestamp 1698431365
transform 1 0 28784 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_249
timestamp 1698431365
transform 1 0 29232 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_253
timestamp 1698431365
transform 1 0 29680 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_257
timestamp 1698431365
transform 1 0 30128 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_261
timestamp 1698431365
transform 1 0 30576 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_286
timestamp 1698431365
transform 1 0 33376 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_2
timestamp 1698431365
transform 1 0 1568 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_45
timestamp 1698431365
transform 1 0 6384 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_49
timestamp 1698431365
transform 1 0 6832 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_86_53
timestamp 1698431365
transform 1 0 7280 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_61
timestamp 1698431365
transform 1 0 8176 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_71
timestamp 1698431365
transform 1 0 9296 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_75
timestamp 1698431365
transform 1 0 9744 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_79
timestamp 1698431365
transform 1 0 10192 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_85
timestamp 1698431365
transform 1 0 10864 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_86_93
timestamp 1698431365
transform 1 0 11760 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_101
timestamp 1698431365
transform 1 0 12656 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_107
timestamp 1698431365
transform 1 0 13328 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_111
timestamp 1698431365
transform 1 0 13776 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_115
timestamp 1698431365
transform 1 0 14224 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_86_152
timestamp 1698431365
transform 1 0 18368 0 1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_168
timestamp 1698431365
transform 1 0 20160 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_172
timestamp 1698431365
transform 1 0 20608 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_174
timestamp 1698431365
transform 1 0 20832 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_177
timestamp 1698431365
transform 1 0 21168 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_181
timestamp 1698431365
transform 1 0 21616 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_183
timestamp 1698431365
transform 1 0 21840 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_222
timestamp 1698431365
transform 1 0 26208 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_224
timestamp 1698431365
transform 1 0 26432 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_229
timestamp 1698431365
transform 1 0 26992 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_231
timestamp 1698431365
transform 1 0 27216 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_243
timestamp 1698431365
transform 1 0 28560 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_255
timestamp 1698431365
transform 1 0 29904 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_277
timestamp 1698431365
transform 1 0 32368 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_288
timestamp 1698431365
transform 1 0 33600 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_290
timestamp 1698431365
transform 1 0 33824 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_327
timestamp 1698431365
transform 1 0 37968 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_87_2
timestamp 1698431365
transform 1 0 1568 0 -1 70560
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_87_34
timestamp 1698431365
transform 1 0 5152 0 -1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_64
timestamp 1698431365
transform 1 0 8512 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_68
timestamp 1698431365
transform 1 0 8960 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_72
timestamp 1698431365
transform 1 0 9408 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_87_74
timestamp 1698431365
transform 1 0 9632 0 -1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_122
timestamp 1698431365
transform 1 0 15008 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_131
timestamp 1698431365
transform 1 0 16016 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_135
timestamp 1698431365
transform 1 0 16464 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_87_139
timestamp 1698431365
transform 1 0 16912 0 -1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_142
timestamp 1698431365
transform 1 0 17248 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_87_146
timestamp 1698431365
transform 1 0 17696 0 -1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_184
timestamp 1698431365
transform 1 0 21952 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_87_188
timestamp 1698431365
transform 1 0 22400 0 -1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_204
timestamp 1698431365
transform 1 0 24192 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_208
timestamp 1698431365
transform 1 0 24640 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_212
timestamp 1698431365
transform 1 0 25088 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_216
timestamp 1698431365
transform 1 0 25536 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_229
timestamp 1698431365
transform 1 0 26992 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_269
timestamp 1698431365
transform 1 0 31472 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_277
timestamp 1698431365
transform 1 0 32368 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_87_279
timestamp 1698431365
transform 1 0 32592 0 -1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_324
timestamp 1698431365
transform 1 0 37632 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_328
timestamp 1698431365
transform 1 0 38080 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_87_330
timestamp 1698431365
transform 1 0 38304 0 -1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_88_2
timestamp 1698431365
transform 1 0 1568 0 1 70560
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_34
timestamp 1698431365
transform 1 0 5152 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_43
timestamp 1698431365
transform 1 0 6160 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_115
timestamp 1698431365
transform 1 0 14224 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_149
timestamp 1698431365
transform 1 0 18032 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_154
timestamp 1698431365
transform 1 0 18592 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_88_158
timestamp 1698431365
transform 1 0 19040 0 1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_174
timestamp 1698431365
transform 1 0 20832 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_203
timestamp 1698431365
transform 1 0 24080 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_207
timestamp 1698431365
transform 1 0 24528 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_209
timestamp 1698431365
transform 1 0 24752 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_220
timestamp 1698431365
transform 1 0 25984 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_222
timestamp 1698431365
transform 1 0 26208 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_244
timestamp 1698431365
transform 1 0 28672 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_89_2
timestamp 1698431365
transform 1 0 1568 0 -1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_89_34
timestamp 1698431365
transform 1 0 5152 0 -1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_89_50
timestamp 1698431365
transform 1 0 6944 0 -1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_58
timestamp 1698431365
transform 1 0 7840 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_89_62
timestamp 1698431365
transform 1 0 8288 0 -1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_89_69
timestamp 1698431365
transform 1 0 9072 0 -1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_72
timestamp 1698431365
transform 1 0 9408 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_78
timestamp 1698431365
transform 1 0 10080 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_82
timestamp 1698431365
transform 1 0 10528 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_89_84
timestamp 1698431365
transform 1 0 10752 0 -1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_114
timestamp 1698431365
transform 1 0 14112 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_89_118
timestamp 1698431365
transform 1 0 14560 0 -1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_134
timestamp 1698431365
transform 1 0 16352 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_138
timestamp 1698431365
transform 1 0 16800 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_142
timestamp 1698431365
transform 1 0 17248 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_89_146
timestamp 1698431365
transform 1 0 17696 0 -1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_89_154
timestamp 1698431365
transform 1 0 18592 0 -1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_212
timestamp 1698431365
transform 1 0 25088 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_89_214
timestamp 1698431365
transform 1 0 25312 0 -1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_275
timestamp 1698431365
transform 1 0 32144 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_89_279
timestamp 1698431365
transform 1 0 32592 0 -1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_282
timestamp 1698431365
transform 1 0 32928 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_302
timestamp 1698431365
transform 1 0 35168 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_314
timestamp 1698431365
transform 1 0 36512 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_318
timestamp 1698431365
transform 1 0 36960 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_322
timestamp 1698431365
transform 1 0 37408 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_326
timestamp 1698431365
transform 1 0 37856 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_89_330
timestamp 1698431365
transform 1 0 38304 0 -1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_90_2
timestamp 1698431365
transform 1 0 1568 0 1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_34
timestamp 1698431365
transform 1 0 5152 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_90_37
timestamp 1698431365
transform 1 0 5488 0 1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_90_69
timestamp 1698431365
transform 1 0 9072 0 1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_85
timestamp 1698431365
transform 1 0 10864 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_89
timestamp 1698431365
transform 1 0 11312 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_90_96
timestamp 1698431365
transform 1 0 12096 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_104
timestamp 1698431365
transform 1 0 12992 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_113
timestamp 1698431365
transform 1 0 14000 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_117
timestamp 1698431365
transform 1 0 14448 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_168
timestamp 1698431365
transform 1 0 20160 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_172
timestamp 1698431365
transform 1 0 20608 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_174
timestamp 1698431365
transform 1 0 20832 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_90_177
timestamp 1698431365
transform 1 0 21168 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_185
timestamp 1698431365
transform 1 0 22064 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_243
timestamp 1698431365
transform 1 0 28560 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_265
timestamp 1698431365
transform 1 0 31024 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_269
timestamp 1698431365
transform 1 0 31472 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_90_275
timestamp 1698431365
transform 1 0 32144 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_283
timestamp 1698431365
transform 1 0 33040 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_287
timestamp 1698431365
transform 1 0 33488 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_290
timestamp 1698431365
transform 1 0 33824 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_294
timestamp 1698431365
transform 1 0 34272 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_304
timestamp 1698431365
transform 1 0 35392 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_308
timestamp 1698431365
transform 1 0 35840 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_312
timestamp 1698431365
transform 1 0 36288 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_314
timestamp 1698431365
transform 1 0 36512 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_90_317
timestamp 1698431365
transform 1 0 36848 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_325
timestamp 1698431365
transform 1 0 37744 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_329
timestamp 1698431365
transform 1 0 38192 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_91_2
timestamp 1698431365
transform 1 0 1568 0 -1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_34
timestamp 1698431365
transform 1 0 5152 0 -1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_37
timestamp 1698431365
transform 1 0 5488 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_41
timestamp 1698431365
transform 1 0 5936 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_91_45
timestamp 1698431365
transform 1 0 6384 0 -1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_91_61
timestamp 1698431365
transform 1 0 8176 0 -1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_69
timestamp 1698431365
transform 1 0 9072 0 -1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_91_72
timestamp 1698431365
transform 1 0 9408 0 -1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_104
timestamp 1698431365
transform 1 0 12992 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_108
timestamp 1698431365
transform 1 0 13440 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_110
timestamp 1698431365
transform 1 0 13664 0 -1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_150
timestamp 1698431365
transform 1 0 18144 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_154
timestamp 1698431365
transform 1 0 18592 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_158
timestamp 1698431365
transform 1 0 19040 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_212
timestamp 1698431365
transform 1 0 25088 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_214
timestamp 1698431365
transform 1 0 25312 0 -1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_263
timestamp 1698431365
transform 1 0 30800 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_267
timestamp 1698431365
transform 1 0 31248 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_91_271
timestamp 1698431365
transform 1 0 31696 0 -1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_279
timestamp 1698431365
transform 1 0 32592 0 -1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_91_282
timestamp 1698431365
transform 1 0 32928 0 -1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_91_314
timestamp 1698431365
transform 1 0 36512 0 -1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_330
timestamp 1698431365
transform 1 0 38304 0 -1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_2
timestamp 1698431365
transform 1 0 1568 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_37
timestamp 1698431365
transform 1 0 5488 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_43
timestamp 1698431365
transform 1 0 6160 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_45
timestamp 1698431365
transform 1 0 6384 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_51
timestamp 1698431365
transform 1 0 7056 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_55
timestamp 1698431365
transform 1 0 7504 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_59
timestamp 1698431365
transform 1 0 7952 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_92_65
timestamp 1698431365
transform 1 0 8624 0 1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_92_97
timestamp 1698431365
transform 1 0 12208 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_107
timestamp 1698431365
transform 1 0 13328 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_111
timestamp 1698431365
transform 1 0 13776 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_113
timestamp 1698431365
transform 1 0 14000 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_152
timestamp 1698431365
transform 1 0 18368 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_156
timestamp 1698431365
transform 1 0 18816 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_160
timestamp 1698431365
transform 1 0 19264 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_172
timestamp 1698431365
transform 1 0 20608 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_174
timestamp 1698431365
transform 1 0 20832 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_177
timestamp 1698431365
transform 1 0 21168 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_181
timestamp 1698431365
transform 1 0 21616 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_243
timestamp 1698431365
transform 1 0 28560 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_252
timestamp 1698431365
transform 1 0 29568 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_256
timestamp 1698431365
transform 1 0 30016 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_260
timestamp 1698431365
transform 1 0 30464 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_92_264
timestamp 1698431365
transform 1 0 30912 0 1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_280
timestamp 1698431365
transform 1 0 32704 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_284
timestamp 1698431365
transform 1 0 33152 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_293
timestamp 1698431365
transform 1 0 34160 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_297
timestamp 1698431365
transform 1 0 34608 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_299
timestamp 1698431365
transform 1 0 34832 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_314
timestamp 1698431365
transform 1 0 36512 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_92_317
timestamp 1698431365
transform 1 0 36848 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_325
timestamp 1698431365
transform 1 0 37744 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_93_2
timestamp 1698431365
transform 1 0 1568 0 -1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_93_18
timestamp 1698431365
transform 1 0 3360 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_63
timestamp 1698431365
transform 1 0 8400 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_67
timestamp 1698431365
transform 1 0 8848 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_69
timestamp 1698431365
transform 1 0 9072 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_93_72
timestamp 1698431365
transform 1 0 9408 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_80
timestamp 1698431365
transform 1 0 10304 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_84
timestamp 1698431365
transform 1 0 10752 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_93_114
timestamp 1698431365
transform 1 0 14112 0 -1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_93_130
timestamp 1698431365
transform 1 0 15904 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_138
timestamp 1698431365
transform 1 0 16800 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_142
timestamp 1698431365
transform 1 0 17248 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_144
timestamp 1698431365
transform 1 0 17472 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_155
timestamp 1698431365
transform 1 0 18704 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_185
timestamp 1698431365
transform 1 0 22064 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_187
timestamp 1698431365
transform 1 0 22288 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_204
timestamp 1698431365
transform 1 0 24192 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_220
timestamp 1698431365
transform 1 0 25984 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_268
timestamp 1698431365
transform 1 0 31360 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_270
timestamp 1698431365
transform 1 0 31584 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_273
timestamp 1698431365
transform 1 0 31920 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_277
timestamp 1698431365
transform 1 0 32368 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_288
timestamp 1698431365
transform 1 0 33600 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_322
timestamp 1698431365
transform 1 0 37408 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_94_2
timestamp 1698431365
transform 1 0 1568 0 1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_94_34
timestamp 1698431365
transform 1 0 5152 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_94_37
timestamp 1698431365
transform 1 0 5488 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_94_47
timestamp 1698431365
transform 1 0 6608 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_94_51
timestamp 1698431365
transform 1 0 7056 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_94_84
timestamp 1698431365
transform 1 0 10752 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_94_88
timestamp 1698431365
transform 1 0 11200 0 1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_94_104
timestamp 1698431365
transform 1 0 12992 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_94_107
timestamp 1698431365
transform 1 0 13328 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_94_115
timestamp 1698431365
transform 1 0 14224 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_94_117
timestamp 1698431365
transform 1 0 14448 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_94_120
timestamp 1698431365
transform 1 0 14784 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_94_124
timestamp 1698431365
transform 1 0 15232 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_94_128
timestamp 1698431365
transform 1 0 15680 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_94_170
timestamp 1698431365
transform 1 0 20384 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_94_172
timestamp 1698431365
transform 1 0 20608 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_94_247
timestamp 1698431365
transform 1 0 29008 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_94_251
timestamp 1698431365
transform 1 0 29456 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_94_253
timestamp 1698431365
transform 1 0 29680 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_94_279
timestamp 1698431365
transform 1 0 32592 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_94_283
timestamp 1698431365
transform 1 0 33040 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_94_285
timestamp 1698431365
transform 1 0 33264 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_94_314
timestamp 1698431365
transform 1 0 36512 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_94_325
timestamp 1698431365
transform 1 0 37744 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_94_329
timestamp 1698431365
transform 1 0 38192 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_95_2
timestamp 1698431365
transform 1 0 1568 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_95_34
timestamp 1698431365
transform 1 0 5152 0 -1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_95_50
timestamp 1698431365
transform 1 0 6944 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_95_58
timestamp 1698431365
transform 1 0 7840 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_81
timestamp 1698431365
transform 1 0 10416 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_85
timestamp 1698431365
transform 1 0 10864 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_95_118
timestamp 1698431365
transform 1 0 14560 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_124
timestamp 1698431365
transform 1 0 15232 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_128
timestamp 1698431365
transform 1 0 15680 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_150
timestamp 1698431365
transform 1 0 18144 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_95_152
timestamp 1698431365
transform 1 0 18368 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_203
timestamp 1698431365
transform 1 0 24080 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_207
timestamp 1698431365
transform 1 0 24528 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_95_209
timestamp 1698431365
transform 1 0 24752 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_220
timestamp 1698431365
transform 1 0 25984 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_243
timestamp 1698431365
transform 1 0 28560 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_95_245
timestamp 1698431365
transform 1 0 28784 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_273
timestamp 1698431365
transform 1 0 31920 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_282
timestamp 1698431365
transform 1 0 32928 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_95_300
timestamp 1698431365
transform 1 0 34944 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_329
timestamp 1698431365
transform 1 0 38192 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_96_2
timestamp 1698431365
transform 1 0 1568 0 1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_96_34
timestamp 1698431365
transform 1 0 5152 0 1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_96_37
timestamp 1698431365
transform 1 0 5488 0 1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_96_45
timestamp 1698431365
transform 1 0 6384 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_96_49
timestamp 1698431365
transform 1 0 6832 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_96_51
timestamp 1698431365
transform 1 0 7056 0 1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_96_81
timestamp 1698431365
transform 1 0 10416 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_96_85
timestamp 1698431365
transform 1 0 10864 0 1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_96_93
timestamp 1698431365
transform 1 0 11760 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_96_107
timestamp 1698431365
transform 1 0 13328 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_96_243
timestamp 1698431365
transform 1 0 28560 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_96_247
timestamp 1698431365
transform 1 0 29008 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_96_251
timestamp 1698431365
transform 1 0 29456 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_96_255
timestamp 1698431365
transform 1 0 29904 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_96_259
timestamp 1698431365
transform 1 0 30352 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_96_263
timestamp 1698431365
transform 1 0 30800 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_96_281
timestamp 1698431365
transform 1 0 32816 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_96_290
timestamp 1698431365
transform 1 0 33824 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_97_2
timestamp 1698431365
transform 1 0 1568 0 -1 78400
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_97_18
timestamp 1698431365
transform 1 0 3360 0 -1 78400
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_97_48
timestamp 1698431365
transform 1 0 6720 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_97_52
timestamp 1698431365
transform 1 0 7168 0 -1 78400
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_97_78
timestamp 1698431365
transform 1 0 10080 0 -1 78400
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_97_94
timestamp 1698431365
transform 1 0 11872 0 -1 78400
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_97_102
timestamp 1698431365
transform 1 0 12768 0 -1 78400
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_97_134
timestamp 1698431365
transform 1 0 16352 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_97_150
timestamp 1698431365
transform 1 0 18144 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_97_206
timestamp 1698431365
transform 1 0 24416 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_97_236
timestamp 1698431365
transform 1 0 27776 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_97_240
timestamp 1698431365
transform 1 0 28224 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_97_244
timestamp 1698431365
transform 1 0 28672 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_97_273
timestamp 1698431365
transform 1 0 31920 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_97_277
timestamp 1698431365
transform 1 0 32368 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_97_279
timestamp 1698431365
transform 1 0 32592 0 -1 78400
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_97_282
timestamp 1698431365
transform 1 0 32928 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_97_286
timestamp 1698431365
transform 1 0 33376 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_97_290
timestamp 1698431365
transform 1 0 33824 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_97_322
timestamp 1698431365
transform 1 0 37408 0 -1 78400
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_97_330
timestamp 1698431365
transform 1 0 38304 0 -1 78400
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_98_2
timestamp 1698431365
transform 1 0 1568 0 1 78400
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_98_34
timestamp 1698431365
transform 1 0 5152 0 1 78400
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98_37
timestamp 1698431365
transform 1 0 5488 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_98_39
timestamp 1698431365
transform 1 0 5712 0 1 78400
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98_48
timestamp 1698431365
transform 1 0 6720 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98_85
timestamp 1698431365
transform 1 0 10864 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98_89
timestamp 1698431365
transform 1 0 11312 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_98_101
timestamp 1698431365
transform 1 0 12656 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_98_107
timestamp 1698431365
transform 1 0 13328 0 1 78400
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_98_125
timestamp 1698431365
transform 1 0 15344 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_98_160
timestamp 1698431365
transform 1 0 19264 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_98_164
timestamp 1698431365
transform 1 0 19712 0 1 78400
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98_177
timestamp 1698431365
transform 1 0 21168 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98_195
timestamp 1698431365
transform 1 0 23184 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_98_199
timestamp 1698431365
transform 1 0 23632 0 1 78400
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98_224
timestamp 1698431365
transform 1 0 26432 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_98_226
timestamp 1698431365
transform 1 0 26656 0 1 78400
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98_255
timestamp 1698431365
transform 1 0 29904 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_98_257
timestamp 1698431365
transform 1 0 30128 0 1 78400
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98_275
timestamp 1698431365
transform 1 0 32144 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98_279
timestamp 1698431365
transform 1 0 32592 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98_283
timestamp 1698431365
transform 1 0 33040 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98_287
timestamp 1698431365
transform 1 0 33488 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_98_291
timestamp 1698431365
transform 1 0 33936 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98_295
timestamp 1698431365
transform 1 0 34384 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98_302
timestamp 1698431365
transform 1 0 35168 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98_312
timestamp 1698431365
transform 1 0 36288 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_98_314
timestamp 1698431365
transform 1 0 36512 0 1 78400
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_98_317
timestamp 1698431365
transform 1 0 36848 0 1 78400
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_98_325
timestamp 1698431365
transform 1 0 37744 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98_329
timestamp 1698431365
transform 1 0 38192 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_99_2
timestamp 1698431365
transform 1 0 1568 0 -1 79968
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_99_34
timestamp 1698431365
transform 1 0 5152 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_99_45
timestamp 1698431365
transform 1 0 6384 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_99_47
timestamp 1698431365
transform 1 0 6608 0 -1 79968
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_99_50
timestamp 1698431365
transform 1 0 6944 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_99_54
timestamp 1698431365
transform 1 0 7392 0 -1 79968
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_99_72
timestamp 1698431365
transform 1 0 9408 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_99_76
timestamp 1698431365
transform 1 0 9856 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_99_80
timestamp 1698431365
transform 1 0 10304 0 -1 79968
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_99_112
timestamp 1698431365
transform 1 0 13888 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_99_116
timestamp 1698431365
transform 1 0 14336 0 -1 79968
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_99_124
timestamp 1698431365
transform 1 0 15232 0 -1 79968
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_99_127
timestamp 1698431365
transform 1 0 15568 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_99_131
timestamp 1698431365
transform 1 0 16016 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_99_133
timestamp 1698431365
transform 1 0 16240 0 -1 79968
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_99_136
timestamp 1698431365
transform 1 0 16576 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_99_142
timestamp 1698431365
transform 1 0 17248 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_99_144
timestamp 1698431365
transform 1 0 17472 0 -1 79968
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_99_203
timestamp 1698431365
transform 1 0 24080 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_99_207
timestamp 1698431365
transform 1 0 24528 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_99_209
timestamp 1698431365
transform 1 0 24752 0 -1 79968
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_99_277
timestamp 1698431365
transform 1 0 32368 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_99_279
timestamp 1698431365
transform 1 0 32592 0 -1 79968
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_99_282
timestamp 1698431365
transform 1 0 32928 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_99_286
timestamp 1698431365
transform 1 0 33376 0 -1 79968
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_99_318
timestamp 1698431365
transform 1 0 36960 0 -1 79968
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_99_326
timestamp 1698431365
transform 1 0 37856 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_99_330
timestamp 1698431365
transform 1 0 38304 0 -1 79968
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_100_2
timestamp 1698431365
transform 1 0 1568 0 1 79968
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_100_34
timestamp 1698431365
transform 1 0 5152 0 1 79968
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_100_37
timestamp 1698431365
transform 1 0 5488 0 1 79968
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_100_69
timestamp 1698431365
transform 1 0 9072 0 1 79968
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_100_85
timestamp 1698431365
transform 1 0 10864 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_100_89
timestamp 1698431365
transform 1 0 11312 0 1 79968
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_100_96
timestamp 1698431365
transform 1 0 12096 0 1 79968
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_100_104
timestamp 1698431365
transform 1 0 12992 0 1 79968
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_100_107
timestamp 1698431365
transform 1 0 13328 0 1 79968
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_100_123
timestamp 1698431365
transform 1 0 15120 0 1 79968
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_100_131
timestamp 1698431365
transform 1 0 16016 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_100_177
timestamp 1698431365
transform 1 0 21168 0 1 79968
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_100_244
timestamp 1698431365
transform 1 0 28672 0 1 79968
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_100_247
timestamp 1698431365
transform 1 0 29008 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_100_266
timestamp 1698431365
transform 1 0 31136 0 1 79968
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_100_298
timestamp 1698431365
transform 1 0 34720 0 1 79968
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_100_314
timestamp 1698431365
transform 1 0 36512 0 1 79968
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_100_317
timestamp 1698431365
transform 1 0 36848 0 1 79968
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_100_325
timestamp 1698431365
transform 1 0 37744 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_100_329
timestamp 1698431365
transform 1 0 38192 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_101_2
timestamp 1698431365
transform 1 0 1568 0 -1 81536
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_101_18
timestamp 1698431365
transform 1 0 3360 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_101_49
timestamp 1698431365
transform 1 0 6832 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_101_53
timestamp 1698431365
transform 1 0 7280 0 -1 81536
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_101_61
timestamp 1698431365
transform 1 0 8176 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_101_65
timestamp 1698431365
transform 1 0 8624 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_101_67
timestamp 1698431365
transform 1 0 8848 0 -1 81536
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_101_81
timestamp 1698431365
transform 1 0 10416 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_101_85
timestamp 1698431365
transform 1 0 10864 0 -1 81536
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_101_93
timestamp 1698431365
transform 1 0 11760 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_101_97
timestamp 1698431365
transform 1 0 12208 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_101_111
timestamp 1698431365
transform 1 0 13776 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_101_115
timestamp 1698431365
transform 1 0 14224 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_101_119
timestamp 1698431365
transform 1 0 14672 0 -1 81536
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_101_127
timestamp 1698431365
transform 1 0 15568 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_101_131
timestamp 1698431365
transform 1 0 16016 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_101_133
timestamp 1698431365
transform 1 0 16240 0 -1 81536
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_101_136
timestamp 1698431365
transform 1 0 16576 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_101_222
timestamp 1698431365
transform 1 0 26208 0 -1 81536
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_101_247
timestamp 1698431365
transform 1 0 29008 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_101_251
timestamp 1698431365
transform 1 0 29456 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_101_268
timestamp 1698431365
transform 1 0 31360 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_101_272
timestamp 1698431365
transform 1 0 31808 0 -1 81536
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_101_282
timestamp 1698431365
transform 1 0 32928 0 -1 81536
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_101_314
timestamp 1698431365
transform 1 0 36512 0 -1 81536
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_101_330
timestamp 1698431365
transform 1 0 38304 0 -1 81536
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_102_2
timestamp 1698431365
transform 1 0 1568 0 1 81536
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_102_18
timestamp 1698431365
transform 1 0 3360 0 1 81536
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102_26
timestamp 1698431365
transform 1 0 4256 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102_37
timestamp 1698431365
transform 1 0 5488 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102_49
timestamp 1698431365
transform 1 0 6832 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_102_51
timestamp 1698431365
transform 1 0 7056 0 1 81536
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102_89
timestamp 1698431365
transform 1 0 11312 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_102_93
timestamp 1698431365
transform 1 0 11760 0 1 81536
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102_101
timestamp 1698431365
transform 1 0 12656 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102_107
timestamp 1698431365
transform 1 0 13328 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_102_109
timestamp 1698431365
transform 1 0 13552 0 1 81536
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102_118
timestamp 1698431365
transform 1 0 14560 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102_122
timestamp 1698431365
transform 1 0 15008 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_102_126
timestamp 1698431365
transform 1 0 15456 0 1 81536
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_102_134
timestamp 1698431365
transform 1 0 16352 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102_138
timestamp 1698431365
transform 1 0 16800 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102_173
timestamp 1698431365
transform 1 0 20720 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102_247
timestamp 1698431365
transform 1 0 29008 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_102_249
timestamp 1698431365
transform 1 0 29232 0 1 81536
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102_291
timestamp 1698431365
transform 1 0 33936 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_102_295
timestamp 1698431365
transform 1 0 34384 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102_299
timestamp 1698431365
transform 1 0 34832 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102_309
timestamp 1698431365
transform 1 0 35952 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102_313
timestamp 1698431365
transform 1 0 36400 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_102_317
timestamp 1698431365
transform 1 0 36848 0 1 81536
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_102_325
timestamp 1698431365
transform 1 0 37744 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102_329
timestamp 1698431365
transform 1 0 38192 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_103_2
timestamp 1698431365
transform 1 0 1568 0 -1 83104
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_103_34
timestamp 1698431365
transform 1 0 5152 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_103_38
timestamp 1698431365
transform 1 0 5600 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_103_40
timestamp 1698431365
transform 1 0 5824 0 -1 83104
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_103_81
timestamp 1698431365
transform 1 0 10416 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_103_85
timestamp 1698431365
transform 1 0 10864 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_103_89
timestamp 1698431365
transform 1 0 11312 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_103_124
timestamp 1698431365
transform 1 0 15232 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_103_128
timestamp 1698431365
transform 1 0 15680 0 -1 83104
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_103_136
timestamp 1698431365
transform 1 0 16576 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_103_142
timestamp 1698431365
transform 1 0 17248 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_103_144
timestamp 1698431365
transform 1 0 17472 0 -1 83104
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_103_147
timestamp 1698431365
transform 1 0 17808 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_103_149
timestamp 1698431365
transform 1 0 18032 0 -1 83104
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_103_208
timestamp 1698431365
transform 1 0 24640 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_103_259
timestamp 1698431365
transform 1 0 30352 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_103_263
timestamp 1698431365
transform 1 0 30800 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_103_277
timestamp 1698431365
transform 1 0 32368 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_103_279
timestamp 1698431365
transform 1 0 32592 0 -1 83104
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_103_282
timestamp 1698431365
transform 1 0 32928 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_103_286
timestamp 1698431365
transform 1 0 33376 0 -1 83104
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_103_294
timestamp 1698431365
transform 1 0 34272 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_103_296
timestamp 1698431365
transform 1 0 34496 0 -1 83104
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_103_330
timestamp 1698431365
transform 1 0 38304 0 -1 83104
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_104_2
timestamp 1698431365
transform 1 0 1568 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104_4
timestamp 1698431365
transform 1 0 1792 0 1 83104
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_104_28
timestamp 1698431365
transform 1 0 4480 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_104_32
timestamp 1698431365
transform 1 0 4928 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104_34
timestamp 1698431365
transform 1 0 5152 0 1 83104
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_104_37
timestamp 1698431365
transform 1 0 5488 0 1 83104
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_104_53
timestamp 1698431365
transform 1 0 7280 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_104_57
timestamp 1698431365
transform 1 0 7728 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_104_65
timestamp 1698431365
transform 1 0 8624 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104_69
timestamp 1698431365
transform 1 0 9072 0 1 83104
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_104_72
timestamp 1698431365
transform 1 0 9408 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_104_76
timestamp 1698431365
transform 1 0 9856 0 1 83104
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_104_92
timestamp 1698431365
transform 1 0 11648 0 1 83104
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_104_100
timestamp 1698431365
transform 1 0 12544 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104_102
timestamp 1698431365
transform 1 0 12768 0 1 83104
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_104_107
timestamp 1698431365
transform 1 0 13328 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104_109
timestamp 1698431365
transform 1 0 13552 0 1 83104
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_104_130
timestamp 1698431365
transform 1 0 15904 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_104_134
timestamp 1698431365
transform 1 0 16352 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_104_138
timestamp 1698431365
transform 1 0 16800 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104_140
timestamp 1698431365
transform 1 0 17024 0 1 83104
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_104_143
timestamp 1698431365
transform 1 0 17360 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_104_254
timestamp 1698431365
transform 1 0 29792 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_104_258
timestamp 1698431365
transform 1 0 30240 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_104_262
timestamp 1698431365
transform 1 0 30688 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_104_266
timestamp 1698431365
transform 1 0 31136 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_104_270
timestamp 1698431365
transform 1 0 31584 0 1 83104
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_104_286
timestamp 1698431365
transform 1 0 33376 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104_290
timestamp 1698431365
transform 1 0 33824 0 1 83104
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_104_313
timestamp 1698431365
transform 1 0 36400 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_104_326
timestamp 1698431365
transform 1 0 37856 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104_330
timestamp 1698431365
transform 1 0 38304 0 1 83104
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_105_2
timestamp 1698431365
transform 1 0 1568 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_105_4
timestamp 1698431365
transform 1 0 1792 0 -1 84672
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_105_28
timestamp 1698431365
transform 1 0 4480 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_105_32
timestamp 1698431365
transform 1 0 4928 0 -1 84672
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_105_64
timestamp 1698431365
transform 1 0 8512 0 -1 84672
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_105_67
timestamp 1698431365
transform 1 0 8848 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_105_69
timestamp 1698431365
transform 1 0 9072 0 -1 84672
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_105_72
timestamp 1698431365
transform 1 0 9408 0 -1 84672
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_105_88
timestamp 1698431365
transform 1 0 11200 0 -1 84672
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_105_96
timestamp 1698431365
transform 1 0 12096 0 -1 84672
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_105_128
timestamp 1698431365
transform 1 0 15680 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_105_132
timestamp 1698431365
transform 1 0 16128 0 -1 84672
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_105_142
timestamp 1698431365
transform 1 0 17248 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_105_144
timestamp 1698431365
transform 1 0 17472 0 -1 84672
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_105_147
timestamp 1698431365
transform 1 0 17808 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_105_151
timestamp 1698431365
transform 1 0 18256 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_105_162
timestamp 1698431365
transform 1 0 19488 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_105_164
timestamp 1698431365
transform 1 0 19712 0 -1 84672
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_105_208
timestamp 1698431365
transform 1 0 24640 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_105_245
timestamp 1698431365
transform 1 0 28784 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_105_255
timestamp 1698431365
transform 1 0 29904 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_105_259
timestamp 1698431365
transform 1 0 30352 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_105_263
timestamp 1698431365
transform 1 0 30800 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_105_267
timestamp 1698431365
transform 1 0 31248 0 -1 84672
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_105_275
timestamp 1698431365
transform 1 0 32144 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_105_279
timestamp 1698431365
transform 1 0 32592 0 -1 84672
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_105_282
timestamp 1698431365
transform 1 0 32928 0 -1 84672
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_106_2
timestamp 1698431365
transform 1 0 1568 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_106_4
timestamp 1698431365
transform 1 0 1792 0 1 84672
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_106_28
timestamp 1698431365
transform 1 0 4480 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_106_32
timestamp 1698431365
transform 1 0 4928 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_106_34
timestamp 1698431365
transform 1 0 5152 0 1 84672
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_106_37
timestamp 1698431365
transform 1 0 5488 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_106_101
timestamp 1698431365
transform 1 0 12656 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_106_107
timestamp 1698431365
transform 1 0 13328 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_106_125
timestamp 1698431365
transform 1 0 15344 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_106_129
timestamp 1698431365
transform 1 0 15792 0 1 84672
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_106_145
timestamp 1698431365
transform 1 0 17584 0 1 84672
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_106_153
timestamp 1698431365
transform 1 0 18480 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_106_157
timestamp 1698431365
transform 1 0 18928 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_106_161
timestamp 1698431365
transform 1 0 19376 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_106_165
timestamp 1698431365
transform 1 0 19824 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_106_177
timestamp 1698431365
transform 1 0 21168 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_106_239
timestamp 1698431365
transform 1 0 28112 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_106_243
timestamp 1698431365
transform 1 0 28560 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_106_257
timestamp 1698431365
transform 1 0 30128 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_106_261
timestamp 1698431365
transform 1 0 30576 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_106_265
timestamp 1698431365
transform 1 0 31024 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_106_283
timestamp 1698431365
transform 1 0 33040 0 1 84672
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_106_312
timestamp 1698431365
transform 1 0 36288 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_106_314
timestamp 1698431365
transform 1 0 36512 0 1 84672
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_106_317
timestamp 1698431365
transform 1 0 36848 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_106_321
timestamp 1698431365
transform 1 0 37296 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_106_325
timestamp 1698431365
transform 1 0 37744 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_106_329
timestamp 1698431365
transform 1 0 38192 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_107_2
timestamp 1698431365
transform 1 0 1568 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_107_4
timestamp 1698431365
transform 1 0 1792 0 -1 86240
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_107_51
timestamp 1698431365
transform 1 0 7056 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_107_55
timestamp 1698431365
transform 1 0 7504 0 -1 86240
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_107_63
timestamp 1698431365
transform 1 0 8400 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_107_67
timestamp 1698431365
transform 1 0 8848 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_107_69
timestamp 1698431365
transform 1 0 9072 0 -1 86240
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_107_72
timestamp 1698431365
transform 1 0 9408 0 -1 86240
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_107_88
timestamp 1698431365
transform 1 0 11200 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_107_94
timestamp 1698431365
transform 1 0 11872 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_107_98
timestamp 1698431365
transform 1 0 12320 0 -1 86240
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_107_106
timestamp 1698431365
transform 1 0 13216 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_107_110
timestamp 1698431365
transform 1 0 13664 0 -1 86240
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_107_119
timestamp 1698431365
transform 1 0 14672 0 -1 86240
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_107_135
timestamp 1698431365
transform 1 0 16464 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_107_139
timestamp 1698431365
transform 1 0 16912 0 -1 86240
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_107_142
timestamp 1698431365
transform 1 0 17248 0 -1 86240
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_107_158
timestamp 1698431365
transform 1 0 19040 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_107_274
timestamp 1698431365
transform 1 0 32032 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_107_290
timestamp 1698431365
transform 1 0 33824 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_107_294
timestamp 1698431365
transform 1 0 34272 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_107_296
timestamp 1698431365
transform 1 0 34496 0 -1 86240
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_107_315
timestamp 1698431365
transform 1 0 36624 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_107_319
timestamp 1698431365
transform 1 0 37072 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_107_323
timestamp 1698431365
transform 1 0 37520 0 -1 86240
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_108_2
timestamp 1698431365
transform 1 0 1568 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_108_4
timestamp 1698431365
transform 1 0 1792 0 1 86240
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_108_28
timestamp 1698431365
transform 1 0 4480 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_108_32
timestamp 1698431365
transform 1 0 4928 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_108_34
timestamp 1698431365
transform 1 0 5152 0 1 86240
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_108_37
timestamp 1698431365
transform 1 0 5488 0 1 86240
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_108_45
timestamp 1698431365
transform 1 0 6384 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_108_49
timestamp 1698431365
transform 1 0 6832 0 1 86240
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_108_73
timestamp 1698431365
transform 1 0 9520 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_108_103
timestamp 1698431365
transform 1 0 12880 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_108_107
timestamp 1698431365
transform 1 0 13328 0 1 86240
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_108_123
timestamp 1698431365
transform 1 0 15120 0 1 86240
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_108_133
timestamp 1698431365
transform 1 0 16240 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_108_149
timestamp 1698431365
transform 1 0 18032 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_108_153
timestamp 1698431365
transform 1 0 18480 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_108_157
timestamp 1698431365
transform 1 0 18928 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_108_161
timestamp 1698431365
transform 1 0 19376 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_108_192
timestamp 1698431365
transform 1 0 22848 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_108_210
timestamp 1698431365
transform 1 0 24864 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_108_243
timestamp 1698431365
transform 1 0 28560 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_108_309
timestamp 1698431365
transform 1 0 35952 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_108_313
timestamp 1698431365
transform 1 0 36400 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_108_317
timestamp 1698431365
transform 1 0 36848 0 1 86240
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_108_325
timestamp 1698431365
transform 1 0 37744 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_108_329
timestamp 1698431365
transform 1 0 38192 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_109_2
timestamp 1698431365
transform 1 0 1568 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_109_4
timestamp 1698431365
transform 1 0 1792 0 -1 87808
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_109_28
timestamp 1698431365
transform 1 0 4480 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_109_32
timestamp 1698431365
transform 1 0 4928 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_109_36
timestamp 1698431365
transform 1 0 5376 0 -1 87808
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_109_44
timestamp 1698431365
transform 1 0 6272 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_109_46
timestamp 1698431365
transform 1 0 6496 0 -1 87808
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_109_114
timestamp 1698431365
transform 1 0 14112 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_109_118
timestamp 1698431365
transform 1 0 14560 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_109_122
timestamp 1698431365
transform 1 0 15008 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_109_139
timestamp 1698431365
transform 1 0 16912 0 -1 87808
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_109_142
timestamp 1698431365
transform 1 0 17248 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_109_159
timestamp 1698431365
transform 1 0 19152 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_109_165
timestamp 1698431365
transform 1 0 19824 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_109_169
timestamp 1698431365
transform 1 0 20272 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_109_188
timestamp 1698431365
transform 1 0 22400 0 -1 87808
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_109_272
timestamp 1698431365
transform 1 0 31808 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_109_276
timestamp 1698431365
transform 1 0 32256 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_109_290
timestamp 1698431365
transform 1 0 33824 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_109_294
timestamp 1698431365
transform 1 0 34272 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_109_327
timestamp 1698431365
transform 1 0 37968 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_110_2
timestamp 1698431365
transform 1 0 1568 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_110_4
timestamp 1698431365
transform 1 0 1792 0 1 87808
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_110_28
timestamp 1698431365
transform 1 0 4480 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_110_32
timestamp 1698431365
transform 1 0 4928 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_110_34
timestamp 1698431365
transform 1 0 5152 0 1 87808
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_110_37
timestamp 1698431365
transform 1 0 5488 0 1 87808
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_110_45
timestamp 1698431365
transform 1 0 6384 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_110_49
timestamp 1698431365
transform 1 0 6832 0 1 87808
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_110_104
timestamp 1698431365
transform 1 0 12992 0 1 87808
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_110_107
timestamp 1698431365
transform 1 0 13328 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_110_167
timestamp 1698431365
transform 1 0 20048 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_110_177
timestamp 1698431365
transform 1 0 21168 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_110_276
timestamp 1698431365
transform 1 0 32256 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_110_280
timestamp 1698431365
transform 1 0 32704 0 1 87808
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_110_296
timestamp 1698431365
transform 1 0 34496 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_110_300
timestamp 1698431365
transform 1 0 34944 0 1 87808
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_110_308
timestamp 1698431365
transform 1 0 35840 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_110_312
timestamp 1698431365
transform 1 0 36288 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_110_314
timestamp 1698431365
transform 1 0 36512 0 1 87808
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_110_317
timestamp 1698431365
transform 1 0 36848 0 1 87808
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_110_325
timestamp 1698431365
transform 1 0 37744 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_110_329
timestamp 1698431365
transform 1 0 38192 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_111_2
timestamp 1698431365
transform 1 0 1568 0 -1 89376
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_111_34
timestamp 1698431365
transform 1 0 5152 0 -1 89376
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_111_42
timestamp 1698431365
transform 1 0 6048 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_111_46
timestamp 1698431365
transform 1 0 6496 0 -1 89376
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_111_72
timestamp 1698431365
transform 1 0 9408 0 -1 89376
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_111_88
timestamp 1698431365
transform 1 0 11200 0 -1 89376
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_111_96
timestamp 1698431365
transform 1 0 12096 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_111_100
timestamp 1698431365
transform 1 0 12544 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_111_102
timestamp 1698431365
transform 1 0 12768 0 -1 89376
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_111_134
timestamp 1698431365
transform 1 0 16352 0 -1 89376
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_111_142
timestamp 1698431365
transform 1 0 17248 0 -1 89376
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_111_180
timestamp 1698431365
transform 1 0 21504 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_111_182
timestamp 1698431365
transform 1 0 21728 0 -1 89376
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_111_200
timestamp 1698431365
transform 1 0 23744 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_111_262
timestamp 1698431365
transform 1 0 30688 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_111_266
timestamp 1698431365
transform 1 0 31136 0 -1 89376
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_111_274
timestamp 1698431365
transform 1 0 32032 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_111_278
timestamp 1698431365
transform 1 0 32480 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_111_282
timestamp 1698431365
transform 1 0 32928 0 -1 89376
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_111_298
timestamp 1698431365
transform 1 0 34720 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_111_302
timestamp 1698431365
transform 1 0 35168 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_111_304
timestamp 1698431365
transform 1 0 35392 0 -1 89376
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_112_2
timestamp 1698431365
transform 1 0 1568 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_112_29
timestamp 1698431365
transform 1 0 4592 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_112_33
timestamp 1698431365
transform 1 0 5040 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_112_37
timestamp 1698431365
transform 1 0 5488 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_112_85
timestamp 1698431365
transform 1 0 10864 0 1 89376
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_112_101
timestamp 1698431365
transform 1 0 12656 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_112_107
timestamp 1698431365
transform 1 0 13328 0 1 89376
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_112_123
timestamp 1698431365
transform 1 0 15120 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_112_127
timestamp 1698431365
transform 1 0 15568 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_112_129
timestamp 1698431365
transform 1 0 15792 0 1 89376
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_112_132
timestamp 1698431365
transform 1 0 16128 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_112_136
timestamp 1698431365
transform 1 0 16576 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_112_140
timestamp 1698431365
transform 1 0 17024 0 1 89376
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_112_143
timestamp 1698431365
transform 1 0 17360 0 1 89376
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_112_159
timestamp 1698431365
transform 1 0 19152 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_112_161
timestamp 1698431365
transform 1 0 19376 0 1 89376
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_112_164
timestamp 1698431365
transform 1 0 19712 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_112_168
timestamp 1698431365
transform 1 0 20160 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_112_172
timestamp 1698431365
transform 1 0 20608 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_112_174
timestamp 1698431365
transform 1 0 20832 0 1 89376
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_112_177
timestamp 1698431365
transform 1 0 21168 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_112_183
timestamp 1698431365
transform 1 0 21840 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_112_187
timestamp 1698431365
transform 1 0 22288 0 1 89376
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_112_209
timestamp 1698431365
transform 1 0 24752 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_112_213
timestamp 1698431365
transform 1 0 25200 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_112_215
timestamp 1698431365
transform 1 0 25424 0 1 89376
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_112_236
timestamp 1698431365
transform 1 0 27776 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_112_240
timestamp 1698431365
transform 1 0 28224 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_112_244
timestamp 1698431365
transform 1 0 28672 0 1 89376
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_112_247
timestamp 1698431365
transform 1 0 29008 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_112_251
timestamp 1698431365
transform 1 0 29456 0 1 89376
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_112_265
timestamp 1698431365
transform 1 0 31024 0 1 89376
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_112_297
timestamp 1698431365
transform 1 0 34608 0 1 89376
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_112_313
timestamp 1698431365
transform 1 0 36400 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_112_317
timestamp 1698431365
transform 1 0 36848 0 1 89376
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_112_325
timestamp 1698431365
transform 1 0 37744 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_112_329
timestamp 1698431365
transform 1 0 38192 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_113_2
timestamp 1698431365
transform 1 0 1568 0 -1 90944
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_113_10
timestamp 1698431365
transform 1 0 2464 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_113_37
timestamp 1698431365
transform 1 0 5488 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_113_41
timestamp 1698431365
transform 1 0 5936 0 -1 90944
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_113_57
timestamp 1698431365
transform 1 0 7728 0 -1 90944
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_113_65
timestamp 1698431365
transform 1 0 8624 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_113_69
timestamp 1698431365
transform 1 0 9072 0 -1 90944
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_113_72
timestamp 1698431365
transform 1 0 9408 0 -1 90944
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_113_88
timestamp 1698431365
transform 1 0 11200 0 -1 90944
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_113_96
timestamp 1698431365
transform 1 0 12096 0 -1 90944
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_113_103
timestamp 1698431365
transform 1 0 12880 0 -1 90944
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_113_135
timestamp 1698431365
transform 1 0 16464 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_113_139
timestamp 1698431365
transform 1 0 16912 0 -1 90944
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_113_142
timestamp 1698431365
transform 1 0 17248 0 -1 90944
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_113_174
timestamp 1698431365
transform 1 0 20832 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_113_178
timestamp 1698431365
transform 1 0 21280 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_113_180
timestamp 1698431365
transform 1 0 21504 0 -1 90944
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_113_183
timestamp 1698431365
transform 1 0 21840 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_113_187
timestamp 1698431365
transform 1 0 22288 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_113_191
timestamp 1698431365
transform 1 0 22736 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_113_195
timestamp 1698431365
transform 1 0 23184 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_113_199
timestamp 1698431365
transform 1 0 23632 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_113_205
timestamp 1698431365
transform 1 0 24304 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_113_207
timestamp 1698431365
transform 1 0 24528 0 -1 90944
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_113_212
timestamp 1698431365
transform 1 0 25088 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_113_222
timestamp 1698431365
transform 1 0 26208 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_113_226
timestamp 1698431365
transform 1 0 26656 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_113_230
timestamp 1698431365
transform 1 0 27104 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_113_234
timestamp 1698431365
transform 1 0 27552 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_113_238
timestamp 1698431365
transform 1 0 28000 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_113_242
timestamp 1698431365
transform 1 0 28448 0 -1 90944
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_113_250
timestamp 1698431365
transform 1 0 29344 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_113_252
timestamp 1698431365
transform 1 0 29568 0 -1 90944
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_113_260
timestamp 1698431365
transform 1 0 30464 0 -1 90944
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_113_276
timestamp 1698431365
transform 1 0 32256 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_113_282
timestamp 1698431365
transform 1 0 32928 0 -1 90944
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_113_314
timestamp 1698431365
transform 1 0 36512 0 -1 90944
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_113_330
timestamp 1698431365
transform 1 0 38304 0 -1 90944
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_114_2
timestamp 1698431365
transform 1 0 1568 0 1 90944
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_114_10
timestamp 1698431365
transform 1 0 2464 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_114_37
timestamp 1698431365
transform 1 0 5488 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_114_41
timestamp 1698431365
transform 1 0 5936 0 1 90944
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_114_57
timestamp 1698431365
transform 1 0 7728 0 1 90944
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_114_65
timestamp 1698431365
transform 1 0 8624 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_114_69
timestamp 1698431365
transform 1 0 9072 0 1 90944
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_114_85
timestamp 1698431365
transform 1 0 10864 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_114_89
timestamp 1698431365
transform 1 0 11312 0 1 90944
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_114_102
timestamp 1698431365
transform 1 0 12768 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_114_104
timestamp 1698431365
transform 1 0 12992 0 1 90944
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_114_113
timestamp 1698431365
transform 1 0 14000 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_114_117
timestamp 1698431365
transform 1 0 14448 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_114_121
timestamp 1698431365
transform 1 0 14896 0 1 90944
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_114_153
timestamp 1698431365
transform 1 0 18480 0 1 90944
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_114_169
timestamp 1698431365
transform 1 0 20272 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_114_173
timestamp 1698431365
transform 1 0 20720 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_114_177
timestamp 1698431365
transform 1 0 21168 0 1 90944
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_114_185
timestamp 1698431365
transform 1 0 22064 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_114_239
timestamp 1698431365
transform 1 0 28112 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_114_243
timestamp 1698431365
transform 1 0 28560 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_114_247
timestamp 1698431365
transform 1 0 29008 0 1 90944
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_114_263
timestamp 1698431365
transform 1 0 30800 0 1 90944
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_114_271
timestamp 1698431365
transform 1 0 31696 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_114_275
timestamp 1698431365
transform 1 0 32144 0 1 90944
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_114_299
timestamp 1698431365
transform 1 0 34832 0 1 90944
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_114_317
timestamp 1698431365
transform 1 0 36848 0 1 90944
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_114_325
timestamp 1698431365
transform 1 0 37744 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_114_329
timestamp 1698431365
transform 1 0 38192 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_115_2
timestamp 1698431365
transform 1 0 1568 0 -1 92512
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_115_10
timestamp 1698431365
transform 1 0 2464 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_115_36
timestamp 1698431365
transform 1 0 5376 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_115_40
timestamp 1698431365
transform 1 0 5824 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_115_67
timestamp 1698431365
transform 1 0 8848 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_115_69
timestamp 1698431365
transform 1 0 9072 0 -1 92512
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_115_72
timestamp 1698431365
transform 1 0 9408 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_115_121
timestamp 1698431365
transform 1 0 14896 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_115_125
timestamp 1698431365
transform 1 0 15344 0 -1 92512
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_115_133
timestamp 1698431365
transform 1 0 16240 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_115_137
timestamp 1698431365
transform 1 0 16688 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_115_139
timestamp 1698431365
transform 1 0 16912 0 -1 92512
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_115_142
timestamp 1698431365
transform 1 0 17248 0 -1 92512
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_115_158
timestamp 1698431365
transform 1 0 19040 0 -1 92512
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_115_166
timestamp 1698431365
transform 1 0 19936 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_115_170
timestamp 1698431365
transform 1 0 20384 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_115_185
timestamp 1698431365
transform 1 0 22064 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_115_189
timestamp 1698431365
transform 1 0 22512 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_115_193
timestamp 1698431365
transform 1 0 22960 0 -1 92512
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_115_198
timestamp 1698431365
transform 1 0 23520 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_115_202
timestamp 1698431365
transform 1 0 23968 0 -1 92512
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_115_205
timestamp 1698431365
transform 1 0 24304 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_115_207
timestamp 1698431365
transform 1 0 24528 0 -1 92512
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_115_229
timestamp 1698431365
transform 1 0 26992 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_115_239
timestamp 1698431365
transform 1 0 28112 0 -1 92512
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_115_271
timestamp 1698431365
transform 1 0 31696 0 -1 92512
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_115_279
timestamp 1698431365
transform 1 0 32592 0 -1 92512
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_115_305
timestamp 1698431365
transform 1 0 35504 0 -1 92512
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_115_321
timestamp 1698431365
transform 1 0 37296 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_116_2
timestamp 1698431365
transform 1 0 1568 0 1 92512
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_116_10
timestamp 1698431365
transform 1 0 2464 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_116_37
timestamp 1698431365
transform 1 0 5488 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_116_41
timestamp 1698431365
transform 1 0 5936 0 1 92512
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_116_72
timestamp 1698431365
transform 1 0 9408 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_116_76
timestamp 1698431365
transform 1 0 9856 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_116_121
timestamp 1698431365
transform 1 0 14896 0 1 92512
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_116_137
timestamp 1698431365
transform 1 0 16688 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_116_152
timestamp 1698431365
transform 1 0 18368 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_116_156
timestamp 1698431365
transform 1 0 18816 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_116_158
timestamp 1698431365
transform 1 0 19040 0 1 92512
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_116_163
timestamp 1698431365
transform 1 0 19600 0 1 92512
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_116_171
timestamp 1698431365
transform 1 0 20496 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_116_200
timestamp 1698431365
transform 1 0 23744 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_116_210
timestamp 1698431365
transform 1 0 24864 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_116_214
timestamp 1698431365
transform 1 0 25312 0 1 92512
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_116_219
timestamp 1698431365
transform 1 0 25872 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_116_223
timestamp 1698431365
transform 1 0 26320 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_116_239
timestamp 1698431365
transform 1 0 28112 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_116_243
timestamp 1698431365
transform 1 0 28560 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_116_293
timestamp 1698431365
transform 1 0 34160 0 1 92512
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_116_309
timestamp 1698431365
transform 1 0 35952 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_116_313
timestamp 1698431365
transform 1 0 36400 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_116_317
timestamp 1698431365
transform 1 0 36848 0 1 92512
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_116_325
timestamp 1698431365
transform 1 0 37744 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_116_329
timestamp 1698431365
transform 1 0 38192 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_117_2
timestamp 1698431365
transform 1 0 1568 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_117_27
timestamp 1698431365
transform 1 0 4368 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_117_31
timestamp 1698431365
transform 1 0 4816 0 -1 94080
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_117_72
timestamp 1698431365
transform 1 0 9408 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_117_76
timestamp 1698431365
transform 1 0 9856 0 -1 94080
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_117_109
timestamp 1698431365
transform 1 0 13552 0 -1 94080
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_117_125
timestamp 1698431365
transform 1 0 15344 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_117_129
timestamp 1698431365
transform 1 0 15792 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_117_131
timestamp 1698431365
transform 1 0 16016 0 -1 94080
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_117_165
timestamp 1698431365
transform 1 0 19824 0 -1 94080
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_117_235
timestamp 1698431365
transform 1 0 27664 0 -1 94080
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_117_266
timestamp 1698431365
transform 1 0 31136 0 -1 94080
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_117_274
timestamp 1698431365
transform 1 0 32032 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_117_278
timestamp 1698431365
transform 1 0 32480 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_117_305
timestamp 1698431365
transform 1 0 35504 0 -1 94080
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_117_321
timestamp 1698431365
transform 1 0 37296 0 -1 94080
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_117_329
timestamp 1698431365
transform 1 0 38192 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_118_6
timestamp 1698431365
transform 1 0 2016 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_118_10
timestamp 1698431365
transform 1 0 2464 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_118_37
timestamp 1698431365
transform 1 0 5488 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_118_41
timestamp 1698431365
transform 1 0 5936 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_118_43
timestamp 1698431365
transform 1 0 6160 0 1 94080
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_118_46
timestamp 1698431365
transform 1 0 6496 0 1 94080
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_118_78
timestamp 1698431365
transform 1 0 10080 0 1 94080
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_118_94
timestamp 1698431365
transform 1 0 11872 0 1 94080
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_118_102
timestamp 1698431365
transform 1 0 12768 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_118_104
timestamp 1698431365
transform 1 0 12992 0 1 94080
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_118_107
timestamp 1698431365
transform 1 0 13328 0 1 94080
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_118_123
timestamp 1698431365
transform 1 0 15120 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_118_125
timestamp 1698431365
transform 1 0 15344 0 1 94080
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_118_140
timestamp 1698431365
transform 1 0 17024 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_118_144
timestamp 1698431365
transform 1 0 17472 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_118_148
timestamp 1698431365
transform 1 0 17920 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_118_193
timestamp 1698431365
transform 1 0 22960 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_118_197
timestamp 1698431365
transform 1 0 23408 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_118_201
timestamp 1698431365
transform 1 0 23856 0 1 94080
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_118_220
timestamp 1698431365
transform 1 0 25984 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_118_270
timestamp 1698431365
transform 1 0 31584 0 1 94080
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_118_278
timestamp 1698431365
transform 1 0 32480 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_118_303
timestamp 1698431365
transform 1 0 35280 0 1 94080
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_118_311
timestamp 1698431365
transform 1 0 36176 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_118_317
timestamp 1698431365
transform 1 0 36848 0 1 94080
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_118_325
timestamp 1698431365
transform 1 0 37744 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_118_329
timestamp 1698431365
transform 1 0 38192 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_119_2
timestamp 1698431365
transform 1 0 1568 0 -1 95648
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_119_18
timestamp 1698431365
transform 1 0 3360 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_119_20
timestamp 1698431365
transform 1 0 3584 0 -1 95648
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_119_44
timestamp 1698431365
transform 1 0 6272 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_119_46
timestamp 1698431365
transform 1 0 6496 0 -1 95648
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_119_72
timestamp 1698431365
transform 1 0 9408 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_119_76
timestamp 1698431365
transform 1 0 9856 0 -1 95648
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_119_92
timestamp 1698431365
transform 1 0 11648 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_119_96
timestamp 1698431365
transform 1 0 12096 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_119_121
timestamp 1698431365
transform 1 0 14896 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_119_125
timestamp 1698431365
transform 1 0 15344 0 -1 95648
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_119_133
timestamp 1698431365
transform 1 0 16240 0 -1 95648
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_119_188
timestamp 1698431365
transform 1 0 22400 0 -1 95648
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_119_196
timestamp 1698431365
transform 1 0 23296 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_119_200
timestamp 1698431365
transform 1 0 23744 0 -1 95648
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_119_235
timestamp 1698431365
transform 1 0 27664 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_119_237
timestamp 1698431365
transform 1 0 27888 0 -1 95648
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_119_261
timestamp 1698431365
transform 1 0 30576 0 -1 95648
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_119_277
timestamp 1698431365
transform 1 0 32368 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_119_279
timestamp 1698431365
transform 1 0 32592 0 -1 95648
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_119_328
timestamp 1698431365
transform 1 0 38080 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_119_330
timestamp 1698431365
transform 1 0 38304 0 -1 95648
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_120_2
timestamp 1698431365
transform 1 0 1568 0 1 95648
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_120_10
timestamp 1698431365
transform 1 0 2464 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_120_37
timestamp 1698431365
transform 1 0 5488 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_120_41
timestamp 1698431365
transform 1 0 5936 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_120_45
timestamp 1698431365
transform 1 0 6384 0 1 95648
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_120_93
timestamp 1698431365
transform 1 0 11760 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_120_97
timestamp 1698431365
transform 1 0 12208 0 1 95648
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_120_130
timestamp 1698431365
transform 1 0 15904 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_120_134
timestamp 1698431365
transform 1 0 16352 0 1 95648
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_120_165
timestamp 1698431365
transform 1 0 19824 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_120_169
timestamp 1698431365
transform 1 0 20272 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_120_206
timestamp 1698431365
transform 1 0 24416 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_120_222
timestamp 1698431365
transform 1 0 26208 0 1 95648
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_120_229
timestamp 1698431365
transform 1 0 26992 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_120_233
timestamp 1698431365
transform 1 0 27440 0 1 95648
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_120_241
timestamp 1698431365
transform 1 0 28336 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_120_270
timestamp 1698431365
transform 1 0 31584 0 1 95648
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_120_278
timestamp 1698431365
transform 1 0 32480 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_120_303
timestamp 1698431365
transform 1 0 35280 0 1 95648
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_120_311
timestamp 1698431365
transform 1 0 36176 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_120_317
timestamp 1698431365
transform 1 0 36848 0 1 95648
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_120_325
timestamp 1698431365
transform 1 0 37744 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_120_329
timestamp 1698431365
transform 1 0 38192 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_121_2
timestamp 1698431365
transform 1 0 1568 0 -1 97216
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_121_34
timestamp 1698431365
transform 1 0 5152 0 -1 97216
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_121_42
timestamp 1698431365
transform 1 0 6048 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_121_46
timestamp 1698431365
transform 1 0 6496 0 -1 97216
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_121_72
timestamp 1698431365
transform 1 0 9408 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_121_76
timestamp 1698431365
transform 1 0 9856 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_121_80
timestamp 1698431365
transform 1 0 10304 0 -1 97216
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_121_96
timestamp 1698431365
transform 1 0 12096 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_121_121
timestamp 1698431365
transform 1 0 14896 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_121_125
timestamp 1698431365
transform 1 0 15344 0 -1 97216
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_121_133
timestamp 1698431365
transform 1 0 16240 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_121_137
timestamp 1698431365
transform 1 0 16688 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_121_139
timestamp 1698431365
transform 1 0 16912 0 -1 97216
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_121_142
timestamp 1698431365
transform 1 0 17248 0 -1 97216
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_121_206
timestamp 1698431365
transform 1 0 24416 0 -1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_121_212
timestamp 1698431365
transform 1 0 25088 0 -1 97216
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_121_244
timestamp 1698431365
transform 1 0 28672 0 -1 97216
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_121_252
timestamp 1698431365
transform 1 0 29568 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_121_254
timestamp 1698431365
transform 1 0 29792 0 -1 97216
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_121_278
timestamp 1698431365
transform 1 0 32480 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_121_305
timestamp 1698431365
transform 1 0 35504 0 -1 97216
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_121_321
timestamp 1698431365
transform 1 0 37296 0 -1 97216
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_121_329
timestamp 1698431365
transform 1 0 38192 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_122_6
timestamp 1698431365
transform 1 0 2016 0 1 97216
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_122_22
timestamp 1698431365
transform 1 0 3808 0 1 97216
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_122_27
timestamp 1698431365
transform 1 0 4368 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_122_31
timestamp 1698431365
transform 1 0 4816 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_122_33
timestamp 1698431365
transform 1 0 5040 0 1 97216
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_122_36
timestamp 1698431365
transform 1 0 5376 0 1 97216
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_122_44
timestamp 1698431365
transform 1 0 6272 0 1 97216
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_122_49
timestamp 1698431365
transform 1 0 6832 0 1 97216
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_122_65
timestamp 1698431365
transform 1 0 8624 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_122_67
timestamp 1698431365
transform 1 0 8848 0 1 97216
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_122_74
timestamp 1698431365
transform 1 0 9632 0 1 97216
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_122_82
timestamp 1698431365
transform 1 0 10528 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_122_86
timestamp 1698431365
transform 1 0 10976 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_122_88
timestamp 1698431365
transform 1 0 11200 0 1 97216
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_122_93
timestamp 1698431365
transform 1 0 11760 0 1 97216
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_122_101
timestamp 1698431365
transform 1 0 12656 0 1 97216
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_122_131
timestamp 1698431365
transform 1 0 16016 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_122_135
timestamp 1698431365
transform 1 0 16464 0 1 97216
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_122_142
timestamp 1698431365
transform 1 0 17248 0 1 97216
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_122_150
timestamp 1698431365
transform 1 0 18144 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_122_154
timestamp 1698431365
transform 1 0 18592 0 1 97216
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_122_159
timestamp 1698431365
transform 1 0 19152 0 1 97216
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_122_167
timestamp 1698431365
transform 1 0 20048 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_122_169
timestamp 1698431365
transform 1 0 20272 0 1 97216
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_122_172
timestamp 1698431365
transform 1 0 20608 0 1 97216
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_122_206
timestamp 1698431365
transform 1 0 24416 0 1 97216
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_122_240
timestamp 1698431365
transform 1 0 28224 0 1 97216
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_122_274
timestamp 1698431365
transform 1 0 32032 0 1 97216
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_122_308
timestamp 1698431365
transform 1 0 35840 0 1 97216
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_122_324
timestamp 1698431365
transform 1 0 37632 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_122_328
timestamp 1698431365
transform 1 0 38080 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_122_330
timestamp 1698431365
transform 1 0 38304 0 1 97216
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698431365
transform -1 0 37184 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform -1 0 27888 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698431365
transform 1 0 26432 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698431365
transform 1 0 25760 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform 1 0 25088 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform 1 0 24416 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698431365
transform 1 0 22736 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1698431365
transform 1 0 21840 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1698431365
transform 1 0 20944 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1698431365
transform 1 0 19712 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1698431365
transform 1 0 19040 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1698431365
transform -1 0 36512 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1698431365
transform 1 0 18256 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input14
timestamp 1698431365
transform 1 0 17360 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input15
timestamp 1698431365
transform -1 0 17920 0 -1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input16
timestamp 1698431365
transform 1 0 15232 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input17
timestamp 1698431365
transform 1 0 14560 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input18
timestamp 1698431365
transform 1 0 13776 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input19
timestamp 1698431365
transform 1 0 12096 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input20
timestamp 1698431365
transform 1 0 11424 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input21
timestamp 1698431365
transform -1 0 11424 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input22
timestamp 1698431365
transform -1 0 10752 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input23
timestamp 1698431365
transform -1 0 35056 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input24
timestamp 1698431365
transform 1 0 9296 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input25
timestamp 1698431365
transform 1 0 8288 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input26
timestamp 1698431365
transform 1 0 33488 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input27
timestamp 1698431365
transform 1 0 32704 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input28
timestamp 1698431365
transform 1 0 32032 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input29
timestamp 1698431365
transform 1 0 30800 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input30
timestamp 1698431365
transform 1 0 29904 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input31
timestamp 1698431365
transform -1 0 29680 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input32
timestamp 1698431365
transform 1 0 28224 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input33
timestamp 1698431365
transform 1 0 7504 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input34
timestamp 1698431365
transform 1 0 6608 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input35
timestamp 1698431365
transform 1 0 5712 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  input36
timestamp 1698431365
transform -1 0 38416 0 -1 9408
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input37
timestamp 1698431365
transform -1 0 38416 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  input38
timestamp 1698431365
transform -1 0 38416 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input39
timestamp 1698431365
transform -1 0 38416 0 -1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input40
timestamp 1698431365
transform -1 0 38416 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input41
timestamp 1698431365
transform -1 0 38416 0 -1 92512
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input42
timestamp 1698431365
transform 1 0 3920 0 1 1568
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_123 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 38640 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_124
timestamp 1698431365
transform 1 0 1344 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 38640 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_125
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 38640 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_126
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 38640 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_127
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 38640 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_128
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 38640 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_129
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 38640 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_130
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 38640 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_131
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 38640 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_132
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 38640 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_133
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 38640 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_134
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 38640 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_135
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 38640 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_136
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 38640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_137
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 38640 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_138
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 38640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_139
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 38640 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_140
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 38640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_141
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 38640 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_142
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 38640 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_143
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 38640 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_144
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 38640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_145
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 38640 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_146
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 38640 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_147
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 38640 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_148
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 38640 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_149
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 38640 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_150
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 38640 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_151
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 38640 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_152
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 38640 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_153
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 38640 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_154
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 38640 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_155
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 38640 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_156
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 38640 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_157
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 38640 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_158
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 38640 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_159
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 38640 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_160
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 38640 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_161
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 38640 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_162
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 38640 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_163
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 38640 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_164
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 38640 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_165
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 38640 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_166
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 38640 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_167
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 38640 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_168
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 38640 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_169
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 38640 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_170
timestamp 1698431365
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 38640 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_171
timestamp 1698431365
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 38640 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_172
timestamp 1698431365
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 38640 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_173
timestamp 1698431365
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698431365
transform -1 0 38640 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_174
timestamp 1698431365
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698431365
transform -1 0 38640 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_175
timestamp 1698431365
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1698431365
transform -1 0 38640 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_176
timestamp 1698431365
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1698431365
transform -1 0 38640 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_177
timestamp 1698431365
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1698431365
transform -1 0 38640 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Left_178
timestamp 1698431365
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Right_55
timestamp 1698431365
transform -1 0 38640 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Left_179
timestamp 1698431365
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Right_56
timestamp 1698431365
transform -1 0 38640 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Left_180
timestamp 1698431365
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Right_57
timestamp 1698431365
transform -1 0 38640 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Left_181
timestamp 1698431365
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Right_58
timestamp 1698431365
transform -1 0 38640 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Left_182
timestamp 1698431365
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Right_59
timestamp 1698431365
transform -1 0 38640 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Left_183
timestamp 1698431365
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Right_60
timestamp 1698431365
transform -1 0 38640 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Left_184
timestamp 1698431365
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Right_61
timestamp 1698431365
transform -1 0 38640 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Left_185
timestamp 1698431365
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Right_62
timestamp 1698431365
transform -1 0 38640 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Left_186
timestamp 1698431365
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Right_63
timestamp 1698431365
transform -1 0 38640 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Left_187
timestamp 1698431365
transform 1 0 1344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Right_64
timestamp 1698431365
transform -1 0 38640 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Left_188
timestamp 1698431365
transform 1 0 1344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Right_65
timestamp 1698431365
transform -1 0 38640 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Left_189
timestamp 1698431365
transform 1 0 1344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Right_66
timestamp 1698431365
transform -1 0 38640 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Left_190
timestamp 1698431365
transform 1 0 1344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Right_67
timestamp 1698431365
transform -1 0 38640 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_68_Left_191
timestamp 1698431365
transform 1 0 1344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_68_Right_68
timestamp 1698431365
transform -1 0 38640 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_69_Left_192
timestamp 1698431365
transform 1 0 1344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_69_Right_69
timestamp 1698431365
transform -1 0 38640 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_70_Left_193
timestamp 1698431365
transform 1 0 1344 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_70_Right_70
timestamp 1698431365
transform -1 0 38640 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_71_Left_194
timestamp 1698431365
transform 1 0 1344 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_71_Right_71
timestamp 1698431365
transform -1 0 38640 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_72_Left_195
timestamp 1698431365
transform 1 0 1344 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_72_Right_72
timestamp 1698431365
transform -1 0 38640 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_73_Left_196
timestamp 1698431365
transform 1 0 1344 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_73_Right_73
timestamp 1698431365
transform -1 0 38640 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_74_Left_197
timestamp 1698431365
transform 1 0 1344 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_74_Right_74
timestamp 1698431365
transform -1 0 38640 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_75_Left_198
timestamp 1698431365
transform 1 0 1344 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_75_Right_75
timestamp 1698431365
transform -1 0 38640 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_76_Left_199
timestamp 1698431365
transform 1 0 1344 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_76_Right_76
timestamp 1698431365
transform -1 0 38640 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_77_Left_200
timestamp 1698431365
transform 1 0 1344 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_77_Right_77
timestamp 1698431365
transform -1 0 38640 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_78_Left_201
timestamp 1698431365
transform 1 0 1344 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_78_Right_78
timestamp 1698431365
transform -1 0 38640 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_79_Left_202
timestamp 1698431365
transform 1 0 1344 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_79_Right_79
timestamp 1698431365
transform -1 0 38640 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_80_Left_203
timestamp 1698431365
transform 1 0 1344 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_80_Right_80
timestamp 1698431365
transform -1 0 38640 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_81_Left_204
timestamp 1698431365
transform 1 0 1344 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_81_Right_81
timestamp 1698431365
transform -1 0 38640 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_82_Left_205
timestamp 1698431365
transform 1 0 1344 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_82_Right_82
timestamp 1698431365
transform -1 0 38640 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_83_Left_206
timestamp 1698431365
transform 1 0 1344 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_83_Right_83
timestamp 1698431365
transform -1 0 38640 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_84_Left_207
timestamp 1698431365
transform 1 0 1344 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_84_Right_84
timestamp 1698431365
transform -1 0 38640 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_85_Left_208
timestamp 1698431365
transform 1 0 1344 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_85_Right_85
timestamp 1698431365
transform -1 0 38640 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_86_Left_209
timestamp 1698431365
transform 1 0 1344 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_86_Right_86
timestamp 1698431365
transform -1 0 38640 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_87_Left_210
timestamp 1698431365
transform 1 0 1344 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_87_Right_87
timestamp 1698431365
transform -1 0 38640 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_88_Left_211
timestamp 1698431365
transform 1 0 1344 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_88_Right_88
timestamp 1698431365
transform -1 0 38640 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_89_Left_212
timestamp 1698431365
transform 1 0 1344 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_89_Right_89
timestamp 1698431365
transform -1 0 38640 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_90_Left_213
timestamp 1698431365
transform 1 0 1344 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_90_Right_90
timestamp 1698431365
transform -1 0 38640 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_91_Left_214
timestamp 1698431365
transform 1 0 1344 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_91_Right_91
timestamp 1698431365
transform -1 0 38640 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_92_Left_215
timestamp 1698431365
transform 1 0 1344 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_92_Right_92
timestamp 1698431365
transform -1 0 38640 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_93_Left_216
timestamp 1698431365
transform 1 0 1344 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_93_Right_93
timestamp 1698431365
transform -1 0 38640 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_94_Left_217
timestamp 1698431365
transform 1 0 1344 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_94_Right_94
timestamp 1698431365
transform -1 0 38640 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_95_Left_218
timestamp 1698431365
transform 1 0 1344 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_95_Right_95
timestamp 1698431365
transform -1 0 38640 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_96_Left_219
timestamp 1698431365
transform 1 0 1344 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_96_Right_96
timestamp 1698431365
transform -1 0 38640 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_97_Left_220
timestamp 1698431365
transform 1 0 1344 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_97_Right_97
timestamp 1698431365
transform -1 0 38640 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_98_Left_221
timestamp 1698431365
transform 1 0 1344 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_98_Right_98
timestamp 1698431365
transform -1 0 38640 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_99_Left_222
timestamp 1698431365
transform 1 0 1344 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_99_Right_99
timestamp 1698431365
transform -1 0 38640 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_100_Left_223
timestamp 1698431365
transform 1 0 1344 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_100_Right_100
timestamp 1698431365
transform -1 0 38640 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_101_Left_224
timestamp 1698431365
transform 1 0 1344 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_101_Right_101
timestamp 1698431365
transform -1 0 38640 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_102_Left_225
timestamp 1698431365
transform 1 0 1344 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_102_Right_102
timestamp 1698431365
transform -1 0 38640 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_103_Left_226
timestamp 1698431365
transform 1 0 1344 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_103_Right_103
timestamp 1698431365
transform -1 0 38640 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_104_Left_227
timestamp 1698431365
transform 1 0 1344 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_104_Right_104
timestamp 1698431365
transform -1 0 38640 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_105_Left_228
timestamp 1698431365
transform 1 0 1344 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_105_Right_105
timestamp 1698431365
transform -1 0 38640 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_106_Left_229
timestamp 1698431365
transform 1 0 1344 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_106_Right_106
timestamp 1698431365
transform -1 0 38640 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_107_Left_230
timestamp 1698431365
transform 1 0 1344 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_107_Right_107
timestamp 1698431365
transform -1 0 38640 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_108_Left_231
timestamp 1698431365
transform 1 0 1344 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_108_Right_108
timestamp 1698431365
transform -1 0 38640 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_109_Left_232
timestamp 1698431365
transform 1 0 1344 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_109_Right_109
timestamp 1698431365
transform -1 0 38640 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_110_Left_233
timestamp 1698431365
transform 1 0 1344 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_110_Right_110
timestamp 1698431365
transform -1 0 38640 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_111_Left_234
timestamp 1698431365
transform 1 0 1344 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_111_Right_111
timestamp 1698431365
transform -1 0 38640 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_112_Left_235
timestamp 1698431365
transform 1 0 1344 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_112_Right_112
timestamp 1698431365
transform -1 0 38640 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_113_Left_236
timestamp 1698431365
transform 1 0 1344 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_113_Right_113
timestamp 1698431365
transform -1 0 38640 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_114_Left_237
timestamp 1698431365
transform 1 0 1344 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_114_Right_114
timestamp 1698431365
transform -1 0 38640 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_115_Left_238
timestamp 1698431365
transform 1 0 1344 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_115_Right_115
timestamp 1698431365
transform -1 0 38640 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_116_Left_239
timestamp 1698431365
transform 1 0 1344 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_116_Right_116
timestamp 1698431365
transform -1 0 38640 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_117_Left_240
timestamp 1698431365
transform 1 0 1344 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_117_Right_117
timestamp 1698431365
transform -1 0 38640 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_118_Left_241
timestamp 1698431365
transform 1 0 1344 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_118_Right_118
timestamp 1698431365
transform -1 0 38640 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_119_Left_242
timestamp 1698431365
transform 1 0 1344 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_119_Right_119
timestamp 1698431365
transform -1 0 38640 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_120_Left_243
timestamp 1698431365
transform 1 0 1344 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_120_Right_120
timestamp 1698431365
transform -1 0 38640 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_121_Left_244
timestamp 1698431365
transform 1 0 1344 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_121_Right_121
timestamp 1698431365
transform -1 0 38640 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_122_Left_245
timestamp 1698431365
transform 1 0 1344 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_122_Right_122
timestamp 1698431365
transform -1 0 38640 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  seg1._26_
timestamp 1698431365
transform 1 0 34496 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  seg1._27_
timestamp 1698431365
transform 1 0 36960 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  seg1._28_
timestamp 1698431365
transform 1 0 36848 0 1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  seg1._29_
timestamp 1698431365
transform 1 0 36176 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  seg1._30_
timestamp 1698431365
transform 1 0 34272 0 -1 78400
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  seg1._31_
timestamp 1698431365
transform 1 0 37744 0 1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  seg1._32_
timestamp 1698431365
transform 1 0 36512 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  seg1._33_
timestamp 1698431365
transform -1 0 36288 0 1 78400
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  seg1._34_
timestamp 1698431365
transform -1 0 36176 0 1 76832
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  seg1._35_
timestamp 1698431365
transform 1 0 35056 0 -1 76832
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  seg1._36_
timestamp 1698431365
transform -1 0 35616 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  seg1._37_
timestamp 1698431365
transform -1 0 34272 0 -1 75264
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  seg1._38_
timestamp 1698431365
transform -1 0 36512 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  seg1._39_
timestamp 1698431365
transform 1 0 35616 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  seg1._40_
timestamp 1698431365
transform 1 0 35504 0 1 73696
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  seg1._41_
timestamp 1698431365
transform 1 0 33376 0 1 75264
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  seg1._42_
timestamp 1698431365
transform -1 0 38192 0 -1 76832
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  seg1._43_
timestamp 1698431365
transform -1 0 33824 0 1 76832
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  seg1._44_
timestamp 1698431365
transform 1 0 33152 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  seg1._45_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 35504 0 1 75264
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  seg1._46_
timestamp 1698431365
transform -1 0 36512 0 1 75264
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  seg1._47_
timestamp 1698431365
transform -1 0 34944 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  seg1._48_
timestamp 1698431365
transform -1 0 33600 0 -1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  seg1._49_
timestamp 1698431365
transform 1 0 36848 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  seg1._50_
timestamp 1698431365
transform 1 0 32144 0 -1 76832
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  seg1._51_
timestamp 1698431365
transform 1 0 34944 0 -1 78400
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  seg1._52_
timestamp 1698431365
transform -1 0 35168 0 1 78400
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  seg1._53_
timestamp 1698431365
transform -1 0 35504 0 1 73696
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  seg1._54_
timestamp 1698431365
transform -1 0 35168 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  seg1._55_
timestamp 1698431365
transform -1 0 34160 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  seg1._56_
timestamp 1698431365
transform 1 0 36736 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  seg1._57_
timestamp 1698431365
transform -1 0 36960 0 -1 78400
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  seg1._58_
timestamp 1698431365
transform 1 0 34048 0 1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_246 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_247
timestamp 1698431365
transform 1 0 8960 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_248
timestamp 1698431365
transform 1 0 12768 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_249
timestamp 1698431365
transform 1 0 16576 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_250
timestamp 1698431365
transform 1 0 20384 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_251
timestamp 1698431365
transform 1 0 24192 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_252
timestamp 1698431365
transform 1 0 28000 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_253
timestamp 1698431365
transform 1 0 31808 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_254
timestamp 1698431365
transform 1 0 35616 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_255
timestamp 1698431365
transform 1 0 9184 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_256
timestamp 1698431365
transform 1 0 17024 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_257
timestamp 1698431365
transform 1 0 24864 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_258
timestamp 1698431365
transform 1 0 32704 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_259
timestamp 1698431365
transform 1 0 5264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_260
timestamp 1698431365
transform 1 0 13104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_261
timestamp 1698431365
transform 1 0 20944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_262
timestamp 1698431365
transform 1 0 28784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_263
timestamp 1698431365
transform 1 0 36624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_264
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_265
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_266
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_267
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_268
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_269
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_270
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_271
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_272
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_273
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_274
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_275
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_276
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_277
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_278
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_279
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_280
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_281
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_282
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_283
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_284
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_285
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_286
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_287
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_288
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_289
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_290
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_291
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_292
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_293
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_294
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_295
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_296
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_297
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_298
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_299
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_300
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_301
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_302
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_303
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_304
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_305
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_306
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_307
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_308
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_309
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_310
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_311
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_312
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_313
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_314
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_315
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_316
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_317
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_318
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_319
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_320
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_321
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_322
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_323
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_324
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_325
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_326
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_327
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_328
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_329
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_330
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_331
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_332
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_333
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_334
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_335
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_336
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_337
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_338
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_339
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_340
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_341
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_342
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_343
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_344
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_345
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_346
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_347
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_348
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_349
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_350
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_351
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_352
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_353
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_354
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_355
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_356
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_357
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_358
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_359
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_360
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_361
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_362
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_363
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_364
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_365
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_366
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_367
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_368
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_369
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_370
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_371
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_372
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_373
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_374
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_375
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_376
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_377
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_378
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_379
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_380
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_381
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_382
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_383
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_384
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_385
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_386
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_387
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_388
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_389
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_390
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_391
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_392
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_393
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_394
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_395
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_396
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_397
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_398
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_399
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_400
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_401
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_402
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_403
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_404
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_405
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_406
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_407
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_408
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_409
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_410
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_411
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_412
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_413
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_414
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_415
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_416
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_417
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_418
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_419
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_420
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_421
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_422
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_423
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_424
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_425
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_426
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_427
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_428
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_429
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_430
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_431
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_432
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_433
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_434
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_435
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_436
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_437
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_438
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_439
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_440
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_441
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_442
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_443
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_444
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_445
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_446
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_447
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_448
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_449
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_450
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_451
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_452
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_453
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_454
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_455
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_456
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_457
timestamp 1698431365
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_458
timestamp 1698431365
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_459
timestamp 1698431365
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_460
timestamp 1698431365
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_461
timestamp 1698431365
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_462
timestamp 1698431365
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_463
timestamp 1698431365
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_464
timestamp 1698431365
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_465
timestamp 1698431365
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_466
timestamp 1698431365
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_467
timestamp 1698431365
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_468
timestamp 1698431365
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_469
timestamp 1698431365
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_470
timestamp 1698431365
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_471
timestamp 1698431365
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_472
timestamp 1698431365
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_473
timestamp 1698431365
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_474
timestamp 1698431365
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_475
timestamp 1698431365
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_476
timestamp 1698431365
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_477
timestamp 1698431365
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_478
timestamp 1698431365
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_479
timestamp 1698431365
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_480
timestamp 1698431365
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_481
timestamp 1698431365
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_482
timestamp 1698431365
transform 1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_483
timestamp 1698431365
transform 1 0 32704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_484
timestamp 1698431365
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_485
timestamp 1698431365
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_486
timestamp 1698431365
transform 1 0 20944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_487
timestamp 1698431365
transform 1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_488
timestamp 1698431365
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_489
timestamp 1698431365
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_490
timestamp 1698431365
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_491
timestamp 1698431365
transform 1 0 24864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_492
timestamp 1698431365
transform 1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_493
timestamp 1698431365
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_494
timestamp 1698431365
transform 1 0 13104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_495
timestamp 1698431365
transform 1 0 20944 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_496
timestamp 1698431365
transform 1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_497
timestamp 1698431365
transform 1 0 36624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_498
timestamp 1698431365
transform 1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_499
timestamp 1698431365
transform 1 0 17024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_500
timestamp 1698431365
transform 1 0 24864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_501
timestamp 1698431365
transform 1 0 32704 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_502
timestamp 1698431365
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_503
timestamp 1698431365
transform 1 0 13104 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_504
timestamp 1698431365
transform 1 0 20944 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_505
timestamp 1698431365
transform 1 0 28784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_506
timestamp 1698431365
transform 1 0 36624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_507
timestamp 1698431365
transform 1 0 9184 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_508
timestamp 1698431365
transform 1 0 17024 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_509
timestamp 1698431365
transform 1 0 24864 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_510
timestamp 1698431365
transform 1 0 32704 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_511
timestamp 1698431365
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_512
timestamp 1698431365
transform 1 0 13104 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_513
timestamp 1698431365
transform 1 0 20944 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_514
timestamp 1698431365
transform 1 0 28784 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_515
timestamp 1698431365
transform 1 0 36624 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_516
timestamp 1698431365
transform 1 0 9184 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_517
timestamp 1698431365
transform 1 0 17024 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_518
timestamp 1698431365
transform 1 0 24864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_519
timestamp 1698431365
transform 1 0 32704 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_520
timestamp 1698431365
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_521
timestamp 1698431365
transform 1 0 13104 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_522
timestamp 1698431365
transform 1 0 20944 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_523
timestamp 1698431365
transform 1 0 28784 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_524
timestamp 1698431365
transform 1 0 36624 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_525
timestamp 1698431365
transform 1 0 9184 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_526
timestamp 1698431365
transform 1 0 17024 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_527
timestamp 1698431365
transform 1 0 24864 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_528
timestamp 1698431365
transform 1 0 32704 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_529
timestamp 1698431365
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_530
timestamp 1698431365
transform 1 0 13104 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_531
timestamp 1698431365
transform 1 0 20944 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_532
timestamp 1698431365
transform 1 0 28784 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_533
timestamp 1698431365
transform 1 0 36624 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_534
timestamp 1698431365
transform 1 0 9184 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_535
timestamp 1698431365
transform 1 0 17024 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_536
timestamp 1698431365
transform 1 0 24864 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_537
timestamp 1698431365
transform 1 0 32704 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_538
timestamp 1698431365
transform 1 0 5264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_539
timestamp 1698431365
transform 1 0 13104 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_540
timestamp 1698431365
transform 1 0 20944 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_541
timestamp 1698431365
transform 1 0 28784 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_542
timestamp 1698431365
transform 1 0 36624 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_543
timestamp 1698431365
transform 1 0 9184 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_544
timestamp 1698431365
transform 1 0 17024 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_545
timestamp 1698431365
transform 1 0 24864 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_546
timestamp 1698431365
transform 1 0 32704 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_547
timestamp 1698431365
transform 1 0 5264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_548
timestamp 1698431365
transform 1 0 13104 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_549
timestamp 1698431365
transform 1 0 20944 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_550
timestamp 1698431365
transform 1 0 28784 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_551
timestamp 1698431365
transform 1 0 36624 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_552
timestamp 1698431365
transform 1 0 9184 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_553
timestamp 1698431365
transform 1 0 17024 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_554
timestamp 1698431365
transform 1 0 24864 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_555
timestamp 1698431365
transform 1 0 32704 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_556
timestamp 1698431365
transform 1 0 5264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_557
timestamp 1698431365
transform 1 0 13104 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_558
timestamp 1698431365
transform 1 0 20944 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_559
timestamp 1698431365
transform 1 0 28784 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_560
timestamp 1698431365
transform 1 0 36624 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_561
timestamp 1698431365
transform 1 0 9184 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_562
timestamp 1698431365
transform 1 0 17024 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_563
timestamp 1698431365
transform 1 0 24864 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_564
timestamp 1698431365
transform 1 0 32704 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_565
timestamp 1698431365
transform 1 0 5264 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_566
timestamp 1698431365
transform 1 0 13104 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_567
timestamp 1698431365
transform 1 0 20944 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_568
timestamp 1698431365
transform 1 0 28784 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_569
timestamp 1698431365
transform 1 0 36624 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_570
timestamp 1698431365
transform 1 0 9184 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_571
timestamp 1698431365
transform 1 0 17024 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_572
timestamp 1698431365
transform 1 0 24864 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_573
timestamp 1698431365
transform 1 0 32704 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_574
timestamp 1698431365
transform 1 0 5264 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_575
timestamp 1698431365
transform 1 0 13104 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_576
timestamp 1698431365
transform 1 0 20944 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_577
timestamp 1698431365
transform 1 0 28784 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_578
timestamp 1698431365
transform 1 0 36624 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_579
timestamp 1698431365
transform 1 0 9184 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_580
timestamp 1698431365
transform 1 0 17024 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_581
timestamp 1698431365
transform 1 0 24864 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_582
timestamp 1698431365
transform 1 0 32704 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_583
timestamp 1698431365
transform 1 0 5264 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_584
timestamp 1698431365
transform 1 0 13104 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_585
timestamp 1698431365
transform 1 0 20944 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_586
timestamp 1698431365
transform 1 0 28784 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_587
timestamp 1698431365
transform 1 0 36624 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_588
timestamp 1698431365
transform 1 0 9184 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_589
timestamp 1698431365
transform 1 0 17024 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_590
timestamp 1698431365
transform 1 0 24864 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_591
timestamp 1698431365
transform 1 0 32704 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_592
timestamp 1698431365
transform 1 0 5264 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_593
timestamp 1698431365
transform 1 0 13104 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_594
timestamp 1698431365
transform 1 0 20944 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_595
timestamp 1698431365
transform 1 0 28784 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_596
timestamp 1698431365
transform 1 0 36624 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_597
timestamp 1698431365
transform 1 0 9184 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_598
timestamp 1698431365
transform 1 0 17024 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_599
timestamp 1698431365
transform 1 0 24864 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_600
timestamp 1698431365
transform 1 0 32704 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_601
timestamp 1698431365
transform 1 0 5264 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_602
timestamp 1698431365
transform 1 0 13104 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_603
timestamp 1698431365
transform 1 0 20944 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_604
timestamp 1698431365
transform 1 0 28784 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_605
timestamp 1698431365
transform 1 0 36624 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_606
timestamp 1698431365
transform 1 0 9184 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_607
timestamp 1698431365
transform 1 0 17024 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_608
timestamp 1698431365
transform 1 0 24864 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_609
timestamp 1698431365
transform 1 0 32704 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_610
timestamp 1698431365
transform 1 0 5264 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_611
timestamp 1698431365
transform 1 0 13104 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_612
timestamp 1698431365
transform 1 0 20944 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_613
timestamp 1698431365
transform 1 0 28784 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_614
timestamp 1698431365
transform 1 0 36624 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_615
timestamp 1698431365
transform 1 0 9184 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_616
timestamp 1698431365
transform 1 0 17024 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_617
timestamp 1698431365
transform 1 0 24864 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_618
timestamp 1698431365
transform 1 0 32704 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_619
timestamp 1698431365
transform 1 0 5264 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_620
timestamp 1698431365
transform 1 0 13104 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_621
timestamp 1698431365
transform 1 0 20944 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_622
timestamp 1698431365
transform 1 0 28784 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_623
timestamp 1698431365
transform 1 0 36624 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_624
timestamp 1698431365
transform 1 0 9184 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_625
timestamp 1698431365
transform 1 0 17024 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_626
timestamp 1698431365
transform 1 0 24864 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_627
timestamp 1698431365
transform 1 0 32704 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_628
timestamp 1698431365
transform 1 0 5264 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_629
timestamp 1698431365
transform 1 0 13104 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_630
timestamp 1698431365
transform 1 0 20944 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_631
timestamp 1698431365
transform 1 0 28784 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_632
timestamp 1698431365
transform 1 0 36624 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_633
timestamp 1698431365
transform 1 0 9184 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_634
timestamp 1698431365
transform 1 0 17024 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_635
timestamp 1698431365
transform 1 0 24864 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_636
timestamp 1698431365
transform 1 0 32704 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_637
timestamp 1698431365
transform 1 0 5264 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_638
timestamp 1698431365
transform 1 0 13104 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_639
timestamp 1698431365
transform 1 0 20944 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_640
timestamp 1698431365
transform 1 0 28784 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_641
timestamp 1698431365
transform 1 0 36624 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_642
timestamp 1698431365
transform 1 0 9184 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_643
timestamp 1698431365
transform 1 0 17024 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_644
timestamp 1698431365
transform 1 0 24864 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_645
timestamp 1698431365
transform 1 0 32704 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_646
timestamp 1698431365
transform 1 0 5264 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_647
timestamp 1698431365
transform 1 0 13104 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_648
timestamp 1698431365
transform 1 0 20944 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_649
timestamp 1698431365
transform 1 0 28784 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_650
timestamp 1698431365
transform 1 0 36624 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_651
timestamp 1698431365
transform 1 0 9184 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_652
timestamp 1698431365
transform 1 0 17024 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_653
timestamp 1698431365
transform 1 0 24864 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_654
timestamp 1698431365
transform 1 0 32704 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_655
timestamp 1698431365
transform 1 0 5264 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_656
timestamp 1698431365
transform 1 0 13104 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_657
timestamp 1698431365
transform 1 0 20944 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_658
timestamp 1698431365
transform 1 0 28784 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_659
timestamp 1698431365
transform 1 0 36624 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_660
timestamp 1698431365
transform 1 0 9184 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_661
timestamp 1698431365
transform 1 0 17024 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_662
timestamp 1698431365
transform 1 0 24864 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_663
timestamp 1698431365
transform 1 0 32704 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_664
timestamp 1698431365
transform 1 0 5264 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_665
timestamp 1698431365
transform 1 0 13104 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_666
timestamp 1698431365
transform 1 0 20944 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_667
timestamp 1698431365
transform 1 0 28784 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_668
timestamp 1698431365
transform 1 0 36624 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_669
timestamp 1698431365
transform 1 0 9184 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_670
timestamp 1698431365
transform 1 0 17024 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_671
timestamp 1698431365
transform 1 0 24864 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_672
timestamp 1698431365
transform 1 0 32704 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_94_673
timestamp 1698431365
transform 1 0 5264 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_94_674
timestamp 1698431365
transform 1 0 13104 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_94_675
timestamp 1698431365
transform 1 0 20944 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_94_676
timestamp 1698431365
transform 1 0 28784 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_94_677
timestamp 1698431365
transform 1 0 36624 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_95_678
timestamp 1698431365
transform 1 0 9184 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_95_679
timestamp 1698431365
transform 1 0 17024 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_95_680
timestamp 1698431365
transform 1 0 24864 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_95_681
timestamp 1698431365
transform 1 0 32704 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_96_682
timestamp 1698431365
transform 1 0 5264 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_96_683
timestamp 1698431365
transform 1 0 13104 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_96_684
timestamp 1698431365
transform 1 0 20944 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_96_685
timestamp 1698431365
transform 1 0 28784 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_96_686
timestamp 1698431365
transform 1 0 36624 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_97_687
timestamp 1698431365
transform 1 0 9184 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_97_688
timestamp 1698431365
transform 1 0 17024 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_97_689
timestamp 1698431365
transform 1 0 24864 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_97_690
timestamp 1698431365
transform 1 0 32704 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_98_691
timestamp 1698431365
transform 1 0 5264 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_98_692
timestamp 1698431365
transform 1 0 13104 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_98_693
timestamp 1698431365
transform 1 0 20944 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_98_694
timestamp 1698431365
transform 1 0 28784 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_98_695
timestamp 1698431365
transform 1 0 36624 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_99_696
timestamp 1698431365
transform 1 0 9184 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_99_697
timestamp 1698431365
transform 1 0 17024 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_99_698
timestamp 1698431365
transform 1 0 24864 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_99_699
timestamp 1698431365
transform 1 0 32704 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_100_700
timestamp 1698431365
transform 1 0 5264 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_100_701
timestamp 1698431365
transform 1 0 13104 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_100_702
timestamp 1698431365
transform 1 0 20944 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_100_703
timestamp 1698431365
transform 1 0 28784 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_100_704
timestamp 1698431365
transform 1 0 36624 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_101_705
timestamp 1698431365
transform 1 0 9184 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_101_706
timestamp 1698431365
transform 1 0 17024 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_101_707
timestamp 1698431365
transform 1 0 24864 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_101_708
timestamp 1698431365
transform 1 0 32704 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_102_709
timestamp 1698431365
transform 1 0 5264 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_102_710
timestamp 1698431365
transform 1 0 13104 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_102_711
timestamp 1698431365
transform 1 0 20944 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_102_712
timestamp 1698431365
transform 1 0 28784 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_102_713
timestamp 1698431365
transform 1 0 36624 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_103_714
timestamp 1698431365
transform 1 0 9184 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_103_715
timestamp 1698431365
transform 1 0 17024 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_103_716
timestamp 1698431365
transform 1 0 24864 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_103_717
timestamp 1698431365
transform 1 0 32704 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_104_718
timestamp 1698431365
transform 1 0 5264 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_104_719
timestamp 1698431365
transform 1 0 13104 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_104_720
timestamp 1698431365
transform 1 0 20944 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_104_721
timestamp 1698431365
transform 1 0 28784 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_104_722
timestamp 1698431365
transform 1 0 36624 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_105_723
timestamp 1698431365
transform 1 0 9184 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_105_724
timestamp 1698431365
transform 1 0 17024 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_105_725
timestamp 1698431365
transform 1 0 24864 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_105_726
timestamp 1698431365
transform 1 0 32704 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_106_727
timestamp 1698431365
transform 1 0 5264 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_106_728
timestamp 1698431365
transform 1 0 13104 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_106_729
timestamp 1698431365
transform 1 0 20944 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_106_730
timestamp 1698431365
transform 1 0 28784 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_106_731
timestamp 1698431365
transform 1 0 36624 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_107_732
timestamp 1698431365
transform 1 0 9184 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_107_733
timestamp 1698431365
transform 1 0 17024 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_107_734
timestamp 1698431365
transform 1 0 24864 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_107_735
timestamp 1698431365
transform 1 0 32704 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_108_736
timestamp 1698431365
transform 1 0 5264 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_108_737
timestamp 1698431365
transform 1 0 13104 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_108_738
timestamp 1698431365
transform 1 0 20944 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_108_739
timestamp 1698431365
transform 1 0 28784 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_108_740
timestamp 1698431365
transform 1 0 36624 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_109_741
timestamp 1698431365
transform 1 0 9184 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_109_742
timestamp 1698431365
transform 1 0 17024 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_109_743
timestamp 1698431365
transform 1 0 24864 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_109_744
timestamp 1698431365
transform 1 0 32704 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_110_745
timestamp 1698431365
transform 1 0 5264 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_110_746
timestamp 1698431365
transform 1 0 13104 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_110_747
timestamp 1698431365
transform 1 0 20944 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_110_748
timestamp 1698431365
transform 1 0 28784 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_110_749
timestamp 1698431365
transform 1 0 36624 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_111_750
timestamp 1698431365
transform 1 0 9184 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_111_751
timestamp 1698431365
transform 1 0 17024 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_111_752
timestamp 1698431365
transform 1 0 24864 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_111_753
timestamp 1698431365
transform 1 0 32704 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_112_754
timestamp 1698431365
transform 1 0 5264 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_112_755
timestamp 1698431365
transform 1 0 13104 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_112_756
timestamp 1698431365
transform 1 0 20944 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_112_757
timestamp 1698431365
transform 1 0 28784 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_112_758
timestamp 1698431365
transform 1 0 36624 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_113_759
timestamp 1698431365
transform 1 0 9184 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_113_760
timestamp 1698431365
transform 1 0 17024 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_113_761
timestamp 1698431365
transform 1 0 24864 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_113_762
timestamp 1698431365
transform 1 0 32704 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_114_763
timestamp 1698431365
transform 1 0 5264 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_114_764
timestamp 1698431365
transform 1 0 13104 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_114_765
timestamp 1698431365
transform 1 0 20944 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_114_766
timestamp 1698431365
transform 1 0 28784 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_114_767
timestamp 1698431365
transform 1 0 36624 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_115_768
timestamp 1698431365
transform 1 0 9184 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_115_769
timestamp 1698431365
transform 1 0 17024 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_115_770
timestamp 1698431365
transform 1 0 24864 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_115_771
timestamp 1698431365
transform 1 0 32704 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_116_772
timestamp 1698431365
transform 1 0 5264 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_116_773
timestamp 1698431365
transform 1 0 13104 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_116_774
timestamp 1698431365
transform 1 0 20944 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_116_775
timestamp 1698431365
transform 1 0 28784 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_116_776
timestamp 1698431365
transform 1 0 36624 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_117_777
timestamp 1698431365
transform 1 0 9184 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_117_778
timestamp 1698431365
transform 1 0 17024 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_117_779
timestamp 1698431365
transform 1 0 24864 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_117_780
timestamp 1698431365
transform 1 0 32704 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_118_781
timestamp 1698431365
transform 1 0 5264 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_118_782
timestamp 1698431365
transform 1 0 13104 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_118_783
timestamp 1698431365
transform 1 0 20944 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_118_784
timestamp 1698431365
transform 1 0 28784 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_118_785
timestamp 1698431365
transform 1 0 36624 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_119_786
timestamp 1698431365
transform 1 0 9184 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_119_787
timestamp 1698431365
transform 1 0 17024 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_119_788
timestamp 1698431365
transform 1 0 24864 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_119_789
timestamp 1698431365
transform 1 0 32704 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_120_790
timestamp 1698431365
transform 1 0 5264 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_120_791
timestamp 1698431365
transform 1 0 13104 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_120_792
timestamp 1698431365
transform 1 0 20944 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_120_793
timestamp 1698431365
transform 1 0 28784 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_120_794
timestamp 1698431365
transform 1 0 36624 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_121_795
timestamp 1698431365
transform 1 0 9184 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_121_796
timestamp 1698431365
transform 1 0 17024 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_121_797
timestamp 1698431365
transform 1 0 24864 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_121_798
timestamp 1698431365
transform 1 0 32704 0 -1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_122_799
timestamp 1698431365
transform 1 0 5152 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_122_800
timestamp 1698431365
transform 1 0 8960 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_122_801
timestamp 1698431365
transform 1 0 12768 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_122_802
timestamp 1698431365
transform 1 0 16576 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_122_803
timestamp 1698431365
transform 1 0 20384 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_122_804
timestamp 1698431365
transform 1 0 24192 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_122_805
timestamp 1698431365
transform 1 0 28000 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_122_806
timestamp 1698431365
transform 1 0 31808 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_122_807
timestamp 1698431365
transform 1 0 35616 0 1 97216
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  temp1.dac._4_
timestamp 1698431365
transform -1 0 14896 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  temp1.dac._5_
timestamp 1698431365
transform 1 0 13328 0 1 90944
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  temp1.dac.parallel_cells\[0\].vdac_batch._3_
timestamp 1698431365
transform 1 0 25424 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  temp1.dac.parallel_cells\[0\].vdac_batch._4_
timestamp 1698431365
transform 1 0 23408 0 -1 94080
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  temp1.dac.parallel_cells\[0\].vdac_batch._5_
timestamp 1698431365
transform -1 0 24864 0 1 92512
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  temp1.dac.parallel_cells\[0\].vdac_batch._6_
timestamp 1698431365
transform 1 0 24192 0 1 94080
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  temp1.dac.parallel_cells\[0\].vdac_batch._7_
timestamp 1698431365
transform -1 0 25984 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  temp1.dac.parallel_cells\[0\].vdac_batch._8_
timestamp 1698431365
transform 1 0 24864 0 1 94080
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].pupd open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 -1 94080
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].vref
timestamp 1698431365
transform 1 0 25088 0 -1 95648
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  temp1.dac.parallel_cells\[1\].vdac_batch._3_
timestamp 1698431365
transform -1 0 23520 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  temp1.dac.parallel_cells\[1\].vdac_batch._4_
timestamp 1698431365
transform -1 0 22064 0 -1 92512
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  temp1.dac.parallel_cells\[1\].vdac_batch._5_
timestamp 1698431365
transform 1 0 19936 0 -1 94080
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  temp1.dac.parallel_cells\[1\].vdac_batch._6_
timestamp 1698431365
transform -1 0 21840 0 1 94080
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  temp1.dac.parallel_cells\[1\].vdac_batch._7_
timestamp 1698431365
transform -1 0 22960 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  temp1.dac.parallel_cells\[1\].vdac_batch._8_
timestamp 1698431365
transform 1 0 21840 0 1 94080
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[0\].pupd
timestamp 1698431365
transform 1 0 20832 0 -1 94080
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[0\].vref
timestamp 1698431365
transform 1 0 21168 0 1 95648
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].pupd
timestamp 1698431365
transform 1 0 21168 0 1 92512
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].vref
timestamp 1698431365
transform -1 0 22400 0 -1 95648
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  temp1.dac.parallel_cells\[2\].vdac_batch._3_
timestamp 1698431365
transform -1 0 19600 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  temp1.dac.parallel_cells\[2\].vdac_batch._4_
timestamp 1698431365
transform -1 0 18368 0 1 92512
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  temp1.dac.parallel_cells\[2\].vdac_batch._5_
timestamp 1698431365
transform -1 0 17024 0 -1 94080
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  temp1.dac.parallel_cells\[2\].vdac_batch._6_
timestamp 1698431365
transform 1 0 16352 0 -1 95648
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  temp1.dac.parallel_cells\[2\].vdac_batch._7_
timestamp 1698431365
transform -1 0 17024 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  temp1.dac.parallel_cells\[2\].vdac_batch._8_
timestamp 1698431365
transform -1 0 16576 0 1 94080
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd
timestamp 1698431365
transform 1 0 17248 0 -1 95648
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].vref
timestamp 1698431365
transform 1 0 13328 0 1 95648
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].pupd
timestamp 1698431365
transform 1 0 17248 0 -1 94080
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref
timestamp 1698431365
transform -1 0 14896 0 -1 95648
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[2\].pupd
timestamp 1698431365
transform 1 0 17248 0 1 95648
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[2\].vref
timestamp 1698431365
transform -1 0 15568 0 1 97216
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].pupd
timestamp 1698431365
transform 1 0 18368 0 1 94080
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].vref
timestamp 1698431365
transform -1 0 14896 0 -1 97216
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  temp1.dac.parallel_cells\[3\].vdac_batch._3_
timestamp 1698431365
transform -1 0 14112 0 -1 87808
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  temp1.dac.parallel_cells\[3\].vdac_batch._4_
timestamp 1698431365
transform -1 0 13440 0 -1 87808
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  temp1.dac.parallel_cells\[3\].vdac_batch._5_
timestamp 1698431365
transform -1 0 12992 0 1 87808
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  temp1.dac.parallel_cells\[3\].vdac_batch._6_
timestamp 1698431365
transform -1 0 10864 0 1 86240
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  temp1.dac.parallel_cells\[3\].vdac_batch._7_
timestamp 1698431365
transform 1 0 11424 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  temp1.dac.parallel_cells\[3\].vdac_batch._8_
timestamp 1698431365
transform 1 0 10864 0 1 86240
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[0\].pupd
timestamp 1698431365
transform 1 0 6608 0 -1 87808
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[0\].vref
timestamp 1698431365
transform -1 0 4480 0 -1 86240
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd
timestamp 1698431365
transform 1 0 6608 0 -1 89376
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref
timestamp 1698431365
transform -1 0 4480 0 1 83104
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[2\].pupd
timestamp 1698431365
transform 1 0 6944 0 1 87808
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[2\].vref
timestamp 1698431365
transform 1 0 4480 0 -1 86240
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[3\].pupd
timestamp 1698431365
transform -1 0 9520 0 1 86240
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[3\].vref
timestamp 1698431365
transform -1 0 4480 0 -1 87808
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd
timestamp 1698431365
transform -1 0 8288 0 1 89376
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref
timestamp 1698431365
transform -1 0 4480 0 1 87808
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[5\].pupd
timestamp 1698431365
transform 1 0 9408 0 -1 87808
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[5\].vref
timestamp 1698431365
transform -1 0 4480 0 1 84672
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[6\].pupd
timestamp 1698431365
transform 1 0 8288 0 1 89376
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[6\].vref
timestamp 1698431365
transform -1 0 4480 0 -1 84672
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd
timestamp 1698431365
transform 1 0 9520 0 1 87808
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref
timestamp 1698431365
transform -1 0 4480 0 1 86240
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  temp1.dac.parallel_cells\[4\].vdac_batch._3_
timestamp 1698431365
transform 1 0 27216 0 -1 92512
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_2  temp1.dac.parallel_cells\[4\].vdac_batch._4_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 26992 0 -1 92512
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  temp1.dac.parallel_cells\[4\].vdac_batch._5_
timestamp 1698431365
transform 1 0 25312 0 -1 90944
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  temp1.dac.parallel_cells\[4\].vdac_batch._6_
timestamp 1698431365
transform 1 0 26544 0 1 92512
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  temp1.dac.parallel_cells\[4\].vdac_batch._7_
timestamp 1698431365
transform 1 0 10080 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  temp1.dac.parallel_cells\[4\].vdac_batch._8_
timestamp 1698431365
transform 1 0 10528 0 -1 92512
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[0\].pupd
timestamp 1698431365
transform 1 0 29008 0 1 92512
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[0\].vref
timestamp 1698431365
transform 1 0 3696 0 -1 95648
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[1\].pupd
timestamp 1698431365
transform -1 0 34832 0 1 90944
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[1\].vref
timestamp 1698431365
transform 1 0 6608 0 -1 95648
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].pupd
timestamp 1698431365
transform -1 0 35504 0 -1 97216
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref
timestamp 1698431365
transform -1 0 9184 0 -1 97216
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[3\].pupd
timestamp 1698431365
transform 1 0 29008 0 1 94080
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[3\].vref
timestamp 1698431365
transform -1 0 4592 0 1 89376
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[4\].pupd
timestamp 1698431365
transform 1 0 29008 0 1 95648
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[4\].vref
timestamp 1698431365
transform 1 0 9184 0 1 95648
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[5\].pupd
timestamp 1698431365
transform 1 0 32704 0 1 94080
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[5\].vref
timestamp 1698431365
transform 1 0 2688 0 1 92512
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[6\].pupd
timestamp 1698431365
transform 1 0 32928 0 -1 92512
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_4  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[6\].vref open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2688 0 -1 92512
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].pupd
timestamp 1698431365
transform 1 0 35504 0 -1 95648
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].vref
timestamp 1698431365
transform 1 0 6608 0 -1 94080
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd
timestamp 1698431365
transform 1 0 32928 0 -1 94080
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].vref
timestamp 1698431365
transform -1 0 4368 0 -1 94080
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[9\].pupd
timestamp 1698431365
transform 1 0 31584 0 1 92512
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[9\].vref
timestamp 1698431365
transform 1 0 2688 0 1 94080
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[10\].pupd
timestamp 1698431365
transform 1 0 32704 0 1 95648
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[10\].vref
timestamp 1698431365
transform 1 0 2912 0 -1 90944
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[11\].pupd
timestamp 1698431365
transform -1 0 32480 0 -1 97216
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[11\].vref
timestamp 1698431365
transform 1 0 2688 0 1 95648
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd
timestamp 1698431365
transform -1 0 28784 0 1 94080
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref
timestamp 1698431365
transform 1 0 6272 0 -1 92512
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd
timestamp 1698431365
transform 1 0 32928 0 -1 95648
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].vref
timestamp 1698431365
transform 1 0 2688 0 1 90944
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[14\].pupd
timestamp 1698431365
transform 1 0 28560 0 -1 94080
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_4  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[14\].vref
timestamp 1698431365
transform 1 0 6496 0 1 95648
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd
timestamp 1698431365
transform 1 0 28000 0 -1 95648
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].vref
timestamp 1698431365
transform 1 0 6832 0 1 92512
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  temp1.dac.vdac_single._3_
timestamp 1698431365
transform -1 0 13552 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  temp1.dac.vdac_single._3__63 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 14448 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  temp1.dac.vdac_single._4__65
timestamp 1698431365
transform -1 0 14896 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  temp1.dac.vdac_single._4_
timestamp 1698431365
transform 1 0 11648 0 -1 94080
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  temp1.dac.vdac_single._4__64
timestamp 1698431365
transform 1 0 10080 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  temp1.dac.vdac_single._5_
timestamp 1698431365
transform 1 0 11872 0 1 90944
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  temp1.dac.vdac_single._6_
timestamp 1698431365
transform -1 0 14000 0 1 92512
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  temp1.dac.vdac_single._7_
timestamp 1698431365
transform 1 0 11424 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  temp1.dac.vdac_single._8_
timestamp 1698431365
transform -1 0 12880 0 -1 90944
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.vdac_single.einvp_batch\[0\].pupd
timestamp 1698431365
transform -1 0 13104 0 1 92512
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  temp1.dac.vdac_single.einvp_batch\[0\].vref open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12544 0 -1 92512
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  temp1.dcdc
timestamp 1698431365
transform 1 0 21840 0 -1 89376
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  temp1.inv1_1
timestamp 1698431365
transform 1 0 20496 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  temp1.inv2_2
timestamp 1698431365
transform -1 0 23632 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  temp1.inv2_3
timestamp 1698431365
transform -1 0 25536 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  temp_sensor_54
timestamp 1698431365
transform -1 0 19152 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  temp_sensor_55
timestamp 1698431365
transform -1 0 17248 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  temp_sensor_56
timestamp 1698431365
transform -1 0 16016 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  temp_sensor_57
timestamp 1698431365
transform -1 0 11760 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  temp_sensor_58
timestamp 1698431365
transform -1 0 9632 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  temp_sensor_59
timestamp 1698431365
transform -1 0 6832 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  temp_sensor_60
timestamp 1698431365
transform -1 0 4368 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  temp_sensor_61
timestamp 1698431365
transform -1 0 2016 0 1 97216
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  temp_sensor_62
timestamp 1698431365
transform -1 0 2016 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  wire4
timestamp 1698431365
transform 1 0 8288 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  wire5
timestamp 1698431365
transform -1 0 11088 0 1 50176
box -86 -86 758 870
<< labels >>
flabel metal4 s 4448 1508 4768 98060 0 FreeSans 1280 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 35168 1508 35488 98060 0 FreeSans 1280 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 19808 1508 20128 98060 0 FreeSans 1280 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal2 s 4704 0 4816 400 0 FreeSans 448 90 0 0 clk
port 2 nsew signal input
flabel metal2 s 36064 0 36176 400 0 FreeSans 448 90 0 0 i_wb_addr[0]
port 3 nsew signal input
flabel metal2 s 27104 0 27216 400 0 FreeSans 448 90 0 0 i_wb_addr[10]
port 4 nsew signal input
flabel metal2 s 26208 0 26320 400 0 FreeSans 448 90 0 0 i_wb_addr[11]
port 5 nsew signal input
flabel metal2 s 25312 0 25424 400 0 FreeSans 448 90 0 0 i_wb_addr[12]
port 6 nsew signal input
flabel metal2 s 24416 0 24528 400 0 FreeSans 448 90 0 0 i_wb_addr[13]
port 7 nsew signal input
flabel metal2 s 23520 0 23632 400 0 FreeSans 448 90 0 0 i_wb_addr[14]
port 8 nsew signal input
flabel metal2 s 22624 0 22736 400 0 FreeSans 448 90 0 0 i_wb_addr[15]
port 9 nsew signal input
flabel metal2 s 21728 0 21840 400 0 FreeSans 448 90 0 0 i_wb_addr[16]
port 10 nsew signal input
flabel metal2 s 20832 0 20944 400 0 FreeSans 448 90 0 0 i_wb_addr[17]
port 11 nsew signal input
flabel metal2 s 19936 0 20048 400 0 FreeSans 448 90 0 0 i_wb_addr[18]
port 12 nsew signal input
flabel metal2 s 19040 0 19152 400 0 FreeSans 448 90 0 0 i_wb_addr[19]
port 13 nsew signal input
flabel metal2 s 35168 0 35280 400 0 FreeSans 448 90 0 0 i_wb_addr[1]
port 14 nsew signal input
flabel metal2 s 18144 0 18256 400 0 FreeSans 448 90 0 0 i_wb_addr[20]
port 15 nsew signal input
flabel metal2 s 17248 0 17360 400 0 FreeSans 448 90 0 0 i_wb_addr[21]
port 16 nsew signal input
flabel metal2 s 16352 0 16464 400 0 FreeSans 448 90 0 0 i_wb_addr[22]
port 17 nsew signal input
flabel metal2 s 15456 0 15568 400 0 FreeSans 448 90 0 0 i_wb_addr[23]
port 18 nsew signal input
flabel metal2 s 14560 0 14672 400 0 FreeSans 448 90 0 0 i_wb_addr[24]
port 19 nsew signal input
flabel metal2 s 13664 0 13776 400 0 FreeSans 448 90 0 0 i_wb_addr[25]
port 20 nsew signal input
flabel metal2 s 12768 0 12880 400 0 FreeSans 448 90 0 0 i_wb_addr[26]
port 21 nsew signal input
flabel metal2 s 11872 0 11984 400 0 FreeSans 448 90 0 0 i_wb_addr[27]
port 22 nsew signal input
flabel metal2 s 10976 0 11088 400 0 FreeSans 448 90 0 0 i_wb_addr[28]
port 23 nsew signal input
flabel metal2 s 10080 0 10192 400 0 FreeSans 448 90 0 0 i_wb_addr[29]
port 24 nsew signal input
flabel metal2 s 34272 0 34384 400 0 FreeSans 448 90 0 0 i_wb_addr[2]
port 25 nsew signal input
flabel metal2 s 9184 0 9296 400 0 FreeSans 448 90 0 0 i_wb_addr[30]
port 26 nsew signal input
flabel metal2 s 8288 0 8400 400 0 FreeSans 448 90 0 0 i_wb_addr[31]
port 27 nsew signal input
flabel metal2 s 33376 0 33488 400 0 FreeSans 448 90 0 0 i_wb_addr[3]
port 28 nsew signal input
flabel metal2 s 32480 0 32592 400 0 FreeSans 448 90 0 0 i_wb_addr[4]
port 29 nsew signal input
flabel metal2 s 31584 0 31696 400 0 FreeSans 448 90 0 0 i_wb_addr[5]
port 30 nsew signal input
flabel metal2 s 30688 0 30800 400 0 FreeSans 448 90 0 0 i_wb_addr[6]
port 31 nsew signal input
flabel metal2 s 29792 0 29904 400 0 FreeSans 448 90 0 0 i_wb_addr[7]
port 32 nsew signal input
flabel metal2 s 28896 0 29008 400 0 FreeSans 448 90 0 0 i_wb_addr[8]
port 33 nsew signal input
flabel metal2 s 28000 0 28112 400 0 FreeSans 448 90 0 0 i_wb_addr[9]
port 34 nsew signal input
flabel metal2 s 7392 0 7504 400 0 FreeSans 448 90 0 0 i_wb_cyc
port 35 nsew signal input
flabel metal2 s 6496 0 6608 400 0 FreeSans 448 90 0 0 i_wb_stb
port 36 nsew signal input
flabel metal2 s 5600 0 5712 400 0 FreeSans 448 90 0 0 i_wb_we
port 37 nsew signal input
flabel metal3 s 39600 8512 40000 8624 0 FreeSans 448 0 0 0 io_in[0]
port 38 nsew signal input
flabel metal3 s 39600 25088 40000 25200 0 FreeSans 448 0 0 0 io_in[1]
port 39 nsew signal input
flabel metal3 s 39600 41664 40000 41776 0 FreeSans 448 0 0 0 io_in[2]
port 40 nsew signal input
flabel metal3 s 39600 58240 40000 58352 0 FreeSans 448 0 0 0 io_in[3]
port 41 nsew signal input
flabel metal3 s 39600 74816 40000 74928 0 FreeSans 448 0 0 0 io_in[4]
port 42 nsew signal input
flabel metal3 s 39600 91392 40000 91504 0 FreeSans 448 0 0 0 io_in[5]
port 43 nsew signal input
flabel metal2 s 18592 99600 18704 100000 0 FreeSans 448 90 0 0 io_oeb[0]
port 44 nsew signal tristate
flabel metal2 s 16128 99600 16240 100000 0 FreeSans 448 90 0 0 io_oeb[1]
port 45 nsew signal tristate
flabel metal2 s 13664 99600 13776 100000 0 FreeSans 448 90 0 0 io_oeb[2]
port 46 nsew signal tristate
flabel metal2 s 11200 99600 11312 100000 0 FreeSans 448 90 0 0 io_oeb[3]
port 47 nsew signal tristate
flabel metal2 s 8736 99600 8848 100000 0 FreeSans 448 90 0 0 io_oeb[4]
port 48 nsew signal tristate
flabel metal2 s 6272 99600 6384 100000 0 FreeSans 448 90 0 0 io_oeb[5]
port 49 nsew signal tristate
flabel metal2 s 3808 99600 3920 100000 0 FreeSans 448 90 0 0 io_oeb[6]
port 50 nsew signal tristate
flabel metal2 s 1344 99600 1456 100000 0 FreeSans 448 90 0 0 io_oeb[7]
port 51 nsew signal tristate
flabel metal2 s 38304 99600 38416 100000 0 FreeSans 448 90 0 0 io_out[0]
port 52 nsew signal tristate
flabel metal2 s 35840 99600 35952 100000 0 FreeSans 448 90 0 0 io_out[1]
port 53 nsew signal tristate
flabel metal2 s 33376 99600 33488 100000 0 FreeSans 448 90 0 0 io_out[2]
port 54 nsew signal tristate
flabel metal2 s 30912 99600 31024 100000 0 FreeSans 448 90 0 0 io_out[3]
port 55 nsew signal tristate
flabel metal2 s 28448 99600 28560 100000 0 FreeSans 448 90 0 0 io_out[4]
port 56 nsew signal tristate
flabel metal2 s 25984 99600 26096 100000 0 FreeSans 448 90 0 0 io_out[5]
port 57 nsew signal tristate
flabel metal2 s 23520 99600 23632 100000 0 FreeSans 448 90 0 0 io_out[6]
port 58 nsew signal tristate
flabel metal2 s 21056 99600 21168 100000 0 FreeSans 448 90 0 0 io_out[7]
port 59 nsew signal tristate
flabel metal3 s 0 5600 400 5712 0 FreeSans 448 0 0 0 o_wb_ack
port 60 nsew signal tristate
flabel metal3 s 0 15456 400 15568 0 FreeSans 448 0 0 0 o_wb_data[0]
port 61 nsew signal tristate
flabel metal3 s 0 25312 400 25424 0 FreeSans 448 0 0 0 o_wb_data[1]
port 62 nsew signal tristate
flabel metal3 s 0 35168 400 35280 0 FreeSans 448 0 0 0 o_wb_data[2]
port 63 nsew signal tristate
flabel metal3 s 0 45024 400 45136 0 FreeSans 448 0 0 0 o_wb_data[3]
port 64 nsew signal tristate
flabel metal3 s 0 54880 400 54992 0 FreeSans 448 0 0 0 o_wb_data[4]
port 65 nsew signal tristate
flabel metal3 s 0 64736 400 64848 0 FreeSans 448 0 0 0 o_wb_data[5]
port 66 nsew signal tristate
flabel metal3 s 0 74592 400 74704 0 FreeSans 448 0 0 0 o_wb_data[6]
port 67 nsew signal tristate
flabel metal3 s 0 84448 400 84560 0 FreeSans 448 0 0 0 o_wb_data[7]
port 68 nsew signal tristate
flabel metal3 s 0 94304 400 94416 0 FreeSans 448 0 0 0 o_wb_stall
port 69 nsew signal tristate
flabel metal2 s 3808 0 3920 400 0 FreeSans 448 90 0 0 reset
port 70 nsew signal input
rlabel metal1 19992 98000 19992 98000 0 VDD
rlabel via1 19992 97216 19992 97216 0 VSS
rlabel metal3 10304 81816 10304 81816 0 _0000_
rlabel metal2 5880 81312 5880 81312 0 _0001_
rlabel metal2 5992 77896 5992 77896 0 _0002_
rlabel metal3 7336 74760 7336 74760 0 _0003_
rlabel metal2 4312 74928 4312 74928 0 _0004_
rlabel metal2 9464 77560 9464 77560 0 _0005_
rlabel metal2 9800 75880 9800 75880 0 _0006_
rlabel metal2 8288 82824 8288 82824 0 _0007_
rlabel metal2 7784 4648 7784 4648 0 _0008_
rlabel metal2 37464 26600 37464 26600 0 _0009_
rlabel metal2 26488 32480 26488 32480 0 _0010_
rlabel metal2 27608 32704 27608 32704 0 _0011_
rlabel metal2 28056 38668 28056 38668 0 _0012_
rlabel metal2 29736 52864 29736 52864 0 _0013_
rlabel metal2 28112 55272 28112 55272 0 _0014_
rlabel metal2 27384 53256 27384 53256 0 _0015_
rlabel metal2 10808 35224 10808 35224 0 _0016_
rlabel metal2 12600 32872 12600 32872 0 _0017_
rlabel metal2 16688 30296 16688 30296 0 _0018_
rlabel metal2 20552 29736 20552 29736 0 _0019_
rlabel metal2 13496 29736 13496 29736 0 _0020_
rlabel metal2 9856 17752 9856 17752 0 _0021_
rlabel metal2 5432 14056 5432 14056 0 _0022_
rlabel metal2 6440 11480 6440 11480 0 _0023_
rlabel metal2 9912 11032 9912 11032 0 _0024_
rlabel metal2 11144 46872 11144 46872 0 _0025_
rlabel metal2 10472 49336 10472 49336 0 _0026_
rlabel metal2 3864 51800 3864 51800 0 _0027_
rlabel metal2 2856 58296 2856 58296 0 _0028_
rlabel metal2 2856 67396 2856 67396 0 _0029_
rlabel metal2 3640 65800 3640 65800 0 _0030_
rlabel metal2 6552 62664 6552 62664 0 _0031_
rlabel metal2 9240 58520 9240 58520 0 _0032_
rlabel metal2 10024 62776 10024 62776 0 _0033_
rlabel metal2 10808 71680 10808 71680 0 _0034_
rlabel metal2 12712 70840 12712 70840 0 _0035_
rlabel metal2 14728 58632 14728 58632 0 _0036_
rlabel metal2 18200 55384 18200 55384 0 _0037_
rlabel metal3 21784 52248 21784 52248 0 _0038_
rlabel metal2 24808 28840 24808 28840 0 _0039_
rlabel metal2 28168 28168 28168 28168 0 _0040_
rlabel metal2 30408 29736 30408 29736 0 _0041_
rlabel metal2 32592 33208 32592 33208 0 _0042_
rlabel metal2 27384 42784 27384 42784 0 _0043_
rlabel metal2 25368 48888 25368 48888 0 _0044_
rlabel metal2 25312 60984 25312 60984 0 _0045_
rlabel metal2 16296 69048 16296 69048 0 _0046_
rlabel metal2 17976 68264 17976 68264 0 _0047_
rlabel metal2 18648 63840 18648 63840 0 _0048_
rlabel metal2 18648 58576 18648 58576 0 _0049_
rlabel metal2 15176 53088 15176 53088 0 _0050_
rlabel metal2 2520 53256 2520 53256 0 _0051_
rlabel metal2 2800 56280 2800 56280 0 _0052_
rlabel metal2 2856 61824 2856 61824 0 _0053_
rlabel metal2 4648 59528 4648 59528 0 _0054_
rlabel metal2 6552 56000 6552 56000 0 _0055_
rlabel metal3 8232 54600 8232 54600 0 _0056_
rlabel metal2 2520 50680 2520 50680 0 _0057_
rlabel metal2 2968 44576 2968 44576 0 _0058_
rlabel metal2 2632 43876 2632 43876 0 _0059_
rlabel metal2 7336 43456 7336 43456 0 _0060_
rlabel metal2 10864 41272 10864 41272 0 _0061_
rlabel metal2 17752 38780 17752 38780 0 _0062_
rlabel metal3 25200 36344 25200 36344 0 _0063_
rlabel metal2 33880 31416 33880 31416 0 _0064_
rlabel metal2 37408 29512 37408 29512 0 _0065_
rlabel metal2 37408 37912 37408 37912 0 _0066_
rlabel metal2 37408 42056 37408 42056 0 _0067_
rlabel metal2 31752 43848 31752 43848 0 _0068_
rlabel metal3 32144 39704 32144 39704 0 _0069_
rlabel metal3 32200 34776 32200 34776 0 _0070_
rlabel metal2 37464 32872 37464 32872 0 _0071_
rlabel metal2 36456 36736 36456 36736 0 _0072_
rlabel metal2 34888 42392 34888 42392 0 _0073_
rlabel metal2 28224 45192 28224 45192 0 _0074_
rlabel metal2 29512 47712 29512 47712 0 _0075_
rlabel metal3 32088 47320 32088 47320 0 _0076_
rlabel metal3 36960 46760 36960 46760 0 _0077_
rlabel metal2 37408 48328 37408 48328 0 _0078_
rlabel metal2 33880 49504 33880 49504 0 _0079_
rlabel metal2 25592 49616 25592 49616 0 _0080_
rlabel metal2 27216 48440 27216 48440 0 _0081_
rlabel metal2 31248 52248 31248 52248 0 _0082_
rlabel metal2 33208 54208 33208 54208 0 _0083_
rlabel metal2 36344 53984 36344 53984 0 _0084_
rlabel metal2 37408 53032 37408 53032 0 _0085_
rlabel metal2 13496 53704 13496 53704 0 _0086_
rlabel metal2 10976 57848 10976 57848 0 _0087_
rlabel metal2 7112 65520 7112 65520 0 _0088_
rlabel metal2 7896 67928 7896 67928 0 _0089_
rlabel metal2 3304 69048 3304 69048 0 _0090_
rlabel metal2 6216 70504 6216 70504 0 _0091_
rlabel metal2 7560 71456 7560 71456 0 _0092_
rlabel metal2 11648 69272 11648 69272 0 _0093_
rlabel metal2 15960 70616 15960 70616 0 _0094_
rlabel metal3 19096 70056 19096 70056 0 _0095_
rlabel metal2 20832 67144 20832 67144 0 _0096_
rlabel metal2 22120 58632 22120 58632 0 _0097_
rlabel metal2 21616 38920 21616 38920 0 _0098_
rlabel metal2 15512 38668 15512 38668 0 _0099_
rlabel metal2 12824 36568 12824 36568 0 _0100_
rlabel metal2 15344 33432 15344 33432 0 _0101_
rlabel metal2 18648 33824 18648 33824 0 _0102_
rlabel metal3 22456 31864 22456 31864 0 _0103_
rlabel metal2 22400 27944 22400 27944 0 _0104_
rlabel metal2 23464 18368 23464 18368 0 _0105_
rlabel metal2 23912 10528 23912 10528 0 _0106_
rlabel metal2 27888 7560 27888 7560 0 _0107_
rlabel metal2 30856 7728 30856 7728 0 _0108_
rlabel metal2 31416 11032 31416 11032 0 _0109_
rlabel metal2 25928 18312 25928 18312 0 _0110_
rlabel metal3 10136 37912 10136 37912 0 _0111_
rlabel metal2 2520 37576 2520 37576 0 _0112_
rlabel metal2 2520 34440 2520 34440 0 _0113_
rlabel metal2 7560 35392 7560 35392 0 _0114_
rlabel metal2 10472 39648 10472 39648 0 _0115_
rlabel metal2 12376 43008 12376 43008 0 _0116_
rlabel metal2 12152 58128 12152 58128 0 _0117_
rlabel metal2 12152 64232 12152 64232 0 _0118_
rlabel metal2 13608 65072 13608 65072 0 _0119_
rlabel metal2 14280 60704 14280 60704 0 _0120_
rlabel metal2 13048 55608 13048 55608 0 _0121_
rlabel metal2 13608 49392 13608 49392 0 _0122_
rlabel metal3 15792 19320 15792 19320 0 _0123_
rlabel metal2 12992 10696 12992 10696 0 _0124_
rlabel metal2 14336 9912 14336 9912 0 _0125_
rlabel metal2 15736 10248 15736 10248 0 _0126_
rlabel metal2 17920 15960 17920 15960 0 _0127_
rlabel metal2 15064 26712 15064 26712 0 _0128_
rlabel metal2 8344 26684 8344 26684 0 _0129_
rlabel metal2 2632 23576 2632 23576 0 _0130_
rlabel metal2 3304 20132 3304 20132 0 _0131_
rlabel metal2 7000 21056 7000 21056 0 _0132_
rlabel metal2 10024 24192 10024 24192 0 _0133_
rlabel metal2 14168 23464 14168 23464 0 _0134_
rlabel metal2 20776 24192 20776 24192 0 _0135_
rlabel metal2 27776 24808 27776 24808 0 _0136_
rlabel metal3 30856 23800 30856 23800 0 _0137_
rlabel metal2 35112 24416 35112 24416 0 _0138_
rlabel metal2 27384 23464 27384 23464 0 _0139_
rlabel metal2 25032 22568 25032 22568 0 _0140_
rlabel metal2 28392 19320 28392 19320 0 _0141_
rlabel metal2 31192 17864 31192 17864 0 _0142_
rlabel metal2 33824 16968 33824 16968 0 _0143_
rlabel metal2 37352 19488 37352 19488 0 _0144_
rlabel metal2 31528 21056 31528 21056 0 _0145_
rlabel metal2 22680 23296 22680 23296 0 _0146_
rlabel metal2 20048 17752 20048 17752 0 _0147_
rlabel metal2 21224 8344 21224 8344 0 _0148_
rlabel metal2 19656 5152 19656 5152 0 _0149_
rlabel metal2 22120 4648 22120 4648 0 _0150_
rlabel metal2 22568 11648 22568 11648 0 _0151_
rlabel metal2 21896 17192 21896 17192 0 _0152_
rlabel metal2 22680 15260 22680 15260 0 _0153_
rlabel metal2 23856 3640 23856 3640 0 _0154_
rlabel metal2 24696 4760 24696 4760 0 _0155_
rlabel metal2 25816 8512 25816 8512 0 _0156_
rlabel metal2 28056 11648 28056 11648 0 _0157_
rlabel metal2 27384 15736 27384 15736 0 _0158_
rlabel metal2 29680 14392 29680 14392 0 _0159_
rlabel metal2 33096 14168 33096 14168 0 _0160_
rlabel metal2 36680 17696 36680 17696 0 _0161_
rlabel metal2 36120 21056 36120 21056 0 _0162_
rlabel metal2 35784 25032 35784 25032 0 _0163_
rlabel metal2 24584 34552 24584 34552 0 _0164_
rlabel metal2 23912 56504 23912 56504 0 _0165_
rlabel metal2 22680 65912 22680 65912 0 _0166_
rlabel metal2 25592 66920 25592 66920 0 _0167_
rlabel metal2 25928 62300 25928 62300 0 _0168_
rlabel metal2 24584 57344 24584 57344 0 _0169_
rlabel metal3 24808 39704 24808 39704 0 _0170_
rlabel metal2 8176 27944 8176 27944 0 _0171_
rlabel metal2 2520 23632 2520 23632 0 _0172_
rlabel metal2 3304 17920 3304 17920 0 _0173_
rlabel metal2 6104 17192 6104 17192 0 _0174_
rlabel metal2 9576 22008 9576 22008 0 _0175_
rlabel metal2 11592 22456 11592 22456 0 _0176_
rlabel metal2 9352 17304 9352 17304 0 _0177_
rlabel metal2 8344 13440 8344 13440 0 _0178_
rlabel metal2 8008 7336 8008 7336 0 _0179_
rlabel metal2 10248 5768 10248 5768 0 _0180_
rlabel metal2 12096 4872 12096 4872 0 _0181_
rlabel metal2 12600 17192 12600 17192 0 _0182_
rlabel metal2 13944 16408 13944 16408 0 _0183_
rlabel metal2 14280 5376 14280 5376 0 _0184_
rlabel metal2 15848 4984 15848 4984 0 _0185_
rlabel metal2 17080 5600 17080 5600 0 _0186_
rlabel metal2 18200 20832 18200 20832 0 _0187_
rlabel metal3 19096 22232 19096 22232 0 _0188_
rlabel metal2 2632 26152 2632 26152 0 _0189_
rlabel metal2 3080 28896 3080 28896 0 _0190_
rlabel metal2 3528 30464 3528 30464 0 _0191_
rlabel metal2 6776 42224 6776 42224 0 _0192_
rlabel metal2 7448 47096 7448 47096 0 _0193_
rlabel metal2 6776 48552 6776 48552 0 _0194_
rlabel metal2 2968 47936 2968 47936 0 _0195_
rlabel metal2 2520 39144 2520 39144 0 _0196_
rlabel metal2 4648 33096 4648 33096 0 _0197_
rlabel metal2 8008 31416 8008 31416 0 _0198_
rlabel metal2 10864 28728 10864 28728 0 _0199_
rlabel metal2 17752 27272 17752 27272 0 _0200_
rlabel metal2 17752 78456 17752 78456 0 _0201_
rlabel metal2 14056 78456 14056 78456 0 _0202_
rlabel metal2 12264 76608 12264 76608 0 _0203_
rlabel metal3 16800 75096 16800 75096 0 _0204_
rlabel metal3 18928 74760 18928 74760 0 _0205_
rlabel metal2 22568 72296 22568 72296 0 _0206_
rlabel metal2 18256 81256 18256 81256 0 _0207_
rlabel metal2 19544 88536 19544 88536 0 _0208_
rlabel metal2 18144 82040 18144 82040 0 _0209_
rlabel metal2 11368 79912 11368 79912 0 _0210_
rlabel metal2 12712 83048 12712 83048 0 _0211_
rlabel metal2 14728 84616 14728 84616 0 _0212_
rlabel metal2 14056 88536 14056 88536 0 _0213_
rlabel metal3 16856 88312 16856 88312 0 _0214_
rlabel metal2 24360 87584 24360 87584 0 _0215_
rlabel metal2 30016 88312 30016 88312 0 _0216_
rlabel metal2 31752 85848 31752 85848 0 _0217_
rlabel metal2 35000 87024 35000 87024 0 _0218_
rlabel metal2 35560 87528 35560 87528 0 _0219_
rlabel metal3 36624 83720 36624 83720 0 _0220_
rlabel metal2 36344 84224 36344 84224 0 _0221_
rlabel metal2 3080 56112 3080 56112 0 _0222_
rlabel metal2 3192 67452 3192 67452 0 _0223_
rlabel metal2 3864 65072 3864 65072 0 _0224_
rlabel metal2 6440 62580 6440 62580 0 _0225_
rlabel metal2 10080 59416 10080 59416 0 _0226_
rlabel metal2 10360 61656 10360 61656 0 _0227_
rlabel metal2 11592 71120 11592 71120 0 _0228_
rlabel metal2 13552 71176 13552 71176 0 _0229_
rlabel metal2 15736 59136 15736 59136 0 _0230_
rlabel metal2 17528 56392 17528 56392 0 _0231_
rlabel metal2 21336 54208 21336 54208 0 _0232_
rlabel metal2 24136 30464 24136 30464 0 _0233_
rlabel metal2 28112 28616 28112 28616 0 _0234_
rlabel metal2 30464 28840 30464 28840 0 _0235_
rlabel metal2 32200 31696 32200 31696 0 _0236_
rlabel metal2 26600 40544 26600 40544 0 _0237_
rlabel metal2 26264 47096 26264 47096 0 _0238_
rlabel metal2 25368 60480 25368 60480 0 _0239_
rlabel metal3 17752 53032 17752 53032 0 _0240_
rlabel metal2 6328 53368 6328 53368 0 _0241_
rlabel metal2 3192 55384 3192 55384 0 _0242_
rlabel metal3 18312 38696 18312 38696 0 _0243_
rlabel metal2 3416 61208 3416 61208 0 _0244_
rlabel metal3 5376 59976 5376 59976 0 _0245_
rlabel metal2 6776 56840 6776 56840 0 _0246_
rlabel metal2 8568 53984 8568 53984 0 _0247_
rlabel metal2 3528 52080 3528 52080 0 _0248_
rlabel metal2 3304 44968 3304 44968 0 _0249_
rlabel metal3 2968 44296 2968 44296 0 _0250_
rlabel metal3 6440 42952 6440 42952 0 _0251_
rlabel metal2 22680 40936 22680 40936 0 _0252_
rlabel metal2 10584 41888 10584 41888 0 _0253_
rlabel metal2 17416 39536 17416 39536 0 _0254_
rlabel metal3 23520 36456 23520 36456 0 _0255_
rlabel metal3 32480 32648 32480 32648 0 _0256_
rlabel metal3 36624 31640 36624 31640 0 _0257_
rlabel metal2 37576 37296 37576 37296 0 _0258_
rlabel metal2 36456 42000 36456 42000 0 _0259_
rlabel metal3 31080 42952 31080 42952 0 _0260_
rlabel metal2 31584 41160 31584 41160 0 _0261_
rlabel metal2 31416 35168 31416 35168 0 _0262_
rlabel metal3 36456 33208 36456 33208 0 _0263_
rlabel metal2 36400 35896 36400 35896 0 _0264_
rlabel metal2 35000 41664 35000 41664 0 _0265_
rlabel metal2 29624 47152 29624 47152 0 _0266_
rlabel metal2 31304 47544 31304 47544 0 _0267_
rlabel metal2 36232 47376 36232 47376 0 _0268_
rlabel metal2 37576 46648 37576 46648 0 _0269_
rlabel metal2 33992 49728 33992 49728 0 _0270_
rlabel metal2 24248 49112 24248 49112 0 _0271_
rlabel metal2 26824 48440 26824 48440 0 _0272_
rlabel metal2 30744 52248 30744 52248 0 _0273_
rlabel metal2 33208 53144 33208 53144 0 _0274_
rlabel metal2 35952 52360 35952 52360 0 _0275_
rlabel metal2 37016 52976 37016 52976 0 _0276_
rlabel metal2 12376 53368 12376 53368 0 _0277_
rlabel metal2 11256 56504 11256 56504 0 _0278_
rlabel metal2 7896 65184 7896 65184 0 _0279_
rlabel metal2 8400 66920 8400 66920 0 _0280_
rlabel metal2 3864 68544 3864 68544 0 _0281_
rlabel metal2 5656 70224 5656 70224 0 _0282_
rlabel metal2 9128 70672 9128 70672 0 _0283_
rlabel metal2 11256 69552 11256 69552 0 _0284_
rlabel metal2 20888 40712 20888 40712 0 _0285_
rlabel metal3 17584 38808 17584 38808 0 _0286_
rlabel metal2 18536 23632 18536 23632 0 _0287_
rlabel metal2 13832 37408 13832 37408 0 _0288_
rlabel metal2 15064 34440 15064 34440 0 _0289_
rlabel metal2 18424 33432 18424 33432 0 _0290_
rlabel metal3 21896 22456 21896 22456 0 _0291_
rlabel metal2 21224 32816 21224 32816 0 _0292_
rlabel metal2 22792 29736 22792 29736 0 _0293_
rlabel metal2 23296 19208 23296 19208 0 _0294_
rlabel metal2 24360 12040 24360 12040 0 _0295_
rlabel metal2 26712 7728 26712 7728 0 _0296_
rlabel metal2 30632 7728 30632 7728 0 _0297_
rlabel metal2 31192 10304 31192 10304 0 _0298_
rlabel metal2 25984 17080 25984 17080 0 _0299_
rlabel metal2 20776 37744 20776 37744 0 _0300_
rlabel metal2 3304 37856 3304 37856 0 _0301_
rlabel metal2 3304 35168 3304 35168 0 _0302_
rlabel metal2 6552 33712 6552 33712 0 _0303_
rlabel metal2 10136 38136 10136 38136 0 _0304_
rlabel metal2 12600 42448 12600 42448 0 _0305_
rlabel metal2 13496 47488 13496 47488 0 _0306_
rlabel metal2 13832 13608 13832 13608 0 _0307_
rlabel metal2 15400 11424 15400 11424 0 _0308_
rlabel metal2 15512 8960 15512 8960 0 _0309_
rlabel metal2 17640 14224 17640 14224 0 _0310_
rlabel metal3 15344 26264 15344 26264 0 _0311_
rlabel metal3 8848 27608 8848 27608 0 _0312_
rlabel metal2 4312 25032 4312 25032 0 _0313_
rlabel metal2 4200 21224 4200 21224 0 _0314_
rlabel metal2 6496 20664 6496 20664 0 _0315_
rlabel metal2 10136 23408 10136 23408 0 _0316_
rlabel metal2 13608 24192 13608 24192 0 _0317_
rlabel metal2 20440 23744 20440 23744 0 _0318_
rlabel metal2 27048 25312 27048 25312 0 _0319_
rlabel metal2 31416 24640 31416 24640 0 _0320_
rlabel metal2 33096 24640 33096 24640 0 _0321_
rlabel metal3 28616 23352 28616 23352 0 _0322_
rlabel metal2 24472 23520 24472 23520 0 _0323_
rlabel metal2 27832 20328 27832 20328 0 _0324_
rlabel metal2 32088 18368 32088 18368 0 _0325_
rlabel metal2 33600 17864 33600 17864 0 _0326_
rlabel metal2 37016 19040 37016 19040 0 _0327_
rlabel metal2 31864 21056 31864 21056 0 _0328_
rlabel metal2 21896 23240 21896 23240 0 _0329_
rlabel metal2 21000 20944 21000 20944 0 _0330_
rlabel metal2 20328 9296 20328 9296 0 _0331_
rlabel metal2 19432 4592 19432 4592 0 _0332_
rlabel metal2 22176 5096 22176 5096 0 _0333_
rlabel metal2 22904 18144 22904 18144 0 _0334_
rlabel metal2 22456 11088 22456 11088 0 _0335_
rlabel metal2 21336 16520 21336 16520 0 _0336_
rlabel metal2 22456 15568 22456 15568 0 _0337_
rlabel metal2 23576 5376 23576 5376 0 _0338_
rlabel metal2 24472 4704 24472 4704 0 _0339_
rlabel metal3 26320 8232 26320 8232 0 _0340_
rlabel metal2 27496 11032 27496 11032 0 _0341_
rlabel metal2 27160 15204 27160 15204 0 _0342_
rlabel metal2 29176 15484 29176 15484 0 _0343_
rlabel metal2 33320 14000 33320 14000 0 _0344_
rlabel metal2 35560 16352 35560 16352 0 _0345_
rlabel metal2 36064 19432 36064 19432 0 _0346_
rlabel metal2 36120 24360 36120 24360 0 _0347_
rlabel metal2 24080 34104 24080 34104 0 _0348_
rlabel metal2 23912 55384 23912 55384 0 _0349_
rlabel metal2 23016 65184 23016 65184 0 _0350_
rlabel metal2 25816 65744 25816 65744 0 _0351_
rlabel metal2 25704 63392 25704 63392 0 _0352_
rlabel metal2 24192 57736 24192 57736 0 _0353_
rlabel metal2 23800 29008 23800 29008 0 _0354_
rlabel metal3 17920 23016 17920 23016 0 _0355_
rlabel metal2 3640 25424 3640 25424 0 _0356_
rlabel metal2 3640 18312 3640 18312 0 _0357_
rlabel metal2 6496 17640 6496 17640 0 _0358_
rlabel metal2 9016 21280 9016 21280 0 _0359_
rlabel metal2 11816 22848 11816 22848 0 _0360_
rlabel metal2 10696 18816 10696 18816 0 _0361_
rlabel metal2 9912 14448 9912 14448 0 _0362_
rlabel metal2 9016 8232 9016 8232 0 _0363_
rlabel metal3 10248 6664 10248 6664 0 _0364_
rlabel metal2 12152 5768 12152 5768 0 _0365_
rlabel metal2 13552 16296 13552 16296 0 _0366_
rlabel metal2 15064 17136 15064 17136 0 _0367_
rlabel metal2 14504 5768 14504 5768 0 _0368_
rlabel metal2 15904 4312 15904 4312 0 _0369_
rlabel metal2 17472 4536 17472 4536 0 _0370_
rlabel metal2 17752 19320 17752 19320 0 _0371_
rlabel metal2 19992 22456 19992 22456 0 _0372_
rlabel metal3 4872 24136 4872 24136 0 _0373_
rlabel metal2 3640 28616 3640 28616 0 _0374_
rlabel metal2 4872 29624 4872 29624 0 _0375_
rlabel metal2 6552 41440 6552 41440 0 _0376_
rlabel metal2 8008 45976 8008 45976 0 _0377_
rlabel metal2 7280 48888 7280 48888 0 _0378_
rlabel metal2 4424 48216 4424 48216 0 _0379_
rlabel metal2 3192 39984 3192 39984 0 _0380_
rlabel metal2 5208 34776 5208 34776 0 _0381_
rlabel metal2 7672 31696 7672 31696 0 _0382_
rlabel metal2 10696 30464 10696 30464 0 _0383_
rlabel metal3 17024 26488 17024 26488 0 _0384_
rlabel metal2 19880 83720 19880 83720 0 _0385_
rlabel metal2 16520 80808 16520 80808 0 _0386_
rlabel metal2 16744 79240 16744 79240 0 _0387_
rlabel metal2 16744 77336 16744 77336 0 _0388_
rlabel metal2 15064 78064 15064 78064 0 _0389_
rlabel metal3 13384 77336 13384 77336 0 _0390_
rlabel metal2 17864 74984 17864 74984 0 _0391_
rlabel metal2 19992 74256 19992 74256 0 _0392_
rlabel metal3 23464 74872 23464 74872 0 _0393_
rlabel metal2 19432 83440 19432 83440 0 _0394_
rlabel metal2 12264 79968 12264 79968 0 _0395_
rlabel metal2 11928 79632 11928 79632 0 _0396_
rlabel metal2 15176 82880 15176 82880 0 _0397_
rlabel metal2 14280 85400 14280 85400 0 _0398_
rlabel metal2 14392 88032 14392 88032 0 _0399_
rlabel metal2 15792 87192 15792 87192 0 _0400_
rlabel metal2 16856 87864 16856 87864 0 _0401_
rlabel metal3 25648 87416 25648 87416 0 _0402_
rlabel metal2 30296 90272 30296 90272 0 _0403_
rlabel metal2 31528 85876 31528 85876 0 _0404_
rlabel metal3 33264 86072 33264 86072 0 _0405_
rlabel metal2 35728 88088 35728 88088 0 _0406_
rlabel metal2 36008 83944 36008 83944 0 _0407_
rlabel metal3 36624 83384 36624 83384 0 _0408_
rlabel metal3 36120 83272 36120 83272 0 _0409_
rlabel metal2 34776 84056 34776 84056 0 _0410_
rlabel metal2 36064 85848 36064 85848 0 _0411_
rlabel metal2 29344 86408 29344 86408 0 _0412_
rlabel metal3 20664 87640 20664 87640 0 _0413_
rlabel metal2 20272 87976 20272 87976 0 _0414_
rlabel metal2 21560 80080 21560 80080 0 _0415_
rlabel metal2 22792 90440 22792 90440 0 _0416_
rlabel metal2 20272 84280 20272 84280 0 _0417_
rlabel metal2 15400 83608 15400 83608 0 _0418_
rlabel metal3 16744 87416 16744 87416 0 _0419_
rlabel metal2 27384 88872 27384 88872 0 _0420_
rlabel metal2 31192 87584 31192 87584 0 _0421_
rlabel metal2 31808 87192 31808 87192 0 _0422_
rlabel metal2 33544 85848 33544 85848 0 _0423_
rlabel metal2 35056 84504 35056 84504 0 _0424_
rlabel metal2 24248 46928 24248 46928 0 _0425_
rlabel metal2 22680 48888 22680 48888 0 _0426_
rlabel metal2 30408 67088 30408 67088 0 _0427_
rlabel metal2 20720 44408 20720 44408 0 _0428_
rlabel metal2 24696 48496 24696 48496 0 _0429_
rlabel metal2 29176 64064 29176 64064 0 _0430_
rlabel metal2 32872 35840 32872 35840 0 _0431_
rlabel metal3 23632 48888 23632 48888 0 _0432_
rlabel metal2 22120 41720 22120 41720 0 _0433_
rlabel metal2 23576 47936 23576 47936 0 _0434_
rlabel metal2 24248 41888 24248 41888 0 _0435_
rlabel metal2 21784 44352 21784 44352 0 _0436_
rlabel metal2 19264 21000 19264 21000 0 _0437_
rlabel metal2 21224 62328 21224 62328 0 _0438_
rlabel metal2 26264 42392 26264 42392 0 _0439_
rlabel metal2 25480 23576 25480 23576 0 _0440_
rlabel metal2 19096 42896 19096 42896 0 _0441_
rlabel metal2 16408 40880 16408 40880 0 _0442_
rlabel metal2 18200 66304 18200 66304 0 _0443_
rlabel metal2 22792 23156 22792 23156 0 _0444_
rlabel metal2 30744 21112 30744 21112 0 _0445_
rlabel via2 33768 34776 33768 34776 0 _0446_
rlabel metal3 24248 63952 24248 63952 0 _0447_
rlabel metal2 26600 45136 26600 45136 0 _0448_
rlabel metal3 29176 44072 29176 44072 0 _0449_
rlabel metal2 31024 34216 31024 34216 0 _0450_
rlabel metal2 18032 48328 18032 48328 0 _0451_
rlabel metal2 19432 48832 19432 48832 0 _0452_
rlabel metal2 16016 45864 16016 45864 0 _0453_
rlabel metal2 22512 53592 22512 53592 0 _0454_
rlabel metal2 31360 41832 31360 41832 0 _0455_
rlabel metal2 24696 45024 24696 45024 0 _0456_
rlabel metal2 26432 26152 26432 26152 0 _0457_
rlabel metal2 27496 29288 27496 29288 0 _0458_
rlabel metal2 23520 26488 23520 26488 0 _0459_
rlabel metal2 26712 28448 26712 28448 0 _0460_
rlabel metal2 28168 31864 28168 31864 0 _0461_
rlabel metal3 31080 34328 31080 34328 0 _0462_
rlabel metal2 20216 48664 20216 48664 0 _0463_
rlabel metal2 17528 40488 17528 40488 0 _0464_
rlabel metal2 17640 41552 17640 41552 0 _0465_
rlabel metal3 16408 40936 16408 40936 0 _0466_
rlabel metal3 16184 38136 16184 38136 0 _0467_
rlabel metal2 16520 40712 16520 40712 0 _0468_
rlabel metal3 16744 42560 16744 42560 0 _0469_
rlabel metal2 5824 38808 5824 38808 0 _0470_
rlabel metal2 17080 50176 17080 50176 0 _0471_
rlabel metal2 17528 45752 17528 45752 0 _0472_
rlabel metal2 5992 39536 5992 39536 0 _0473_
rlabel metal2 15176 22904 15176 22904 0 _0474_
rlabel metal2 23800 45136 23800 45136 0 _0475_
rlabel metal3 16296 22120 16296 22120 0 _0476_
rlabel metal2 6608 28728 6608 28728 0 _0477_
rlabel metal2 17080 48720 17080 48720 0 _0478_
rlabel metal3 11256 42504 11256 42504 0 _0479_
rlabel metal2 6440 39256 6440 39256 0 _0480_
rlabel metal2 16632 37856 16632 37856 0 _0481_
rlabel metal2 13720 62832 13720 62832 0 _0482_
rlabel metal2 14056 63672 14056 63672 0 _0483_
rlabel metal3 22400 63896 22400 63896 0 _0484_
rlabel metal2 17976 66192 17976 66192 0 _0485_
rlabel metal2 19320 66640 19320 66640 0 _0486_
rlabel metal3 16184 70280 16184 70280 0 _0487_
rlabel metal2 17416 65184 17416 65184 0 _0488_
rlabel metal2 14392 64176 14392 64176 0 _0489_
rlabel metal2 16520 49560 16520 49560 0 _0490_
rlabel metal2 15176 63616 15176 63616 0 _0491_
rlabel metal2 16408 63952 16408 63952 0 _0492_
rlabel metal2 18872 43960 18872 43960 0 _0493_
rlabel metal2 19992 18480 19992 18480 0 _0494_
rlabel metal3 18872 15176 18872 15176 0 _0495_
rlabel metal2 23912 16744 23912 16744 0 _0496_
rlabel metal2 25368 16296 25368 16296 0 _0497_
rlabel metal2 18200 15344 18200 15344 0 _0498_
rlabel metal2 15904 21784 15904 21784 0 _0499_
rlabel metal2 11984 16072 11984 16072 0 _0500_
rlabel metal2 12152 15624 12152 15624 0 _0501_
rlabel metal2 19544 23856 19544 23856 0 _0502_
rlabel metal2 17528 19376 17528 19376 0 _0503_
rlabel metal2 17472 15288 17472 15288 0 _0504_
rlabel metal2 17080 37576 17080 37576 0 _0505_
rlabel metal3 22120 37688 22120 37688 0 _0506_
rlabel metal3 31528 65352 31528 65352 0 _0507_
rlabel metal2 29624 65184 29624 65184 0 _0508_
rlabel metal2 29344 33544 29344 33544 0 _0509_
rlabel metal2 33992 23100 33992 23100 0 _0510_
rlabel metal2 33992 33600 33992 33600 0 _0511_
rlabel metal2 33992 43372 33992 43372 0 _0512_
rlabel metal2 31864 29344 31864 29344 0 _0513_
rlabel metal2 31584 27272 31584 27272 0 _0514_
rlabel metal2 32424 29736 32424 29736 0 _0515_
rlabel metal3 33096 33488 33096 33488 0 _0516_
rlabel metal3 16632 35560 16632 35560 0 _0517_
rlabel metal2 5992 36624 5992 36624 0 _0518_
rlabel metal3 4760 37240 4760 37240 0 _0519_
rlabel metal2 5432 23352 5432 23352 0 _0520_
rlabel metal3 5376 38584 5376 38584 0 _0521_
rlabel metal2 6440 36400 6440 36400 0 _0522_
rlabel metal2 20552 65800 20552 65800 0 _0523_
rlabel metal3 22232 65464 22232 65464 0 _0524_
rlabel metal2 17864 68432 17864 68432 0 _0525_
rlabel metal2 18592 70280 18592 70280 0 _0526_
rlabel metal2 19096 66136 19096 66136 0 _0527_
rlabel metal2 14112 66024 14112 66024 0 _0528_
rlabel metal2 15064 65184 15064 65184 0 _0529_
rlabel metal3 16912 65576 16912 65576 0 _0530_
rlabel metal2 18592 39368 18592 39368 0 _0531_
rlabel metal3 19488 10808 19488 10808 0 _0532_
rlabel metal2 25312 10472 25312 10472 0 _0533_
rlabel metal2 17976 11984 17976 11984 0 _0534_
rlabel metal3 16912 12152 16912 12152 0 _0535_
rlabel metal3 17528 35672 17528 35672 0 _0536_
rlabel metal2 27384 34832 27384 34832 0 _0537_
rlabel metal2 29288 45864 29288 45864 0 _0538_
rlabel metal2 29624 60480 29624 60480 0 _0539_
rlabel metal2 28504 36176 28504 36176 0 _0540_
rlabel metal3 35504 20104 35504 20104 0 _0541_
rlabel metal2 35448 34608 35448 34608 0 _0542_
rlabel metal3 36232 42952 36232 42952 0 _0543_
rlabel metal2 33096 29680 33096 29680 0 _0544_
rlabel metal2 32648 28616 32648 28616 0 _0545_
rlabel metal2 33768 29624 33768 29624 0 _0546_
rlabel metal2 34552 34496 34552 34496 0 _0547_
rlabel metal2 17752 34608 17752 34608 0 _0548_
rlabel metal2 6104 34384 6104 34384 0 _0549_
rlabel metal2 6552 40936 6552 40936 0 _0550_
rlabel metal2 6384 22456 6384 22456 0 _0551_
rlabel metal2 6384 40040 6384 40040 0 _0552_
rlabel metal2 18088 34552 18088 34552 0 _0553_
rlabel metal2 19544 65128 19544 65128 0 _0554_
rlabel metal3 22456 64680 22456 64680 0 _0555_
rlabel metal2 19432 65800 19432 65800 0 _0556_
rlabel metal2 20664 68040 20664 68040 0 _0557_
rlabel metal2 18648 65576 18648 65576 0 _0558_
rlabel metal2 14672 63672 14672 63672 0 _0559_
rlabel metal2 16520 62608 16520 62608 0 _0560_
rlabel metal2 16632 63336 16632 63336 0 _0561_
rlabel metal3 18928 34776 18928 34776 0 _0562_
rlabel metal2 18872 10640 18872 10640 0 _0563_
rlabel metal3 22568 9912 22568 9912 0 _0564_
rlabel metal2 11032 10248 11032 10248 0 _0565_
rlabel metal2 17640 10080 17640 10080 0 _0566_
rlabel metal2 19488 21000 19488 21000 0 _0567_
rlabel metal2 27048 35168 27048 35168 0 _0568_
rlabel metal2 28784 58632 28784 58632 0 _0569_
rlabel metal3 29568 59976 29568 59976 0 _0570_
rlabel metal2 29736 40488 29736 40488 0 _0571_
rlabel metal2 34888 23408 34888 23408 0 _0572_
rlabel metal2 35224 39592 35224 39592 0 _0573_
rlabel metal2 35000 39928 35000 39928 0 _0574_
rlabel metal2 32816 38696 32816 38696 0 _0575_
rlabel metal2 33320 38416 33320 38416 0 _0576_
rlabel metal2 33656 39424 33656 39424 0 _0577_
rlabel metal3 32424 39816 32424 39816 0 _0578_
rlabel metal2 19544 35000 19544 35000 0 _0579_
rlabel metal2 9016 36176 9016 36176 0 _0580_
rlabel metal3 8064 36568 8064 36568 0 _0581_
rlabel metal2 8960 31640 8960 31640 0 _0582_
rlabel metal3 9744 42504 9744 42504 0 _0583_
rlabel metal2 19712 35784 19712 35784 0 _0584_
rlabel metal3 20160 59416 20160 59416 0 _0585_
rlabel metal2 22792 59472 22792 59472 0 _0586_
rlabel metal2 19432 60424 19432 60424 0 _0587_
rlabel metal2 21784 63700 21784 63700 0 _0588_
rlabel metal2 19096 59696 19096 59696 0 _0589_
rlabel metal2 16072 58296 16072 58296 0 _0590_
rlabel metal2 18088 58520 18088 58520 0 _0591_
rlabel metal3 18536 59304 18536 59304 0 _0592_
rlabel metal2 20944 35896 20944 35896 0 _0593_
rlabel metal3 20832 11368 20832 11368 0 _0594_
rlabel metal2 26824 11032 26824 11032 0 _0595_
rlabel metal2 19768 11424 19768 11424 0 _0596_
rlabel metal2 19656 11648 19656 11648 0 _0597_
rlabel metal2 18816 21000 18816 21000 0 _0598_
rlabel metal2 20552 36288 20552 36288 0 _0599_
rlabel metal2 29008 43176 29008 43176 0 _0600_
rlabel metal3 30464 58520 30464 58520 0 _0601_
rlabel metal3 30688 54712 30688 54712 0 _0602_
rlabel metal2 19656 24696 19656 24696 0 _0603_
rlabel metal2 22008 24472 22008 24472 0 _0604_
rlabel metal2 25144 29232 25144 29232 0 _0605_
rlabel metal3 23352 26376 23352 26376 0 _0606_
rlabel metal2 24472 25760 24472 25760 0 _0607_
rlabel metal3 25144 39480 25144 39480 0 _0608_
rlabel metal3 21672 27944 21672 27944 0 _0609_
rlabel metal3 26152 26488 26152 26488 0 _0610_
rlabel metal2 25648 39592 25648 39592 0 _0611_
rlabel metal3 31360 42728 31360 42728 0 _0612_
rlabel metal2 27272 44240 27272 44240 0 _0613_
rlabel metal2 26824 42280 26824 42280 0 _0614_
rlabel metal2 28056 18312 28056 18312 0 _0615_
rlabel metal2 27160 42280 27160 42280 0 _0616_
rlabel metal2 25648 48440 25648 48440 0 _0617_
rlabel metal2 25144 42056 25144 42056 0 _0618_
rlabel metal2 26152 31864 26152 31864 0 _0619_
rlabel metal3 20216 39256 20216 39256 0 _0620_
rlabel metal2 26040 39200 26040 39200 0 _0621_
rlabel metal2 30128 46760 30128 46760 0 _0622_
rlabel metal2 15960 49392 15960 49392 0 _0623_
rlabel metal2 14504 49112 14504 49112 0 _0624_
rlabel metal2 15512 48664 15512 48664 0 _0625_
rlabel metal3 18928 50904 18928 50904 0 _0626_
rlabel metal2 22232 44744 22232 44744 0 _0627_
rlabel metal2 19992 51464 19992 51464 0 _0628_
rlabel metal2 19264 45304 19264 45304 0 _0629_
rlabel metal2 20440 52024 20440 52024 0 _0630_
rlabel metal2 20776 51352 20776 51352 0 _0631_
rlabel metal2 22120 53256 22120 53256 0 _0632_
rlabel metal2 22624 46984 22624 46984 0 _0633_
rlabel metal2 22008 51800 22008 51800 0 _0634_
rlabel metal2 22456 52248 22456 52248 0 _0635_
rlabel metal3 21840 41160 21840 41160 0 _0636_
rlabel metal2 21448 42560 21448 42560 0 _0637_
rlabel metal2 17864 48328 17864 48328 0 _0638_
rlabel metal3 22064 51464 22064 51464 0 _0639_
rlabel metal2 24584 52864 24584 52864 0 _0640_
rlabel metal2 30016 64120 30016 64120 0 _0641_
rlabel metal3 29064 64904 29064 64904 0 _0642_
rlabel metal3 30184 62552 30184 62552 0 _0643_
rlabel metal2 16072 22232 16072 22232 0 _0644_
rlabel metal2 15624 23184 15624 23184 0 _0645_
rlabel metal3 16744 47208 16744 47208 0 _0646_
rlabel metal2 16296 52416 16296 52416 0 _0647_
rlabel metal2 15736 50960 15736 50960 0 _0648_
rlabel metal2 15624 49896 15624 49896 0 _0649_
rlabel metal3 17248 50344 17248 50344 0 _0650_
rlabel metal2 14728 47824 14728 47824 0 _0651_
rlabel metal3 21112 26824 21112 26824 0 _0652_
rlabel metal2 16408 48664 16408 48664 0 _0653_
rlabel metal2 16520 47768 16520 47768 0 _0654_
rlabel metal2 19824 18200 19824 18200 0 _0655_
rlabel metal2 15456 42616 15456 42616 0 _0656_
rlabel metal2 15736 32452 15736 32452 0 _0657_
rlabel metal2 16296 43848 16296 43848 0 _0658_
rlabel metal2 26936 48384 26936 48384 0 _0659_
rlabel metal2 22232 38388 22232 38388 0 _0660_
rlabel metal2 22456 39592 22456 39592 0 _0661_
rlabel metal2 22792 42672 22792 42672 0 _0662_
rlabel metal2 21560 44128 21560 44128 0 _0663_
rlabel metal2 22960 41832 22960 41832 0 _0664_
rlabel metal3 23352 44408 23352 44408 0 _0665_
rlabel metal2 23800 39984 23800 39984 0 _0666_
rlabel metal2 25480 41496 25480 41496 0 _0667_
rlabel metal2 24248 39480 24248 39480 0 _0668_
rlabel metal2 26264 44688 26264 44688 0 _0669_
rlabel metal2 23688 45864 23688 45864 0 _0670_
rlabel metal2 23576 45136 23576 45136 0 _0671_
rlabel metal3 25368 45752 25368 45752 0 _0672_
rlabel metal2 27944 56728 27944 56728 0 _0673_
rlabel metal2 31080 57456 31080 57456 0 _0674_
rlabel metal2 19544 83384 19544 83384 0 _0675_
rlabel metal2 32256 81816 32256 81816 0 _0676_
rlabel metal2 24248 84504 24248 84504 0 _0677_
rlabel metal2 22904 83216 22904 83216 0 _0678_
rlabel metal2 22792 86688 22792 86688 0 _0679_
rlabel metal2 21784 88984 21784 88984 0 _0680_
rlabel metal2 22120 88760 22120 88760 0 _0681_
rlabel metal2 26152 73192 26152 73192 0 _0682_
rlabel metal2 26264 70560 26264 70560 0 _0683_
rlabel metal2 26152 69776 26152 69776 0 _0684_
rlabel metal2 26544 70392 26544 70392 0 _0685_
rlabel metal2 27048 82544 27048 82544 0 _0686_
rlabel metal2 26824 69776 26824 69776 0 _0687_
rlabel metal3 27272 73192 27272 73192 0 _0688_
rlabel metal2 25816 76384 25816 76384 0 _0689_
rlabel metal3 28728 73304 28728 73304 0 _0690_
rlabel metal2 25256 76272 25256 76272 0 _0691_
rlabel metal2 27944 72324 27944 72324 0 _0692_
rlabel metal2 28616 68264 28616 68264 0 _0693_
rlabel metal2 30296 69664 30296 69664 0 _0694_
rlabel metal2 31696 69384 31696 69384 0 _0695_
rlabel metal3 33152 70168 33152 70168 0 _0696_
rlabel metal3 32984 70392 32984 70392 0 _0697_
rlabel metal2 28952 70728 28952 70728 0 _0698_
rlabel metal2 31528 78960 31528 78960 0 _0699_
rlabel metal2 30520 78848 30520 78848 0 _0700_
rlabel metal2 30184 72184 30184 72184 0 _0701_
rlabel metal2 29736 80752 29736 80752 0 _0702_
rlabel metal3 27832 81144 27832 81144 0 _0703_
rlabel metal2 29624 70280 29624 70280 0 _0704_
rlabel metal2 26488 74928 26488 74928 0 _0705_
rlabel metal2 27496 81312 27496 81312 0 _0706_
rlabel metal2 26600 82040 26600 82040 0 _0707_
rlabel metal3 28112 82936 28112 82936 0 _0708_
rlabel metal3 28560 83720 28560 83720 0 _0709_
rlabel metal3 29456 63896 29456 63896 0 _0710_
rlabel metal2 31024 64008 31024 64008 0 _0711_
rlabel metal2 31304 77280 31304 77280 0 _0712_
rlabel metal2 30072 77896 30072 77896 0 _0713_
rlabel metal3 28672 81256 28672 81256 0 _0714_
rlabel metal2 28280 82040 28280 82040 0 _0715_
rlabel metal3 24248 86072 24248 86072 0 _0716_
rlabel metal2 23744 86072 23744 86072 0 _0717_
rlabel metal2 27776 86408 27776 86408 0 _0718_
rlabel metal2 28896 84504 28896 84504 0 _0719_
rlabel metal2 22792 87696 22792 87696 0 _0720_
rlabel metal2 23184 86632 23184 86632 0 _0721_
rlabel metal3 22400 86408 22400 86408 0 _0722_
rlabel metal2 22344 84784 22344 84784 0 _0723_
rlabel metal3 23072 86184 23072 86184 0 _0724_
rlabel metal2 24752 95928 24752 95928 0 _0725_
rlabel metal2 28448 60536 28448 60536 0 _0726_
rlabel metal2 28728 70168 28728 70168 0 _0727_
rlabel metal3 30968 77224 30968 77224 0 _0728_
rlabel metal2 29400 78848 29400 78848 0 _0729_
rlabel metal2 28504 80640 28504 80640 0 _0730_
rlabel metal3 28672 78904 28672 78904 0 _0731_
rlabel metal2 27160 78792 27160 78792 0 _0732_
rlabel metal3 18312 79632 18312 79632 0 _0733_
rlabel metal3 21056 79576 21056 79576 0 _0734_
rlabel metal2 22568 87640 22568 87640 0 _0735_
rlabel metal2 18424 79128 18424 79128 0 _0736_
rlabel metal3 21392 80136 21392 80136 0 _0737_
rlabel metal2 23632 95144 23632 95144 0 _0738_
rlabel metal2 29512 63784 29512 63784 0 _0739_
rlabel metal2 30912 70056 30912 70056 0 _0740_
rlabel metal3 31304 75656 31304 75656 0 _0741_
rlabel metal2 30072 75992 30072 75992 0 _0742_
rlabel metal3 28504 76440 28504 76440 0 _0743_
rlabel metal2 27048 76664 27048 76664 0 _0744_
rlabel metal2 24136 77616 24136 77616 0 _0745_
rlabel metal3 24976 76664 24976 76664 0 _0746_
rlabel metal2 26824 82208 26824 82208 0 _0747_
rlabel metal3 23576 78568 23576 78568 0 _0748_
rlabel metal2 25592 77728 25592 77728 0 _0749_
rlabel metal2 24864 75656 24864 75656 0 _0750_
rlabel metal2 25200 86072 25200 86072 0 _0751_
rlabel metal2 29512 58912 29512 58912 0 _0752_
rlabel metal2 31360 70952 31360 70952 0 _0753_
rlabel metal2 31416 77112 31416 77112 0 _0754_
rlabel metal2 31528 78232 31528 78232 0 _0755_
rlabel metal2 27720 79072 27720 79072 0 _0756_
rlabel metal3 27664 78792 27664 78792 0 _0757_
rlabel metal2 27272 77392 27272 77392 0 _0758_
rlabel metal2 26600 77560 26600 77560 0 _0759_
rlabel metal3 26824 89544 26824 89544 0 _0760_
rlabel metal2 22120 78176 22120 78176 0 _0761_
rlabel metal2 27440 95816 27440 95816 0 _0762_
rlabel metal2 32200 69776 32200 69776 0 _0763_
rlabel metal2 30016 66472 30016 66472 0 _0764_
rlabel metal2 27608 69160 27608 69160 0 _0765_
rlabel metal2 29624 72576 29624 72576 0 _0766_
rlabel metal2 26712 70336 26712 70336 0 _0767_
rlabel metal2 27048 70168 27048 70168 0 _0768_
rlabel metal2 29400 69328 29400 69328 0 _0769_
rlabel metal2 25928 71064 25928 71064 0 _0770_
rlabel metal2 24472 75320 24472 75320 0 _0771_
rlabel metal2 25592 72240 25592 72240 0 _0772_
rlabel metal2 26152 72352 26152 72352 0 _0773_
rlabel metal3 25480 75096 25480 75096 0 _0774_
rlabel metal3 26320 86408 26320 86408 0 _0775_
rlabel metal2 26824 75544 26824 75544 0 _0776_
rlabel metal3 29064 73528 29064 73528 0 _0777_
rlabel metal2 28952 57512 28952 57512 0 _0778_
rlabel metal2 31080 75880 31080 75880 0 _0779_
rlabel metal2 29064 75600 29064 75600 0 _0780_
rlabel metal2 28504 74816 28504 74816 0 _0781_
rlabel metal2 27440 81928 27440 81928 0 _0782_
rlabel metal2 25480 83328 25480 83328 0 _0783_
rlabel metal3 24808 87864 24808 87864 0 _0784_
rlabel metal2 29288 67200 29288 67200 0 _0785_
rlabel metal2 25816 70560 25816 70560 0 _0786_
rlabel metal2 25424 77000 25424 77000 0 _0787_
rlabel metal2 25704 81032 25704 81032 0 _0788_
rlabel metal2 24192 86744 24192 86744 0 _0789_
rlabel metal3 22232 86632 22232 86632 0 _0790_
rlabel metal2 20440 85064 20440 85064 0 _0791_
rlabel metal2 21784 20944 21784 20944 0 _0792_
rlabel metal2 21672 64400 21672 64400 0 _0793_
rlabel metal3 6888 3416 6888 3416 0 _0794_
rlabel metal2 7728 49224 7728 49224 0 _0795_
rlabel metal2 15064 1848 15064 1848 0 _0796_
rlabel metal2 16296 2464 16296 2464 0 _0797_
rlabel metal2 10472 3976 10472 3976 0 _0798_
rlabel metal3 12320 3304 12320 3304 0 _0799_
rlabel metal2 13720 2408 13720 2408 0 _0800_
rlabel metal2 11592 2520 11592 2520 0 _0801_
rlabel metal2 33096 3024 33096 3024 0 _0802_
rlabel metal2 33992 3472 33992 3472 0 _0803_
rlabel metal3 16548 2632 16548 2632 0 _0804_
rlabel metal3 26320 3304 26320 3304 0 _0805_
rlabel metal2 25928 3640 25928 3640 0 _0806_
rlabel metal2 10584 2632 10584 2632 0 _0807_
rlabel metal2 19768 78568 19768 78568 0 _0808_
rlabel metal3 10360 81368 10360 81368 0 _0809_
rlabel metal2 6328 81984 6328 81984 0 _0810_
rlabel metal2 21224 83048 21224 83048 0 _0811_
rlabel metal2 6328 79184 6328 79184 0 _0812_
rlabel metal3 13608 78680 13608 78680 0 _0813_
rlabel metal2 7000 74256 7000 74256 0 _0814_
rlabel metal3 22904 75040 22904 75040 0 _0815_
rlabel metal2 6104 74816 6104 74816 0 _0816_
rlabel metal2 22008 77224 22008 77224 0 _0817_
rlabel metal2 9912 78512 9912 78512 0 _0818_
rlabel metal2 9464 76216 9464 76216 0 _0819_
rlabel metal2 9688 82768 9688 82768 0 _0820_
rlabel metal2 5320 11032 5320 11032 0 _0821_
rlabel metal2 17920 26040 17920 26040 0 _0822_
rlabel metal2 10136 2912 10136 2912 0 _0823_
rlabel metal3 9408 4088 9408 4088 0 _0824_
rlabel metal2 37016 26320 37016 26320 0 _0825_
rlabel metal2 13832 86968 13832 86968 0 _0826_
rlabel metal2 26824 53816 26824 53816 0 _0827_
rlabel metal3 32536 87416 32536 87416 0 _0828_
rlabel metal2 11704 36680 11704 36680 0 _0829_
rlabel metal2 12600 33600 12600 33600 0 _0830_
rlabel metal2 16240 31080 16240 31080 0 _0831_
rlabel metal3 24080 47880 24080 47880 0 _0832_
rlabel metal2 20104 30016 20104 30016 0 _0833_
rlabel metal3 13104 28840 13104 28840 0 _0834_
rlabel metal2 10192 22680 10192 22680 0 _0835_
rlabel metal2 6552 14784 6552 14784 0 _0836_
rlabel metal2 6104 12320 6104 12320 0 _0837_
rlabel metal2 9576 11312 9576 11312 0 _0838_
rlabel metal2 11424 45304 11424 45304 0 _0839_
rlabel metal2 11368 48608 11368 48608 0 _0840_
rlabel metal2 6328 51072 6328 51072 0 _0841_
rlabel metal2 26712 10248 26712 10248 0 cal_lut\[100\]
rlabel metal2 26320 15512 26320 15512 0 cal_lut\[101\]
rlabel metal2 23800 21280 23800 21280 0 cal_lut\[102\]
rlabel metal3 6160 38136 6160 38136 0 cal_lut\[103\]
rlabel metal2 4480 37128 4480 37128 0 cal_lut\[104\]
rlabel metal2 5880 34160 5880 34160 0 cal_lut\[105\]
rlabel metal2 9576 36456 9576 36456 0 cal_lut\[106\]
rlabel metal3 14112 47320 14112 47320 0 cal_lut\[107\]
rlabel metal2 15624 48216 15624 48216 0 cal_lut\[108\]
rlabel metal2 13832 60256 13832 60256 0 cal_lut\[109\]
rlabel metal2 19264 30296 19264 30296 0 cal_lut\[10\]
rlabel metal2 14224 63784 14224 63784 0 cal_lut\[110\]
rlabel metal2 14616 64680 14616 64680 0 cal_lut\[111\]
rlabel metal2 16184 58912 16184 58912 0 cal_lut\[112\]
rlabel metal2 14728 53312 14728 53312 0 cal_lut\[113\]
rlabel metal2 14616 49000 14616 49000 0 cal_lut\[114\]
rlabel metal2 16184 18088 16184 18088 0 cal_lut\[115\]
rlabel metal2 14336 11256 14336 11256 0 cal_lut\[116\]
rlabel metal2 17192 9856 17192 9856 0 cal_lut\[117\]
rlabel metal2 18536 12152 18536 12152 0 cal_lut\[118\]
rlabel metal2 16464 26152 16464 26152 0 cal_lut\[119\]
rlabel metal2 18424 29008 18424 29008 0 cal_lut\[11\]
rlabel metal2 16296 28728 16296 28728 0 cal_lut\[120\]
rlabel metal2 6216 26236 6216 26236 0 cal_lut\[121\]
rlabel metal2 5320 22344 5320 22344 0 cal_lut\[122\]
rlabel metal2 5768 21560 5768 21560 0 cal_lut\[123\]
rlabel metal2 8904 22288 8904 22288 0 cal_lut\[124\]
rlabel metal2 13048 24920 13048 24920 0 cal_lut\[125\]
rlabel metal2 16296 23296 16296 23296 0 cal_lut\[126\]
rlabel metal3 25200 25368 25200 25368 0 cal_lut\[127\]
rlabel metal2 30296 24976 30296 24976 0 cal_lut\[128\]
rlabel metal2 31864 24976 31864 24976 0 cal_lut\[129\]
rlabel metal2 11368 29400 11368 29400 0 cal_lut\[12\]
rlabel metal3 31416 24024 31416 24024 0 cal_lut\[130\]
rlabel metal2 26096 24024 26096 24024 0 cal_lut\[131\]
rlabel metal2 26376 26656 26376 26656 0 cal_lut\[132\]
rlabel metal2 30464 18312 30464 18312 0 cal_lut\[133\]
rlabel metal2 33320 18424 33320 18424 0 cal_lut\[134\]
rlabel metal2 34664 18760 34664 18760 0 cal_lut\[135\]
rlabel metal2 33656 20664 33656 20664 0 cal_lut\[136\]
rlabel metal2 22456 21896 22456 21896 0 cal_lut\[137\]
rlabel metal3 21280 21672 21280 21672 0 cal_lut\[138\]
rlabel metal2 19656 15848 19656 15848 0 cal_lut\[139\]
rlabel metal2 7112 15624 7112 15624 0 cal_lut\[13\]
rlabel metal3 19768 7336 19768 7336 0 cal_lut\[140\]
rlabel metal2 21784 7672 21784 7672 0 cal_lut\[141\]
rlabel metal2 21896 10304 21896 10304 0 cal_lut\[142\]
rlabel metal3 21392 15176 21392 15176 0 cal_lut\[143\]
rlabel metal2 19768 16464 19768 16464 0 cal_lut\[144\]
rlabel metal2 24472 15204 24472 15204 0 cal_lut\[145\]
rlabel metal2 25760 5880 25760 5880 0 cal_lut\[146\]
rlabel metal2 27608 8400 27608 8400 0 cal_lut\[147\]
rlabel metal2 28056 9688 28056 9688 0 cal_lut\[148\]
rlabel metal2 26712 15204 26712 15204 0 cal_lut\[149\]
rlabel metal2 7224 11312 7224 11312 0 cal_lut\[14\]
rlabel metal2 25704 16464 25704 16464 0 cal_lut\[150\]
rlabel metal2 30968 16800 30968 16800 0 cal_lut\[151\]
rlabel metal2 35000 16688 35000 16688 0 cal_lut\[152\]
rlabel metal2 35560 19656 35560 19656 0 cal_lut\[153\]
rlabel metal2 35000 22288 35000 22288 0 cal_lut\[154\]
rlabel metal2 24024 42728 24024 42728 0 cal_lut\[155\]
rlabel metal2 22232 35504 22232 35504 0 cal_lut\[156\]
rlabel metal2 23632 64680 23632 64680 0 cal_lut\[157\]
rlabel metal3 24640 65464 24640 65464 0 cal_lut\[158\]
rlabel metal2 24920 64960 24920 64960 0 cal_lut\[159\]
rlabel metal2 10472 10080 10472 10080 0 cal_lut\[15\]
rlabel metal2 24136 60760 24136 60760 0 cal_lut\[160\]
rlabel metal2 25704 56112 25704 56112 0 cal_lut\[161\]
rlabel metal3 23632 38136 23632 38136 0 cal_lut\[162\]
rlabel metal2 5432 26572 5432 26572 0 cal_lut\[163\]
rlabel metal2 4648 22176 4648 22176 0 cal_lut\[164\]
rlabel metal2 5656 18536 5656 18536 0 cal_lut\[165\]
rlabel metal2 8456 19600 8456 19600 0 cal_lut\[166\]
rlabel metal2 12376 22624 12376 22624 0 cal_lut\[167\]
rlabel metal2 15512 21672 15512 21672 0 cal_lut\[168\]
rlabel metal2 11480 15736 11480 15736 0 cal_lut\[169\]
rlabel metal2 13328 23352 13328 23352 0 cal_lut\[16\]
rlabel metal2 10696 11928 10696 11928 0 cal_lut\[170\]
rlabel metal2 10976 6776 10976 6776 0 cal_lut\[171\]
rlabel metal2 12376 9016 12376 9016 0 cal_lut\[172\]
rlabel metal2 14168 16072 14168 16072 0 cal_lut\[173\]
rlabel metal2 15624 19208 15624 19208 0 cal_lut\[174\]
rlabel metal2 16072 15456 16072 15456 0 cal_lut\[175\]
rlabel metal2 15848 6720 15848 6720 0 cal_lut\[176\]
rlabel metal2 17864 8176 17864 8176 0 cal_lut\[177\]
rlabel metal3 18704 16520 18704 16520 0 cal_lut\[178\]
rlabel metal2 19656 23632 19656 23632 0 cal_lut\[179\]
rlabel metal2 12936 48160 12936 48160 0 cal_lut\[17\]
rlabel metal2 16408 22400 16408 22400 0 cal_lut\[180\]
rlabel metal3 4928 39368 4928 39368 0 cal_lut\[181\]
rlabel metal2 4872 39004 4872 39004 0 cal_lut\[182\]
rlabel metal3 6104 41832 6104 41832 0 cal_lut\[183\]
rlabel metal2 9016 44184 9016 44184 0 cal_lut\[184\]
rlabel metal2 8008 49168 8008 49168 0 cal_lut\[185\]
rlabel metal3 7112 48104 7112 48104 0 cal_lut\[186\]
rlabel metal2 5824 40488 5824 40488 0 cal_lut\[187\]
rlabel metal2 4648 38668 4648 38668 0 cal_lut\[188\]
rlabel metal3 6608 32424 6608 32424 0 cal_lut\[189\]
rlabel metal2 8344 48888 8344 48888 0 cal_lut\[18\]
rlabel metal2 10080 31864 10080 31864 0 cal_lut\[190\]
rlabel metal2 17976 26572 17976 26572 0 cal_lut\[191\]
rlabel metal2 19880 27608 19880 27608 0 cal_lut\[192\]
rlabel metal2 4984 52976 4984 52976 0 cal_lut\[19\]
rlabel metal3 36176 27272 36176 27272 0 cal_lut\[1\]
rlabel metal2 4368 58408 4368 58408 0 cal_lut\[20\]
rlabel metal2 4536 64792 4536 64792 0 cal_lut\[21\]
rlabel metal2 5768 64008 5768 64008 0 cal_lut\[22\]
rlabel via2 8680 59976 8680 59976 0 cal_lut\[23\]
rlabel metal2 11536 46872 11536 46872 0 cal_lut\[24\]
rlabel metal3 15652 63000 15652 63000 0 cal_lut\[25\]
rlabel metal2 15512 69832 15512 69832 0 cal_lut\[26\]
rlabel metal2 14840 63392 14840 63392 0 cal_lut\[27\]
rlabel metal2 17640 58016 17640 58016 0 cal_lut\[28\]
rlabel metal2 21896 53312 21896 53312 0 cal_lut\[29\]
rlabel metal2 28616 32088 28616 32088 0 cal_lut\[2\]
rlabel metal2 24136 43624 24136 43624 0 cal_lut\[30\]
rlabel metal2 26936 29064 26936 29064 0 cal_lut\[31\]
rlabel metal2 31024 28728 31024 28728 0 cal_lut\[32\]
rlabel metal3 32200 30184 32200 30184 0 cal_lut\[33\]
rlabel metal3 28840 39256 28840 39256 0 cal_lut\[34\]
rlabel metal3 26040 43400 26040 43400 0 cal_lut\[35\]
rlabel metal2 26768 49672 26768 49672 0 cal_lut\[36\]
rlabel metal2 26488 64176 26488 64176 0 cal_lut\[37\]
rlabel metal2 17976 69496 17976 69496 0 cal_lut\[38\]
rlabel metal2 19768 68208 19768 68208 0 cal_lut\[39\]
rlabel metal2 29736 32984 29736 32984 0 cal_lut\[3\]
rlabel metal2 20664 63224 20664 63224 0 cal_lut\[40\]
rlabel metal2 20552 55272 20552 55272 0 cal_lut\[41\]
rlabel metal2 16072 52472 16072 52472 0 cal_lut\[42\]
rlabel metal2 4648 53088 4648 53088 0 cal_lut\[43\]
rlabel metal2 4704 58408 4704 58408 0 cal_lut\[44\]
rlabel metal2 4648 62188 4648 62188 0 cal_lut\[45\]
rlabel metal3 7000 58408 7000 58408 0 cal_lut\[46\]
rlabel metal3 8848 53592 8848 53592 0 cal_lut\[47\]
rlabel metal2 9016 54432 9016 54432 0 cal_lut\[48\]
rlabel metal2 4648 49616 4648 49616 0 cal_lut\[49\]
rlabel metal2 30184 39088 30184 39088 0 cal_lut\[4\]
rlabel metal2 4200 41944 4200 41944 0 cal_lut\[50\]
rlabel metal2 5544 42840 5544 42840 0 cal_lut\[51\]
rlabel metal2 9800 42336 9800 42336 0 cal_lut\[52\]
rlabel metal2 15176 40880 15176 40880 0 cal_lut\[53\]
rlabel metal2 21672 37632 21672 37632 0 cal_lut\[54\]
rlabel metal3 29624 35896 29624 35896 0 cal_lut\[55\]
rlabel metal2 35672 31920 35672 31920 0 cal_lut\[56\]
rlabel metal2 37016 36120 37016 36120 0 cal_lut\[57\]
rlabel metal2 35896 40320 35896 40320 0 cal_lut\[58\]
rlabel metal2 29960 42112 29960 42112 0 cal_lut\[59\]
rlabel metal2 32088 54096 32088 54096 0 cal_lut\[5\]
rlabel metal3 30744 44184 30744 44184 0 cal_lut\[60\]
rlabel metal2 30632 36232 30632 36232 0 cal_lut\[61\]
rlabel metal2 34328 33768 34328 33768 0 cal_lut\[62\]
rlabel metal2 37016 35448 37016 35448 0 cal_lut\[63\]
rlabel metal2 36232 39872 36232 39872 0 cal_lut\[64\]
rlabel metal2 33096 43120 33096 43120 0 cal_lut\[65\]
rlabel metal2 30352 44968 30352 44968 0 cal_lut\[66\]
rlabel metal3 30968 48104 30968 48104 0 cal_lut\[67\]
rlabel metal3 36176 47544 36176 47544 0 cal_lut\[68\]
rlabel metal2 35336 46480 35336 46480 0 cal_lut\[69\]
rlabel metal2 29400 54936 29400 54936 0 cal_lut\[6\]
rlabel metal2 35224 49000 35224 49000 0 cal_lut\[70\]
rlabel metal2 23688 47712 23688 47712 0 cal_lut\[71\]
rlabel metal3 20496 49112 20496 49112 0 cal_lut\[72\]
rlabel metal2 30072 49336 30072 49336 0 cal_lut\[73\]
rlabel metal2 33600 50120 33600 50120 0 cal_lut\[74\]
rlabel metal2 35784 48104 35784 48104 0 cal_lut\[75\]
rlabel metal2 37576 52080 37576 52080 0 cal_lut\[76\]
rlabel metal2 22344 52920 22344 52920 0 cal_lut\[77\]
rlabel metal2 12936 53200 12936 53200 0 cal_lut\[78\]
rlabel metal3 8848 63336 8848 63336 0 cal_lut\[79\]
rlabel metal2 25424 48216 25424 48216 0 cal_lut\[7\]
rlabel metal2 8680 66416 8680 66416 0 cal_lut\[80\]
rlabel metal3 10528 68488 10528 68488 0 cal_lut\[81\]
rlabel via2 6216 68824 6216 68824 0 cal_lut\[82\]
rlabel metal2 8344 69664 8344 69664 0 cal_lut\[83\]
rlabel metal2 10136 69384 10136 69384 0 cal_lut\[84\]
rlabel metal2 14448 71064 14448 71064 0 cal_lut\[85\]
rlabel metal2 18088 71064 18088 71064 0 cal_lut\[86\]
rlabel metal2 21224 69384 21224 69384 0 cal_lut\[87\]
rlabel metal2 21896 65296 21896 65296 0 cal_lut\[88\]
rlabel metal2 21560 41216 21560 41216 0 cal_lut\[89\]
rlabel metal2 13160 34552 13160 34552 0 cal_lut\[8\]
rlabel metal2 19544 39088 19544 39088 0 cal_lut\[90\]
rlabel metal3 15484 38024 15484 38024 0 cal_lut\[91\]
rlabel metal2 15400 35224 15400 35224 0 cal_lut\[92\]
rlabel metal2 17416 33488 17416 33488 0 cal_lut\[93\]
rlabel metal2 20776 33488 20776 33488 0 cal_lut\[94\]
rlabel metal2 21336 31808 21336 31808 0 cal_lut\[95\]
rlabel metal2 24136 20048 24136 20048 0 cal_lut\[96\]
rlabel metal2 24024 16632 24024 16632 0 cal_lut\[97\]
rlabel metal2 26040 9744 26040 9744 0 cal_lut\[98\]
rlabel metal2 26600 8456 26600 8456 0 cal_lut\[99\]
rlabel metal2 15624 32312 15624 32312 0 cal_lut\[9\]
rlabel metal2 4760 1246 4760 1246 0 clk
rlabel metal2 23576 80304 23576 80304 0 clknet_0__0385_
rlabel metal2 20664 76888 20664 76888 0 clknet_0__0387_
rlabel metal2 25480 78736 25480 78736 0 clknet_0__0737_
rlabel metal2 26152 76608 26152 76608 0 clknet_0__0750_
rlabel metal2 25032 66584 25032 66584 0 clknet_0_clk
rlabel metal2 25704 86548 25704 86548 0 clknet_0_net66
rlabel metal2 30240 88872 30240 88872 0 clknet_0_temp1.i_precharge_n
rlabel metal2 18872 81592 18872 81592 0 clknet_1_0__leaf__0385_
rlabel metal2 16856 76888 16856 76888 0 clknet_1_0__leaf__0387_
rlabel metal2 20776 77952 20776 77952 0 clknet_1_0__leaf__0737_
rlabel metal2 23072 78568 23072 78568 0 clknet_1_0__leaf__0750_
rlabel metal2 23464 83160 23464 83160 0 clknet_1_0__leaf_net66
rlabel metal2 27496 87472 27496 87472 0 clknet_1_0__leaf_temp1.i_precharge_n
rlabel metal2 19096 84896 19096 84896 0 clknet_1_1__leaf__0385_
rlabel metal3 18928 74088 18928 74088 0 clknet_1_1__leaf__0387_
rlabel metal3 21728 80584 21728 80584 0 clknet_1_1__leaf__0737_
rlabel metal2 25032 79184 25032 79184 0 clknet_1_1__leaf__0750_
rlabel metal2 25368 86744 25368 86744 0 clknet_1_1__leaf_net66
rlabel metal2 23688 88984 23688 88984 0 clknet_1_1__leaf_temp1.i_precharge_n
rlabel metal2 11144 67536 11144 67536 0 clknet_2_0__leaf_clk
rlabel metal2 16072 88200 16072 88200 0 clknet_2_1__leaf_clk
rlabel metal3 19712 71736 19712 71736 0 clknet_2_2__leaf_clk
rlabel metal2 31080 88536 31080 88536 0 clknet_2_3__leaf_clk
rlabel metal2 20440 88928 20440 88928 0 ctr\[0\]
rlabel metal2 32928 86744 32928 86744 0 ctr\[10\]
rlabel metal2 34944 85848 34944 85848 0 ctr\[11\]
rlabel metal2 31920 82488 31920 82488 0 ctr\[12\]
rlabel metal2 19992 83552 19992 83552 0 ctr\[1\]
rlabel metal2 15848 78344 15848 78344 0 ctr\[2\]
rlabel metal2 22344 84168 22344 84168 0 ctr\[3\]
rlabel metal2 13776 85736 13776 85736 0 ctr\[4\]
rlabel metal2 16240 88872 16240 88872 0 ctr\[5\]
rlabel metal2 19208 87752 19208 87752 0 ctr\[6\]
rlabel metal2 27048 88872 27048 88872 0 ctr\[7\]
rlabel metal2 31640 86128 31640 86128 0 ctr\[8\]
rlabel metal2 31864 85792 31864 85792 0 ctr\[9\]
rlabel metal2 19096 79240 19096 79240 0 dbg3\[0\]
rlabel metal2 16184 77336 16184 77336 0 dbg3\[1\]
rlabel metal2 14392 75208 14392 75208 0 dbg3\[2\]
rlabel metal2 18872 71960 18872 71960 0 dbg3\[3\]
rlabel metal2 22064 69384 22064 69384 0 dbg3\[4\]
rlabel metal3 23800 71624 23800 71624 0 dbg3\[5\]
rlabel metal2 33264 68824 33264 68824 0 dec1._000_
rlabel metal2 33432 71176 33432 71176 0 dec1._001_
rlabel metal2 37352 70112 37352 70112 0 dec1._002_
rlabel metal2 33152 67704 33152 67704 0 dec1._003_
rlabel metal2 33320 61040 33320 61040 0 dec1._004_
rlabel metal3 32480 60200 32480 60200 0 dec1._005_
rlabel metal3 35784 60648 35784 60648 0 dec1._006_
rlabel metal3 34664 61768 34664 61768 0 dec1._007_
rlabel metal2 36232 58744 36232 58744 0 dec1._008_
rlabel metal2 32536 58856 32536 58856 0 dec1._009_
rlabel metal2 34888 59248 34888 59248 0 dec1._010_
rlabel metal2 33040 62440 33040 62440 0 dec1._011_
rlabel metal2 36344 59416 36344 59416 0 dec1._012_
rlabel metal2 37240 61376 37240 61376 0 dec1._013_
rlabel metal2 35896 59808 35896 59808 0 dec1._014_
rlabel metal2 32536 62272 32536 62272 0 dec1._015_
rlabel metal2 33880 64568 33880 64568 0 dec1._016_
rlabel metal2 35056 64568 35056 64568 0 dec1._017_
rlabel metal2 37576 65912 37576 65912 0 dec1._018_
rlabel metal2 37352 65800 37352 65800 0 dec1._019_
rlabel metal2 32704 60872 32704 60872 0 dec1._020_
rlabel metal2 33432 64008 33432 64008 0 dec1._021_
rlabel metal2 34104 63420 34104 63420 0 dec1._022_
rlabel metal2 33656 63560 33656 63560 0 dec1._023_
rlabel metal2 37576 60592 37576 60592 0 dec1._024_
rlabel metal2 33544 64456 33544 64456 0 dec1._025_
rlabel metal2 34552 65520 34552 65520 0 dec1._026_
rlabel metal2 35896 64288 35896 64288 0 dec1._027_
rlabel metal2 38248 62776 38248 62776 0 dec1._028_
rlabel metal2 35616 56952 35616 56952 0 dec1._029_
rlabel metal2 37128 64456 37128 64456 0 dec1._030_
rlabel metal3 36680 64792 36680 64792 0 dec1._031_
rlabel metal2 35504 66136 35504 66136 0 dec1._032_
rlabel metal2 35896 65744 35896 65744 0 dec1._033_
rlabel metal2 36120 64064 36120 64064 0 dec1._034_
rlabel metal2 32088 64288 32088 64288 0 dec1._035_
rlabel metal2 35224 63168 35224 63168 0 dec1._036_
rlabel metal2 35616 63112 35616 63112 0 dec1._037_
rlabel metal2 36008 64288 36008 64288 0 dec1._038_
rlabel metal2 37464 65968 37464 65968 0 dec1._039_
rlabel metal2 35560 68320 35560 68320 0 dec1._040_
rlabel metal2 34888 70840 34888 70840 0 dec1._041_
rlabel metal2 31640 67088 31640 67088 0 dec1._042_
rlabel metal2 33656 68152 33656 68152 0 dec1._043_
rlabel metal2 33040 68040 33040 68040 0 dec1._044_
rlabel metal2 33880 68040 33880 68040 0 dec1._045_
rlabel metal2 34776 68656 34776 68656 0 dec1._046_
rlabel metal2 33432 67200 33432 67200 0 dec1._047_
rlabel metal3 33824 65464 33824 65464 0 dec1._048_
rlabel metal2 37912 64960 37912 64960 0 dec1._049_
rlabel metal2 33824 65576 33824 65576 0 dec1._050_
rlabel metal2 33432 68712 33432 68712 0 dec1._051_
rlabel metal3 35504 69384 35504 69384 0 dec1._052_
rlabel metal3 34552 67816 34552 67816 0 dec1._053_
rlabel metal2 37576 68824 37576 68824 0 dec1._054_
rlabel metal3 36456 67592 36456 67592 0 dec1._055_
rlabel metal2 33768 70112 33768 70112 0 dec1._056_
rlabel metal2 35000 65520 35000 65520 0 dec1._057_
rlabel metal2 36904 68824 36904 68824 0 dec1._058_
rlabel metal2 33320 70840 33320 70840 0 dec1._059_
rlabel metal3 33712 68712 33712 68712 0 dec1.i_bin\[0\]
rlabel metal2 33656 66304 33656 66304 0 dec1.i_bin\[1\]
rlabel metal3 33320 62104 33320 62104 0 dec1.i_bin\[2\]
rlabel metal2 33096 60592 33096 60592 0 dec1.i_bin\[3\]
rlabel metal3 33488 61544 33488 61544 0 dec1.i_bin\[4\]
rlabel metal3 31696 61544 31696 61544 0 dec1.i_bin\[5\]
rlabel metal2 32872 59640 32872 59640 0 dec1.i_bin\[6\]
rlabel metal2 29512 69216 29512 69216 0 dec1.i_ones
rlabel metal2 34832 69384 34832 69384 0 dec1.i_tens
rlabel metal2 35840 69944 35840 69944 0 dec1.o_dec\[0\]
rlabel metal2 35672 70028 35672 70028 0 dec1.o_dec\[1\]
rlabel metal2 35056 72408 35056 72408 0 dec1.o_dec\[2\]
rlabel metal2 33656 70784 33656 70784 0 dec1.o_dec\[3\]
rlabel metal2 36904 1848 36904 1848 0 i_wb_addr[0]
rlabel metal2 27608 1680 27608 1680 0 i_wb_addr[10]
rlabel metal2 26600 1680 26600 1680 0 i_wb_addr[11]
rlabel metal2 26096 1960 26096 1960 0 i_wb_addr[12]
rlabel metal2 25200 1848 25200 1848 0 i_wb_addr[13]
rlabel metal2 24584 1680 24584 1680 0 i_wb_addr[14]
rlabel metal2 22904 2632 22904 2632 0 i_wb_addr[15]
rlabel metal3 22848 1960 22848 1960 0 i_wb_addr[16]
rlabel metal2 21112 2632 21112 2632 0 i_wb_addr[17]
rlabel metal2 19880 1792 19880 1792 0 i_wb_addr[18]
rlabel metal2 19152 1848 19152 1848 0 i_wb_addr[19]
rlabel metal2 36232 1904 36232 1904 0 i_wb_addr[1]
rlabel metal2 18312 1848 18312 1848 0 i_wb_addr[20]
rlabel metal2 17696 1960 17696 1960 0 i_wb_addr[21]
rlabel metal3 17024 2744 17024 2744 0 i_wb_addr[22]
rlabel metal2 15512 2254 15512 2254 0 i_wb_addr[23]
rlabel metal2 14616 1834 14616 1834 0 i_wb_addr[24]
rlabel metal2 13776 1624 13776 1624 0 i_wb_addr[25]
rlabel metal2 12376 1736 12376 1736 0 i_wb_addr[26]
rlabel metal2 11704 2632 11704 2632 0 i_wb_addr[27]
rlabel metal2 11256 2632 11256 2632 0 i_wb_addr[28]
rlabel metal2 10472 2296 10472 2296 0 i_wb_addr[29]
rlabel metal2 34888 2296 34888 2296 0 i_wb_addr[2]
rlabel metal2 9352 1848 9352 1848 0 i_wb_addr[30]
rlabel metal2 8344 1078 8344 1078 0 i_wb_addr[31]
rlabel metal3 34552 1960 34552 1960 0 i_wb_addr[3]
rlabel metal2 32872 1680 32872 1680 0 i_wb_addr[4]
rlabel metal2 31640 1022 31640 1022 0 i_wb_addr[5]
rlabel metal2 30856 1848 30856 1848 0 i_wb_addr[6]
rlabel metal2 29960 1848 29960 1848 0 i_wb_addr[7]
rlabel metal2 29400 1736 29400 1736 0 i_wb_addr[8]
rlabel metal2 28224 1848 28224 1848 0 i_wb_addr[9]
rlabel metal2 7560 1848 7560 1848 0 i_wb_cyc
rlabel metal3 5936 1736 5936 1736 0 i_wb_stb
rlabel metal3 4872 1848 4872 1848 0 i_wb_we
rlabel metal2 38360 8456 38360 8456 0 io_in[0]
rlabel metal2 38248 25256 38248 25256 0 io_in[1]
rlabel metal2 38248 41440 38248 41440 0 io_in[2]
rlabel metal2 38248 58016 38248 58016 0 io_in[3]
rlabel metal3 38962 74872 38962 74872 0 io_in[4]
rlabel metal2 38248 91784 38248 91784 0 io_in[5]
rlabel metal3 15120 81312 15120 81312 0 io_out[0]
rlabel metal2 35896 97930 35896 97930 0 io_out[1]
rlabel metal2 33432 97818 33432 97818 0 io_out[2]
rlabel metal2 30968 97706 30968 97706 0 io_out[3]
rlabel metal2 28504 98546 28504 98546 0 io_out[4]
rlabel metal2 26040 98574 26040 98574 0 io_out[5]
rlabel metal3 24360 95480 24360 95480 0 io_out[6]
rlabel metal2 21112 98574 21112 98574 0 io_out[7]
rlabel metal2 36680 2464 36680 2464 0 net1
rlabel metal2 20216 2352 20216 2352 0 net10
rlabel metal2 19768 2296 19768 2296 0 net11
rlabel metal2 36008 2408 36008 2408 0 net12
rlabel metal2 18760 2240 18760 2240 0 net13
rlabel metal3 18256 3416 18256 3416 0 net14
rlabel metal2 17304 2968 17304 2968 0 net15
rlabel metal2 15736 3472 15736 3472 0 net16
rlabel metal2 14896 2744 14896 2744 0 net17
rlabel metal3 14784 2856 14784 2856 0 net18
rlabel metal2 12600 2072 12600 2072 0 net19
rlabel metal2 27384 1960 27384 1960 0 net2
rlabel metal2 11928 2296 11928 2296 0 net20
rlabel metal2 10808 1848 10808 1848 0 net21
rlabel metal2 10248 2464 10248 2464 0 net22
rlabel metal2 34552 3024 34552 3024 0 net23
rlabel metal2 9856 1848 9856 1848 0 net24
rlabel metal3 9576 3528 9576 3528 0 net25
rlabel metal2 34216 1736 34216 1736 0 net26
rlabel metal2 33264 1848 33264 1848 0 net27
rlabel metal3 33096 3416 33096 3416 0 net28
rlabel metal2 31248 1848 31248 1848 0 net29
rlabel metal2 27104 1736 27104 1736 0 net3
rlabel metal2 30856 2856 30856 2856 0 net30
rlabel metal3 28560 1736 28560 1736 0 net31
rlabel metal2 28616 1848 28616 1848 0 net32
rlabel metal2 8008 2604 8008 2604 0 net33
rlabel metal2 7112 2520 7112 2520 0 net34
rlabel metal2 6216 2632 6216 2632 0 net35
rlabel metal2 18312 20944 18312 20944 0 net36
rlabel metal2 37912 25480 37912 25480 0 net37
rlabel metal3 34832 41384 34832 41384 0 net38
rlabel metal2 38304 70840 38304 70840 0 net39
rlabel metal2 26320 1848 26320 1848 0 net4
rlabel metal2 26824 71680 26824 71680 0 net40
rlabel metal2 37912 90608 37912 90608 0 net41
rlabel metal2 4368 1848 4368 1848 0 net42
rlabel metal2 2632 19152 2632 19152 0 net43
rlabel metal2 1848 22736 1848 22736 0 net44
rlabel metal2 16800 23352 16800 23352 0 net45
rlabel metal2 26712 17192 26712 17192 0 net46
rlabel metal2 23968 23016 23968 23016 0 net47
rlabel metal2 29736 24304 29736 24304 0 net48
rlabel metal2 1848 38752 1848 38752 0 net49
rlabel metal2 25592 2352 25592 2352 0 net5
rlabel metal2 1848 58408 1848 58408 0 net50
rlabel metal2 15624 40096 15624 40096 0 net51
rlabel via1 22344 38802 22344 38802 0 net52
rlabel metal3 20664 70168 20664 70168 0 net53
rlabel metal2 18760 97496 18760 97496 0 net54
rlabel metal3 16576 97384 16576 97384 0 net55
rlabel metal2 13720 98546 13720 98546 0 net56
rlabel metal2 11480 97440 11480 97440 0 net57
rlabel metal2 9352 98560 9352 98560 0 net58
rlabel metal2 6552 97440 6552 97440 0 net59
rlabel metal2 24920 2072 24920 2072 0 net6
rlabel metal2 4088 97440 4088 97440 0 net60
rlabel metal2 1680 97384 1680 97384 0 net61
rlabel metal3 1022 94360 1022 94360 0 net62
rlabel metal2 14168 93240 14168 93240 0 net63
rlabel metal2 10360 93240 10360 93240 0 net64
rlabel metal2 14616 93184 14616 93184 0 net65
rlabel metal3 21728 86856 21728 86856 0 net66
rlabel metal3 21672 84392 21672 84392 0 net67
rlabel metal3 23016 85848 23016 85848 0 net68
rlabel metal2 20272 15848 20272 15848 0 net69
rlabel metal2 23240 2296 23240 2296 0 net7
rlabel metal2 10416 18312 10416 18312 0 net70
rlabel metal2 22288 1848 22288 1848 0 net8
rlabel metal2 21448 2352 21448 2352 0 net9
rlabel metal3 406 5656 406 5656 0 o_wb_ack
rlabel metal2 8120 16744 8120 16744 0 o_wb_data[0]
rlabel metal3 1134 25368 1134 25368 0 o_wb_data[1]
rlabel metal2 3304 51464 3304 51464 0 o_wb_data[2]
rlabel metal3 1918 45080 1918 45080 0 o_wb_data[3]
rlabel metal2 3696 65352 3696 65352 0 o_wb_data[4]
rlabel metal2 6776 66864 6776 66864 0 o_wb_data[5]
rlabel metal3 6272 75768 6272 75768 0 o_wb_data[6]
rlabel metal3 5544 82600 5544 82600 0 o_wb_data[7]
rlabel metal2 4088 1512 4088 1512 0 reset
rlabel metal2 35112 73192 35112 73192 0 seg1._00_
rlabel metal3 36568 78008 36568 78008 0 seg1._01_
rlabel metal2 35448 77168 35448 77168 0 seg1._02_
rlabel metal2 34440 77168 34440 77168 0 seg1._03_
rlabel metal2 35168 77448 35168 77448 0 seg1._04_
rlabel metal2 38024 77952 38024 77952 0 seg1._05_
rlabel metal2 36792 76552 36792 76552 0 seg1._06_
rlabel metal2 36008 78008 36008 78008 0 seg1._07_
rlabel metal3 34664 76440 34664 76440 0 seg1._08_
rlabel metal2 35280 75096 35280 75096 0 seg1._09_
rlabel metal2 33712 75096 33712 75096 0 seg1._10_
rlabel metal3 35952 77896 35952 77896 0 seg1._11_
rlabel metal3 36904 75096 36904 75096 0 seg1._12_
rlabel metal3 34272 75544 34272 75544 0 seg1._13_
rlabel metal3 36064 75880 36064 75880 0 seg1._14_
rlabel metal2 37688 76776 37688 76776 0 seg1._15_
rlabel metal2 34552 75712 34552 75712 0 seg1._16_
rlabel metal3 35056 76216 35056 76216 0 seg1._17_
rlabel metal2 33432 75600 33432 75600 0 seg1._18_
rlabel metal3 34720 75768 34720 75768 0 seg1._19_
rlabel metal2 32704 76552 32704 76552 0 seg1._20_
rlabel metal2 35000 78456 35000 78456 0 seg1._21_
rlabel metal2 34776 75264 34776 75264 0 seg1._22_
rlabel metal2 34048 74088 34048 74088 0 seg1._23_
rlabel metal2 37016 76888 37016 76888 0 seg1._24_
rlabel metal2 34776 77336 34776 77336 0 seg1._25_
rlabel metal2 31752 78512 31752 78512 0 seg1.o_segments\[0\]
rlabel metal3 32424 77112 32424 77112 0 seg1.o_segments\[1\]
rlabel metal2 33432 76776 33432 76776 0 seg1.o_segments\[2\]
rlabel metal2 33096 75152 33096 75152 0 seg1.o_segments\[3\]
rlabel metal2 31584 76552 31584 76552 0 seg1.o_segments\[4\]
rlabel metal2 32200 71120 32200 71120 0 seg1.o_segments\[5\]
rlabel metal2 31304 76328 31304 76328 0 seg1.o_segments\[6\]
rlabel metal3 12824 91336 12824 91336 0 temp1.dac._0_
rlabel metal2 13832 91448 13832 91448 0 temp1.dac._1_
rlabel metal2 25592 92624 25592 92624 0 temp1.dac.i_data\[0\]
rlabel metal3 22512 92008 22512 92008 0 temp1.dac.i_data\[1\]
rlabel metal2 22568 89768 22568 89768 0 temp1.dac.i_data\[2\]
rlabel metal2 27160 86912 27160 86912 0 temp1.dac.i_data\[3\]
rlabel metal3 27132 92120 27132 92120 0 temp1.dac.i_data\[4\]
rlabel metal2 28392 91364 28392 91364 0 temp1.dac.i_data\[5\]
rlabel metal2 10136 92232 10136 92232 0 temp1.dac.i_enable
rlabel metal2 25536 94472 25536 94472 0 temp1.dac.parallel_cells\[0\].vdac_batch._0_
rlabel metal2 24584 94024 24584 94024 0 temp1.dac.parallel_cells\[0\].vdac_batch._1_
rlabel metal2 24192 93128 24192 93128 0 temp1.dac.parallel_cells\[0\].vdac_batch._2_
rlabel metal2 24696 93968 24696 93968 0 temp1.dac.parallel_cells\[0\].vdac_batch.en_pupd
rlabel metal2 25368 94976 25368 94976 0 temp1.dac.parallel_cells\[0\].vdac_batch.en_vref
rlabel metal2 25704 93408 25704 93408 0 temp1.dac.parallel_cells\[0\].vdac_batch.npu_pd
rlabel metal2 7672 96432 7672 96432 0 temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
rlabel metal2 22512 94472 22512 94472 0 temp1.dac.parallel_cells\[1\].vdac_batch._0_
rlabel metal2 20328 94024 20328 94024 0 temp1.dac.parallel_cells\[1\].vdac_batch._1_
rlabel metal3 21112 93912 21112 93912 0 temp1.dac.parallel_cells\[1\].vdac_batch._2_
rlabel metal2 21336 93576 21336 93576 0 temp1.dac.parallel_cells\[1\].vdac_batch.en_pupd
rlabel metal2 22232 95536 22232 95536 0 temp1.dac.parallel_cells\[1\].vdac_batch.en_vref
rlabel metal2 22344 92624 22344 92624 0 temp1.dac.parallel_cells\[1\].vdac_batch.npu_pd
rlabel metal2 16464 94472 16464 94472 0 temp1.dac.parallel_cells\[2\].vdac_batch._0_
rlabel metal3 16296 93688 16296 93688 0 temp1.dac.parallel_cells\[2\].vdac_batch._1_
rlabel metal2 16296 93968 16296 93968 0 temp1.dac.parallel_cells\[2\].vdac_batch._2_
rlabel metal2 17528 94080 17528 94080 0 temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd
rlabel metal2 14728 94976 14728 94976 0 temp1.dac.parallel_cells\[2\].vdac_batch.en_vref
rlabel metal2 19320 93800 19320 93800 0 temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd
rlabel metal2 11704 86352 11704 86352 0 temp1.dac.parallel_cells\[3\].vdac_batch._0_
rlabel metal2 12600 87696 12600 87696 0 temp1.dac.parallel_cells\[3\].vdac_batch._1_
rlabel metal2 10696 87304 10696 87304 0 temp1.dac.parallel_cells\[3\].vdac_batch._2_
rlabel metal2 7112 87808 7112 87808 0 temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd
rlabel metal2 4312 86576 4312 86576 0 temp1.dac.parallel_cells\[3\].vdac_batch.en_vref
rlabel metal2 7560 89376 7560 89376 0 temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd
rlabel metal2 10584 91896 10584 91896 0 temp1.dac.parallel_cells\[4\].vdac_batch._0_
rlabel metal2 25704 91336 25704 91336 0 temp1.dac.parallel_cells\[4\].vdac_batch._1_
rlabel metal2 26152 90664 26152 90664 0 temp1.dac.parallel_cells\[4\].vdac_batch._2_
rlabel metal2 31864 92848 31864 92848 0 temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd
rlabel metal2 6776 95648 6776 95648 0 temp1.dac.parallel_cells\[4\].vdac_batch.en_vref
rlabel metal3 30744 96040 30744 96040 0 temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd
rlabel metal2 12376 90608 12376 90608 0 temp1.dac.vdac_single._0_
rlabel metal2 12264 91952 12264 91952 0 temp1.dac.vdac_single._1_
rlabel metal2 12600 92176 12600 92176 0 temp1.dac.vdac_single._2_
rlabel metal2 13496 92848 13496 92848 0 temp1.dac.vdac_single.en_pupd
rlabel metal2 12656 90776 12656 90776 0 temp1.dac.vdac_single.en_vref
rlabel metal2 12152 93352 12152 93352 0 temp1.dac.vdac_single.npu_pd
rlabel metal2 20664 88312 20664 88312 0 temp1.dcdel_capnode_notouch_
rlabel metal2 24696 89544 24696 89544 0 temp1.i_precharge_n
rlabel metal3 19488 81032 19488 81032 0 temp_delay_last
<< properties >>
string FIXED_BBOX 0 0 40000 100000
<< end >>
