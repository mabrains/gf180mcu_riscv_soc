module core_alu (clk,
    i_wb_cyc,
    i_wb_stb,
    i_wb_we,
    o_wb_ack,
    o_wb_stall,
    reset,
    vdd,
    vss,
    i_wb_addr,
    i_wb_data,
    o_wb_data);
 input clk;
 input i_wb_cyc;
 input i_wb_stb;
 input i_wb_we;
 output o_wb_ack;
 output o_wb_stall;
 input reset;
 input vdd;
 input vss;
 input [31:0] i_wb_addr;
 input [25:0] i_wb_data;
 output [7:0] o_wb_data;

 wire net63;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire \add_out_d0[0] ;
 wire \add_out_d0[1] ;
 wire \add_out_d0[2] ;
 wire \add_out_d0[3] ;
 wire \add_out_d0[4] ;
 wire \add_out_d0[5] ;
 wire \add_out_d0[6] ;
 wire \add_out_d0[7] ;
 wire \add_out_d1[0] ;
 wire \add_out_d1[1] ;
 wire \add_out_d1[2] ;
 wire \add_out_d1[3] ;
 wire \add_out_d1[4] ;
 wire \add_out_d1[5] ;
 wire \add_out_d1[6] ;
 wire \add_out_d1[7] ;
 wire \add_out_d2[0] ;
 wire \add_out_d2[1] ;
 wire \add_out_d2[2] ;
 wire \add_out_d2[3] ;
 wire \add_out_d2[4] ;
 wire \add_out_d2[5] ;
 wire \add_out_d2[6] ;
 wire \add_out_d2[7] ;
 wire \add_out_d3[0] ;
 wire \add_out_d3[1] ;
 wire \add_out_d3[2] ;
 wire \add_out_d3[3] ;
 wire \add_out_d3[4] ;
 wire \add_out_d3[5] ;
 wire \add_out_d3[6] ;
 wire \add_out_d3[7] ;
 wire \add_out_d4[0] ;
 wire \add_out_d4[1] ;
 wire \add_out_d4[2] ;
 wire \add_out_d4[3] ;
 wire \add_out_d4[4] ;
 wire \add_out_d4[5] ;
 wire \add_out_d4[6] ;
 wire \add_out_d4[7] ;
 wire \add_out_d5[0] ;
 wire \add_out_d5[1] ;
 wire \add_out_d5[2] ;
 wire \add_out_d5[3] ;
 wire \add_out_d5[4] ;
 wire \add_out_d5[5] ;
 wire \add_out_d5[6] ;
 wire \add_out_d5[7] ;
 wire \add_out_d6[0] ;
 wire \add_out_d6[1] ;
 wire \add_out_d6[2] ;
 wire \add_out_d6[3] ;
 wire \add_out_d6[4] ;
 wire \add_out_d6[5] ;
 wire \add_out_d6[6] ;
 wire \add_out_d6[7] ;
 wire \add_out_d7[0] ;
 wire \add_out_d7[1] ;
 wire \add_out_d7[2] ;
 wire \add_out_d7[3] ;
 wire \add_out_d7[4] ;
 wire \add_out_d7[5] ;
 wire \add_out_d7[6] ;
 wire \add_out_d7[7] ;
 wire \add_u0._000_ ;
 wire \add_u0._001_ ;
 wire \add_u0._002_ ;
 wire \add_u0._003_ ;
 wire \add_u0._004_ ;
 wire \add_u0._005_ ;
 wire \add_u0._006_ ;
 wire \add_u0._007_ ;
 wire \add_u0._008_ ;
 wire \add_u0._009_ ;
 wire \add_u0._010_ ;
 wire \add_u0._011_ ;
 wire \add_u0._012_ ;
 wire \add_u0._013_ ;
 wire \add_u0._014_ ;
 wire \add_u0._015_ ;
 wire \add_u0._016_ ;
 wire \add_u0._017_ ;
 wire \add_u0._018_ ;
 wire \add_u0._019_ ;
 wire \add_u0._020_ ;
 wire \add_u0._021_ ;
 wire \add_u0._022_ ;
 wire \add_u0._023_ ;
 wire \add_u0._024_ ;
 wire \add_u0._025_ ;
 wire \add_u0._026_ ;
 wire \add_u0._027_ ;
 wire \add_u0._028_ ;
 wire \add_u0._029_ ;
 wire \add_u0._030_ ;
 wire \add_u0._031_ ;
 wire \add_u0._032_ ;
 wire \add_u0._033_ ;
 wire \add_u0._034_ ;
 wire \add_u0._035_ ;
 wire \add_u0._036_ ;
 wire \add_u0._037_ ;
 wire \add_u0._038_ ;
 wire \add_u0._039_ ;
 wire \add_u0._040_ ;
 wire \add_u0._041_ ;
 wire \add_u0._042_ ;
 wire \add_u0._043_ ;
 wire \add_u0._044_ ;
 wire \add_u0._045_ ;
 wire \add_u0._046_ ;
 wire \add_u0._047_ ;
 wire \add_u0._048_ ;
 wire \add_u0._049_ ;
 wire \add_u0._050_ ;
 wire \add_u0._051_ ;
 wire \add_u0._052_ ;
 wire \add_u0.a[0] ;
 wire \add_u0.a[1] ;
 wire \add_u0.a[2] ;
 wire \add_u0.a[3] ;
 wire \add_u0.a[4] ;
 wire \add_u0.a[5] ;
 wire \add_u0.a[6] ;
 wire \add_u0.a[7] ;
 wire \add_u0.a_in[0] ;
 wire \add_u0.a_in[1] ;
 wire \add_u0.a_in[2] ;
 wire \add_u0.a_in[3] ;
 wire \add_u0.a_in[4] ;
 wire \add_u0.a_in[5] ;
 wire \add_u0.a_in[6] ;
 wire \add_u0.b[0] ;
 wire \add_u0.b[1] ;
 wire \add_u0.b[2] ;
 wire \add_u0.b[3] ;
 wire \add_u0.b[4] ;
 wire \add_u0.b[5] ;
 wire \add_u0.b[6] ;
 wire \add_u0.b[7] ;
 wire \add_u0.b_in[0] ;
 wire \add_u0.b_in[1] ;
 wire \add_u0.b_in[2] ;
 wire \add_u0.b_in[3] ;
 wire \add_u0.b_in[4] ;
 wire \add_u0.b_in[5] ;
 wire \add_u0.b_in[6] ;
 wire \add_u0.c_in ;
 wire \add_u0.ppa_u0.S[0] ;
 wire \add_u0.ppa_u0.S[1] ;
 wire \add_u0.ppa_u0.S[2] ;
 wire \add_u0.ppa_u0.S[3] ;
 wire \add_u0.ppa_u0.S[4] ;
 wire \add_u0.ppa_u0.S[5] ;
 wire \add_u0.ppa_u0.S[6] ;
 wire \add_u0.ppa_u0.cg21 ;
 wire \add_u0.ppa_u0.cg43 ;
 wire \add_u0.ppa_u0.cg54 ;
 wire \add_u0.ppa_u0.cg[0] ;
 wire \add_u0.ppa_u0.cg[1] ;
 wire \add_u0.ppa_u0.cg[2] ;
 wire \add_u0.ppa_u0.cg[3] ;
 wire \add_u0.ppa_u0.cg[4] ;
 wire \add_u0.ppa_u0.cg[5] ;
 wire \add_u0.ppa_u0.cp21 ;
 wire \add_u0.ppa_u0.cp43 ;
 wire \add_u0.ppa_u0.cp54 ;
 wire \add_u0.ppa_u0.d1_0.a2._0_ ;
 wire \add_u0.ppa_u0.d1_0.a2.in0 ;
 wire \add_u0.ppa_u0.d1_0.a2.out ;
 wire \add_u0.ppa_u0.d1_0.g1 ;
 wire \add_u0.ppa_u0.d1_0.o2._0_ ;
 wire \add_u0.ppa_u0.d2_0.a2._0_ ;
 wire \add_u0.ppa_u0.d2_0.a2.in0 ;
 wire \add_u0.ppa_u0.d2_0.a2.out ;
 wire \add_u0.ppa_u0.d2_0.g1 ;
 wire \add_u0.ppa_u0.d2_0.o2._0_ ;
 wire \add_u0.ppa_u0.d3_0.a1._0_ ;
 wire \add_u0.ppa_u0.d3_0.a1.in0 ;
 wire \add_u0.ppa_u0.d3_0.a2._0_ ;
 wire \add_u0.ppa_u0.d3_0.a2.out ;
 wire \add_u0.ppa_u0.d3_0.g1 ;
 wire \add_u0.ppa_u0.d3_0.o2._0_ ;
 wire \add_u0.ppa_u0.d3_1.a2._0_ ;
 wire \add_u0.ppa_u0.d3_1.a2.out ;
 wire \add_u0.ppa_u0.d3_1.o2._0_ ;
 wire \add_u0.ppa_u0.d4_0.a2._0_ ;
 wire \add_u0.ppa_u0.d4_0.a2.in0 ;
 wire \add_u0.ppa_u0.d4_0.a2.out ;
 wire \add_u0.ppa_u0.d4_0.g1 ;
 wire \add_u0.ppa_u0.d4_0.o2._0_ ;
 wire \add_u0.ppa_u0.d5_0.a1._0_ ;
 wire \add_u0.ppa_u0.d5_0.a1.in0 ;
 wire \add_u0.ppa_u0.d5_0.a2._0_ ;
 wire \add_u0.ppa_u0.d5_0.a2.out ;
 wire \add_u0.ppa_u0.d5_0.g1 ;
 wire \add_u0.ppa_u0.d5_0.o2._0_ ;
 wire \add_u0.ppa_u0.d5_1.a2._0_ ;
 wire \add_u0.ppa_u0.d5_1.a2.out ;
 wire \add_u0.ppa_u0.d5_1.o2._0_ ;
 wire \add_u0.ppa_u0.d6_0.a1._0_ ;
 wire \add_u0.ppa_u0.d6_0.a1.in0 ;
 wire \add_u0.ppa_u0.d6_0.a2._0_ ;
 wire \add_u0.ppa_u0.d6_0.a2.out ;
 wire \add_u0.ppa_u0.d6_0.g1 ;
 wire \add_u0.ppa_u0.d6_0.o2._0_ ;
 wire \add_u0.ppa_u0.d6_1.a2._0_ ;
 wire \add_u0.ppa_u0.d6_1.a2.out ;
 wire \add_u0.ppa_u0.d6_1.o2._0_ ;
 wire \add_u0.ppa_u0.p_0.a._0_ ;
 wire \add_u0.ppa_u0.p_0.o._0_ ;
 wire \add_u0.ppa_u0.p_1.a._0_ ;
 wire \add_u0.ppa_u0.p_1.o._0_ ;
 wire \add_u0.ppa_u0.p_2.a._0_ ;
 wire \add_u0.ppa_u0.p_2.o._0_ ;
 wire \add_u0.ppa_u0.p_3.a._0_ ;
 wire \add_u0.ppa_u0.p_3.o._0_ ;
 wire \add_u0.ppa_u0.p_4.a._0_ ;
 wire \add_u0.ppa_u0.p_4.o._0_ ;
 wire \add_u0.ppa_u0.p_5.a._0_ ;
 wire \add_u0.ppa_u0.p_5.o._0_ ;
 wire \add_u0.ppa_u0.s0.temp ;
 wire \add_u0.ppa_u0.s0.xor2_0._0_ ;
 wire \add_u0.ppa_u0.s0.xor2_1._0_ ;
 wire \add_u0.ppa_u0.s1.temp ;
 wire \add_u0.ppa_u0.s1.xor2_0._0_ ;
 wire \add_u0.ppa_u0.s1.xor2_1._0_ ;
 wire \add_u0.ppa_u0.s2.temp ;
 wire \add_u0.ppa_u0.s2.xor2_0._0_ ;
 wire \add_u0.ppa_u0.s2.xor2_1._0_ ;
 wire \add_u0.ppa_u0.s3.temp ;
 wire \add_u0.ppa_u0.s3.xor2_0._0_ ;
 wire \add_u0.ppa_u0.s3.xor2_1._0_ ;
 wire \add_u0.ppa_u0.s4.temp ;
 wire \add_u0.ppa_u0.s4.xor2_0._0_ ;
 wire \add_u0.ppa_u0.s4.xor2_1._0_ ;
 wire \add_u0.ppa_u0.s5.temp ;
 wire \add_u0.ppa_u0.s5.xor2_0._0_ ;
 wire \add_u0.ppa_u0.s5.xor2_1._0_ ;
 wire \add_u0.ppa_u0.s6.temp ;
 wire \add_u0.ppa_u0.s6.xor2_0._0_ ;
 wire \add_u0.ppa_u0.s6.xor2_1._0_ ;
 wire \add_u0.sign ;
 wire \add_u0.sum[7] ;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_9_clk;
 wire \mul_out_d0[0] ;
 wire \mul_out_d0[1] ;
 wire \mul_out_d0[2] ;
 wire \mul_out_d0[3] ;
 wire \mul_out_d0[4] ;
 wire \mul_out_d0[5] ;
 wire \mul_out_d0[6] ;
 wire \mul_out_d0[7] ;
 wire \mult_add_u0._000_ ;
 wire \mult_add_u0._001_ ;
 wire \mult_add_u0._002_ ;
 wire \mult_add_u0._003_ ;
 wire \mult_add_u0._004_ ;
 wire \mult_add_u0._005_ ;
 wire \mult_add_u0._006_ ;
 wire \mult_add_u0._007_ ;
 wire \mult_add_u0._008_ ;
 wire \mult_add_u0._009_ ;
 wire \mult_add_u0._010_ ;
 wire \mult_add_u0._011_ ;
 wire \mult_add_u0._012_ ;
 wire \mult_add_u0._013_ ;
 wire \mult_add_u0._014_ ;
 wire \mult_add_u0._015_ ;
 wire \mult_add_u0._016_ ;
 wire \mult_add_u0.add0._000_ ;
 wire \mult_add_u0.add0._001_ ;
 wire \mult_add_u0.add0._002_ ;
 wire \mult_add_u0.add0._003_ ;
 wire \mult_add_u0.add0._004_ ;
 wire \mult_add_u0.add0._005_ ;
 wire \mult_add_u0.add0._006_ ;
 wire \mult_add_u0.add0._007_ ;
 wire \mult_add_u0.add0._008_ ;
 wire \mult_add_u0.add0._009_ ;
 wire \mult_add_u0.add0._010_ ;
 wire \mult_add_u0.add0._011_ ;
 wire \mult_add_u0.add0._012_ ;
 wire \mult_add_u0.add0._013_ ;
 wire \mult_add_u0.add0._014_ ;
 wire \mult_add_u0.add0._015_ ;
 wire \mult_add_u0.add0._016_ ;
 wire \mult_add_u0.add0._017_ ;
 wire \mult_add_u0.add0._018_ ;
 wire \mult_add_u0.add0._019_ ;
 wire \mult_add_u0.add0._020_ ;
 wire \mult_add_u0.add0._021_ ;
 wire \mult_add_u0.add0._022_ ;
 wire \mult_add_u0.add0._023_ ;
 wire \mult_add_u0.add0._024_ ;
 wire \mult_add_u0.add0._025_ ;
 wire \mult_add_u0.add0._026_ ;
 wire \mult_add_u0.add0._027_ ;
 wire \mult_add_u0.add0._028_ ;
 wire \mult_add_u0.add0._029_ ;
 wire \mult_add_u0.add0._030_ ;
 wire \mult_add_u0.add0._031_ ;
 wire \mult_add_u0.add0._032_ ;
 wire \mult_add_u0.add0._033_ ;
 wire \mult_add_u0.add0._034_ ;
 wire \mult_add_u0.add0._035_ ;
 wire \mult_add_u0.add0._036_ ;
 wire \mult_add_u0.add0._037_ ;
 wire \mult_add_u0.add0._038_ ;
 wire \mult_add_u0.add0._039_ ;
 wire \mult_add_u0.add0._040_ ;
 wire \mult_add_u0.add0._041_ ;
 wire \mult_add_u0.add0._042_ ;
 wire \mult_add_u0.add0._043_ ;
 wire \mult_add_u0.add0._044_ ;
 wire \mult_add_u0.add0._045_ ;
 wire \mult_add_u0.add0._046_ ;
 wire \mult_add_u0.add0._047_ ;
 wire \mult_add_u0.add0._048_ ;
 wire \mult_add_u0.add0._049_ ;
 wire \mult_add_u0.add0._050_ ;
 wire \mult_add_u0.add0._051_ ;
 wire \mult_add_u0.add0._052_ ;
 wire \mult_add_u0.add0.a[0] ;
 wire \mult_add_u0.add0.a[1] ;
 wire \mult_add_u0.add0.a[2] ;
 wire \mult_add_u0.add0.a[3] ;
 wire \mult_add_u0.add0.a[4] ;
 wire \mult_add_u0.add0.a[5] ;
 wire \mult_add_u0.add0.a[6] ;
 wire \mult_add_u0.add0.a[7] ;
 wire \mult_add_u0.add0.a_in[0] ;
 wire \mult_add_u0.add0.a_in[1] ;
 wire \mult_add_u0.add0.a_in[2] ;
 wire \mult_add_u0.add0.a_in[3] ;
 wire \mult_add_u0.add0.a_in[4] ;
 wire \mult_add_u0.add0.a_in[5] ;
 wire \mult_add_u0.add0.a_in[6] ;
 wire \mult_add_u0.add0.b[0] ;
 wire \mult_add_u0.add0.b[1] ;
 wire \mult_add_u0.add0.b[2] ;
 wire \mult_add_u0.add0.b[3] ;
 wire \mult_add_u0.add0.b[4] ;
 wire \mult_add_u0.add0.b[5] ;
 wire \mult_add_u0.add0.b[6] ;
 wire \mult_add_u0.add0.b[7] ;
 wire \mult_add_u0.add0.b_in[0] ;
 wire \mult_add_u0.add0.b_in[1] ;
 wire \mult_add_u0.add0.b_in[2] ;
 wire \mult_add_u0.add0.b_in[3] ;
 wire \mult_add_u0.add0.b_in[4] ;
 wire \mult_add_u0.add0.b_in[5] ;
 wire \mult_add_u0.add0.b_in[6] ;
 wire \mult_add_u0.add0.c_in ;
 wire \mult_add_u0.add0.ppa_u0.S[0] ;
 wire \mult_add_u0.add0.ppa_u0.S[1] ;
 wire \mult_add_u0.add0.ppa_u0.S[2] ;
 wire \mult_add_u0.add0.ppa_u0.S[3] ;
 wire \mult_add_u0.add0.ppa_u0.S[4] ;
 wire \mult_add_u0.add0.ppa_u0.S[5] ;
 wire \mult_add_u0.add0.ppa_u0.S[6] ;
 wire \mult_add_u0.add0.ppa_u0.cg21 ;
 wire \mult_add_u0.add0.ppa_u0.cg43 ;
 wire \mult_add_u0.add0.ppa_u0.cg54 ;
 wire \mult_add_u0.add0.ppa_u0.cg[0] ;
 wire \mult_add_u0.add0.ppa_u0.cg[1] ;
 wire \mult_add_u0.add0.ppa_u0.cg[2] ;
 wire \mult_add_u0.add0.ppa_u0.cg[3] ;
 wire \mult_add_u0.add0.ppa_u0.cg[4] ;
 wire \mult_add_u0.add0.ppa_u0.cg[5] ;
 wire \mult_add_u0.add0.ppa_u0.cp21 ;
 wire \mult_add_u0.add0.ppa_u0.cp43 ;
 wire \mult_add_u0.add0.ppa_u0.cp54 ;
 wire \mult_add_u0.add0.ppa_u0.d1_0.a2._0_ ;
 wire \mult_add_u0.add0.ppa_u0.d1_0.a2.in0 ;
 wire \mult_add_u0.add0.ppa_u0.d1_0.a2.out ;
 wire \mult_add_u0.add0.ppa_u0.d1_0.g1 ;
 wire \mult_add_u0.add0.ppa_u0.d1_0.o2._0_ ;
 wire \mult_add_u0.add0.ppa_u0.d2_0.a2._0_ ;
 wire \mult_add_u0.add0.ppa_u0.d2_0.a2.in0 ;
 wire \mult_add_u0.add0.ppa_u0.d2_0.a2.out ;
 wire \mult_add_u0.add0.ppa_u0.d2_0.g1 ;
 wire \mult_add_u0.add0.ppa_u0.d2_0.o2._0_ ;
 wire \mult_add_u0.add0.ppa_u0.d3_0.a1._0_ ;
 wire \mult_add_u0.add0.ppa_u0.d3_0.a1.in0 ;
 wire \mult_add_u0.add0.ppa_u0.d3_0.a2._0_ ;
 wire \mult_add_u0.add0.ppa_u0.d3_0.a2.out ;
 wire \mult_add_u0.add0.ppa_u0.d3_0.g1 ;
 wire \mult_add_u0.add0.ppa_u0.d3_0.o2._0_ ;
 wire \mult_add_u0.add0.ppa_u0.d3_1.a2._0_ ;
 wire \mult_add_u0.add0.ppa_u0.d3_1.a2.out ;
 wire \mult_add_u0.add0.ppa_u0.d3_1.o2._0_ ;
 wire \mult_add_u0.add0.ppa_u0.d4_0.a2._0_ ;
 wire \mult_add_u0.add0.ppa_u0.d4_0.a2.in0 ;
 wire \mult_add_u0.add0.ppa_u0.d4_0.a2.out ;
 wire \mult_add_u0.add0.ppa_u0.d4_0.g1 ;
 wire \mult_add_u0.add0.ppa_u0.d4_0.o2._0_ ;
 wire \mult_add_u0.add0.ppa_u0.d5_0.a1._0_ ;
 wire \mult_add_u0.add0.ppa_u0.d5_0.a1.in0 ;
 wire \mult_add_u0.add0.ppa_u0.d5_0.a2._0_ ;
 wire \mult_add_u0.add0.ppa_u0.d5_0.a2.out ;
 wire \mult_add_u0.add0.ppa_u0.d5_0.g1 ;
 wire \mult_add_u0.add0.ppa_u0.d5_0.o2._0_ ;
 wire \mult_add_u0.add0.ppa_u0.d5_1.a2._0_ ;
 wire \mult_add_u0.add0.ppa_u0.d5_1.a2.out ;
 wire \mult_add_u0.add0.ppa_u0.d5_1.o2._0_ ;
 wire \mult_add_u0.add0.ppa_u0.d6_0.a1._0_ ;
 wire \mult_add_u0.add0.ppa_u0.d6_0.a1.in0 ;
 wire \mult_add_u0.add0.ppa_u0.d6_0.a2._0_ ;
 wire \mult_add_u0.add0.ppa_u0.d6_0.a2.out ;
 wire \mult_add_u0.add0.ppa_u0.d6_0.g1 ;
 wire \mult_add_u0.add0.ppa_u0.d6_0.o2._0_ ;
 wire \mult_add_u0.add0.ppa_u0.d6_1.a2._0_ ;
 wire \mult_add_u0.add0.ppa_u0.d6_1.a2.out ;
 wire \mult_add_u0.add0.ppa_u0.d6_1.o2._0_ ;
 wire \mult_add_u0.add0.ppa_u0.p_0.a._0_ ;
 wire \mult_add_u0.add0.ppa_u0.p_0.o._0_ ;
 wire \mult_add_u0.add0.ppa_u0.p_1.a._0_ ;
 wire \mult_add_u0.add0.ppa_u0.p_1.o._0_ ;
 wire \mult_add_u0.add0.ppa_u0.p_2.a._0_ ;
 wire \mult_add_u0.add0.ppa_u0.p_2.o._0_ ;
 wire \mult_add_u0.add0.ppa_u0.p_3.a._0_ ;
 wire \mult_add_u0.add0.ppa_u0.p_3.o._0_ ;
 wire \mult_add_u0.add0.ppa_u0.p_4.a._0_ ;
 wire \mult_add_u0.add0.ppa_u0.p_4.o._0_ ;
 wire \mult_add_u0.add0.ppa_u0.p_5.a._0_ ;
 wire \mult_add_u0.add0.ppa_u0.p_5.o._0_ ;
 wire \mult_add_u0.add0.ppa_u0.s0.temp ;
 wire \mult_add_u0.add0.ppa_u0.s0.xor2_0._0_ ;
 wire \mult_add_u0.add0.ppa_u0.s0.xor2_1._0_ ;
 wire \mult_add_u0.add0.ppa_u0.s1.temp ;
 wire \mult_add_u0.add0.ppa_u0.s1.xor2_0._0_ ;
 wire \mult_add_u0.add0.ppa_u0.s1.xor2_1._0_ ;
 wire \mult_add_u0.add0.ppa_u0.s2.temp ;
 wire \mult_add_u0.add0.ppa_u0.s2.xor2_0._0_ ;
 wire \mult_add_u0.add0.ppa_u0.s2.xor2_1._0_ ;
 wire \mult_add_u0.add0.ppa_u0.s3.temp ;
 wire \mult_add_u0.add0.ppa_u0.s3.xor2_0._0_ ;
 wire \mult_add_u0.add0.ppa_u0.s3.xor2_1._0_ ;
 wire \mult_add_u0.add0.ppa_u0.s4.temp ;
 wire \mult_add_u0.add0.ppa_u0.s4.xor2_0._0_ ;
 wire \mult_add_u0.add0.ppa_u0.s4.xor2_1._0_ ;
 wire \mult_add_u0.add0.ppa_u0.s5.temp ;
 wire \mult_add_u0.add0.ppa_u0.s5.xor2_0._0_ ;
 wire \mult_add_u0.add0.ppa_u0.s5.xor2_1._0_ ;
 wire \mult_add_u0.add0.ppa_u0.s6.temp ;
 wire \mult_add_u0.add0.ppa_u0.s6.xor2_0._0_ ;
 wire \mult_add_u0.add0.ppa_u0.s6.xor2_1._0_ ;
 wire \mult_add_u0.add0.sign ;
 wire \mult_add_u0.add0.sum[7] ;
 wire \mult_add_u0.b_in[0] ;
 wire \mult_add_u0.b_in[1] ;
 wire \mult_add_u0.b_in[2] ;
 wire \mult_add_u0.b_in[3] ;
 wire \mult_add_u0.b_in[4] ;
 wire \mult_add_u0.b_in[5] ;
 wire \mult_add_u0.b_in[6] ;
 wire \mult_add_u0.b_in[7] ;
 wire \mult_add_u0.b_in_d1[0] ;
 wire \mult_add_u0.b_in_d1[1] ;
 wire \mult_add_u0.b_in_d1[2] ;
 wire \mult_add_u0.b_in_d1[3] ;
 wire \mult_add_u0.b_in_d1[4] ;
 wire \mult_add_u0.b_in_d1[5] ;
 wire \mult_add_u0.b_in_d1[6] ;
 wire \mult_add_u0.b_in_d1[7] ;
 wire \mult_add_u0.b_in_d2[0] ;
 wire \mult_add_u0.b_in_d2[1] ;
 wire \mult_add_u0.b_in_d2[2] ;
 wire \mult_add_u0.b_in_d2[3] ;
 wire \mult_add_u0.b_in_d2[4] ;
 wire \mult_add_u0.b_in_d2[5] ;
 wire \mult_add_u0.b_in_d2[6] ;
 wire \mult_add_u0.b_in_d2[7] ;
 wire \mult_add_u0.b_in_d3[0] ;
 wire \mult_add_u0.b_in_d3[1] ;
 wire \mult_add_u0.b_in_d3[2] ;
 wire \mult_add_u0.b_in_d3[3] ;
 wire \mult_add_u0.b_in_d3[4] ;
 wire \mult_add_u0.b_in_d3[5] ;
 wire \mult_add_u0.b_in_d3[6] ;
 wire \mult_add_u0.b_in_d3[7] ;
 wire \mult_add_u0.b_in_d4[0] ;
 wire \mult_add_u0.b_in_d4[1] ;
 wire \mult_add_u0.b_in_d4[2] ;
 wire \mult_add_u0.b_in_d4[3] ;
 wire \mult_add_u0.b_in_d4[4] ;
 wire \mult_add_u0.b_in_d4[5] ;
 wire \mult_add_u0.b_in_d4[6] ;
 wire \mult_add_u0.b_in_d4[7] ;
 wire \mult_add_u0.b_in_d5[0] ;
 wire \mult_add_u0.b_in_d5[1] ;
 wire \mult_add_u0.b_in_d5[2] ;
 wire \mult_add_u0.b_in_d5[3] ;
 wire \mult_add_u0.b_in_d5[4] ;
 wire \mult_add_u0.b_in_d5[5] ;
 wire \mult_add_u0.b_in_d5[6] ;
 wire \mult_add_u0.b_in_d5[7] ;
 wire \mult_add_u0.b_in_d6[0] ;
 wire \mult_add_u0.b_in_d6[1] ;
 wire \mult_add_u0.b_in_d6[2] ;
 wire \mult_add_u0.b_in_d6[3] ;
 wire \mult_add_u0.b_in_d6[4] ;
 wire \mult_add_u0.b_in_d6[5] ;
 wire \mult_add_u0.b_in_d6[6] ;
 wire \mult_add_u0.b_in_d6[7] ;
 wire \mult_add_u0.m[0] ;
 wire \mult_add_u0.m[1] ;
 wire \mult_add_u0.m[2] ;
 wire \mult_add_u0.m[3] ;
 wire \mult_add_u0.m[4] ;
 wire \mult_add_u0.m[5] ;
 wire \mult_add_u0.m[6] ;
 wire \mult_add_u0.m[7] ;
 wire \mult_add_u0.mult0.Q[0][0] ;
 wire \mult_add_u0.mult0.Q[0][1] ;
 wire \mult_add_u0.mult0.Q[0][2] ;
 wire \mult_add_u0.mult0.Q[0][3] ;
 wire \mult_add_u0.mult0.Q[0][4] ;
 wire \mult_add_u0.mult0.Q[0][5] ;
 wire \mult_add_u0.mult0.Q[1][0] ;
 wire \mult_add_u0.mult0.Q[1][1] ;
 wire \mult_add_u0.mult0.Q[1][2] ;
 wire \mult_add_u0.mult0.Q[1][3] ;
 wire \mult_add_u0.mult0.Q[1][4] ;
 wire \mult_add_u0.mult0.Q[2][0] ;
 wire \mult_add_u0.mult0.Q[2][1] ;
 wire \mult_add_u0.mult0.Q[2][2] ;
 wire \mult_add_u0.mult0.Q[2][3] ;
 wire \mult_add_u0.mult0.Q[3][0] ;
 wire \mult_add_u0.mult0.Q[3][1] ;
 wire \mult_add_u0.mult0.Q[3][2] ;
 wire \mult_add_u0.mult0.Q[3][6] ;
 wire \mult_add_u0.mult0.Q[4][0] ;
 wire \mult_add_u0.mult0.Q[4][1] ;
 wire \mult_add_u0.mult0.Q[4][5] ;
 wire \mult_add_u0.mult0.Q[4][6] ;
 wire \mult_add_u0.mult0.Q[5][0] ;
 wire \mult_add_u0.mult0.Q[5][4] ;
 wire \mult_add_u0.mult0.Q[5][5] ;
 wire \mult_add_u0.mult0.Q[5][6] ;
 wire \mult_add_u0.mult0.Q_s1[0] ;
 wire \mult_add_u0.mult0.Q_s1[1] ;
 wire \mult_add_u0.mult0.Q_s1[2] ;
 wire \mult_add_u0.mult0.Q_s1[3] ;
 wire \mult_add_u0.mult0.Q_s1[4] ;
 wire \mult_add_u0.mult0.Q_s1[5] ;
 wire \mult_add_u0.mult0.Q_s2[0] ;
 wire \mult_add_u0.mult0.Q_s2[1] ;
 wire \mult_add_u0.mult0.Q_s2[2] ;
 wire \mult_add_u0.mult0.Q_s2[3] ;
 wire \mult_add_u0.mult0.Q_s2[4] ;
 wire \mult_add_u0.mult0.Q_s3[0] ;
 wire \mult_add_u0.mult0.Q_s3[1] ;
 wire \mult_add_u0.mult0.Q_s3[2] ;
 wire \mult_add_u0.mult0.Q_s3[3] ;
 wire \mult_add_u0.mult0.Q_s4[0] ;
 wire \mult_add_u0.mult0.Q_s4[1] ;
 wire \mult_add_u0.mult0.Q_s4[2] ;
 wire \mult_add_u0.mult0.Q_s4[6] ;
 wire \mult_add_u0.mult0.Q_s5[0] ;
 wire \mult_add_u0.mult0.Q_s5[1] ;
 wire \mult_add_u0.mult0.Q_s5[5] ;
 wire \mult_add_u0.mult0.Q_s5[6] ;
 wire \mult_add_u0.mult0.Q_s6[0] ;
 wire \mult_add_u0.mult0.Q_s6[4] ;
 wire \mult_add_u0.mult0.Q_s6[5] ;
 wire \mult_add_u0.mult0.Q_s6[6] ;
 wire \mult_add_u0.mult0._000_ ;
 wire \mult_add_u0.mult0._001_ ;
 wire \mult_add_u0.mult0._002_ ;
 wire \mult_add_u0.mult0._003_ ;
 wire \mult_add_u0.mult0._004_ ;
 wire \mult_add_u0.mult0._005_ ;
 wire \mult_add_u0.mult0._006_ ;
 wire \mult_add_u0.mult0._007_ ;
 wire \mult_add_u0.mult0._008_ ;
 wire \mult_add_u0.mult0._009_ ;
 wire \mult_add_u0.mult0._010_ ;
 wire \mult_add_u0.mult0._011_ ;
 wire \mult_add_u0.mult0._012_ ;
 wire \mult_add_u0.mult0._013_ ;
 wire \mult_add_u0.mult0._014_ ;
 wire \mult_add_u0.mult0._015_ ;
 wire \mult_add_u0.mult0._016_ ;
 wire \mult_add_u0.mult0.acc[1][0] ;
 wire \mult_add_u0.mult0.acc[1][1] ;
 wire \mult_add_u0.mult0.acc[1][2] ;
 wire \mult_add_u0.mult0.acc[1][3] ;
 wire \mult_add_u0.mult0.acc[1][4] ;
 wire \mult_add_u0.mult0.acc[1][5] ;
 wire \mult_add_u0.mult0.acc[1][6] ;
 wire \mult_add_u0.mult0.acc[2][0] ;
 wire \mult_add_u0.mult0.acc[2][1] ;
 wire \mult_add_u0.mult0.acc[2][2] ;
 wire \mult_add_u0.mult0.acc[2][3] ;
 wire \mult_add_u0.mult0.acc[2][4] ;
 wire \mult_add_u0.mult0.acc[2][5] ;
 wire \mult_add_u0.mult0.acc[2][6] ;
 wire \mult_add_u0.mult0.acc[3][0] ;
 wire \mult_add_u0.mult0.acc[3][1] ;
 wire \mult_add_u0.mult0.acc[3][2] ;
 wire \mult_add_u0.mult0.acc[3][3] ;
 wire \mult_add_u0.mult0.acc[3][4] ;
 wire \mult_add_u0.mult0.acc[3][5] ;
 wire \mult_add_u0.mult0.acc[3][6] ;
 wire \mult_add_u0.mult0.acc[4][0] ;
 wire \mult_add_u0.mult0.acc[4][1] ;
 wire \mult_add_u0.mult0.acc[4][2] ;
 wire \mult_add_u0.mult0.acc[4][3] ;
 wire \mult_add_u0.mult0.acc[4][4] ;
 wire \mult_add_u0.mult0.acc[4][5] ;
 wire \mult_add_u0.mult0.acc[4][6] ;
 wire \mult_add_u0.mult0.acc[5][0] ;
 wire \mult_add_u0.mult0.acc[5][1] ;
 wire \mult_add_u0.mult0.acc[5][2] ;
 wire \mult_add_u0.mult0.acc[5][3] ;
 wire \mult_add_u0.mult0.acc[5][4] ;
 wire \mult_add_u0.mult0.acc[6][0] ;
 wire \mult_add_u0.mult0.acc[6][1] ;
 wire \mult_add_u0.mult0.acc[6][2] ;
 wire \mult_add_u0.mult0.acc[6][3] ;
 wire \mult_add_u0.mult0.acc_s1[0] ;
 wire \mult_add_u0.mult0.acc_s1[1] ;
 wire \mult_add_u0.mult0.acc_s1[2] ;
 wire \mult_add_u0.mult0.acc_s1[3] ;
 wire \mult_add_u0.mult0.acc_s1[4] ;
 wire \mult_add_u0.mult0.acc_s1[5] ;
 wire \mult_add_u0.mult0.acc_s1[6] ;
 wire \mult_add_u0.mult0.acc_s2[0] ;
 wire \mult_add_u0.mult0.acc_s2[1] ;
 wire \mult_add_u0.mult0.acc_s2[2] ;
 wire \mult_add_u0.mult0.acc_s2[3] ;
 wire \mult_add_u0.mult0.acc_s2[4] ;
 wire \mult_add_u0.mult0.acc_s2[5] ;
 wire \mult_add_u0.mult0.acc_s2[6] ;
 wire \mult_add_u0.mult0.acc_s3[0] ;
 wire \mult_add_u0.mult0.acc_s3[1] ;
 wire \mult_add_u0.mult0.acc_s3[2] ;
 wire \mult_add_u0.mult0.acc_s3[3] ;
 wire \mult_add_u0.mult0.acc_s3[4] ;
 wire \mult_add_u0.mult0.acc_s3[5] ;
 wire \mult_add_u0.mult0.acc_s3[6] ;
 wire \mult_add_u0.mult0.acc_s4[0] ;
 wire \mult_add_u0.mult0.acc_s4[1] ;
 wire \mult_add_u0.mult0.acc_s4[2] ;
 wire \mult_add_u0.mult0.acc_s4[3] ;
 wire \mult_add_u0.mult0.acc_s4[4] ;
 wire \mult_add_u0.mult0.acc_s4[5] ;
 wire \mult_add_u0.mult0.acc_s5[0] ;
 wire \mult_add_u0.mult0.acc_s5[1] ;
 wire \mult_add_u0.mult0.acc_s5[2] ;
 wire \mult_add_u0.mult0.acc_s5[3] ;
 wire \mult_add_u0.mult0.acc_s5[4] ;
 wire \mult_add_u0.mult0.acc_s6[0] ;
 wire \mult_add_u0.mult0.acc_s6[1] ;
 wire \mult_add_u0.mult0.acc_s6[2] ;
 wire \mult_add_u0.mult0.acc_s6[3] ;
 wire \mult_add_u0.mult0.mul_sign ;
 wire \mult_add_u0.mult0.mul_sign_s1 ;
 wire \mult_add_u0.mult0.mul_sign_s2 ;
 wire \mult_add_u0.mult0.mul_sign_s3 ;
 wire \mult_add_u0.mult0.mul_sign_s4 ;
 wire \mult_add_u0.mult0.mul_sign_s5 ;
 wire \mult_add_u0.mult0.mul_sign_s6 ;
 wire \mult_add_u0.mult0.multiplicand[0] ;
 wire \mult_add_u0.mult0.multiplicand[1] ;
 wire \mult_add_u0.mult0.multiplicand[2] ;
 wire \mult_add_u0.mult0.multiplicand[3] ;
 wire \mult_add_u0.mult0.multiplicand[4] ;
 wire \mult_add_u0.mult0.multiplicand[5] ;
 wire \mult_add_u0.mult0.multiplicand[6] ;
 wire \mult_add_u0.mult0.multiplicand_s1[0] ;
 wire \mult_add_u0.mult0.multiplicand_s1[1] ;
 wire \mult_add_u0.mult0.multiplicand_s1[2] ;
 wire \mult_add_u0.mult0.multiplicand_s1[3] ;
 wire \mult_add_u0.mult0.multiplicand_s1[4] ;
 wire \mult_add_u0.mult0.multiplicand_s1[5] ;
 wire \mult_add_u0.mult0.multiplicand_s1[6] ;
 wire \mult_add_u0.mult0.multiplicand_s2[0] ;
 wire \mult_add_u0.mult0.multiplicand_s2[1] ;
 wire \mult_add_u0.mult0.multiplicand_s2[2] ;
 wire \mult_add_u0.mult0.multiplicand_s2[3] ;
 wire \mult_add_u0.mult0.multiplicand_s2[4] ;
 wire \mult_add_u0.mult0.multiplicand_s2[5] ;
 wire \mult_add_u0.mult0.multiplicand_s2[6] ;
 wire \mult_add_u0.mult0.multiplicand_s3[0] ;
 wire \mult_add_u0.mult0.multiplicand_s3[1] ;
 wire \mult_add_u0.mult0.multiplicand_s3[2] ;
 wire \mult_add_u0.mult0.multiplicand_s3[3] ;
 wire \mult_add_u0.mult0.multiplicand_s3[4] ;
 wire \mult_add_u0.mult0.multiplicand_s3[5] ;
 wire \mult_add_u0.mult0.multiplicand_s3[6] ;
 wire \mult_add_u0.mult0.multiplicand_s4[0] ;
 wire \mult_add_u0.mult0.multiplicand_s4[1] ;
 wire \mult_add_u0.mult0.multiplicand_s4[2] ;
 wire \mult_add_u0.mult0.multiplicand_s4[3] ;
 wire \mult_add_u0.mult0.multiplicand_s4[4] ;
 wire \mult_add_u0.mult0.multiplicand_s4[5] ;
 wire \mult_add_u0.mult0.multiplicand_s5[0] ;
 wire \mult_add_u0.mult0.multiplicand_s5[1] ;
 wire \mult_add_u0.mult0.multiplicand_s5[2] ;
 wire \mult_add_u0.mult0.multiplicand_s5[3] ;
 wire \mult_add_u0.mult0.multiplicand_s5[4] ;
 wire \mult_add_u0.mult0.multiplicand_s6[0] ;
 wire \mult_add_u0.mult0.multiplicand_s6[1] ;
 wire \mult_add_u0.mult0.multiplicand_s6[2] ;
 wire \mult_add_u0.mult0.multiplicand_s6[3] ;
 wire \mult_add_u0.mult0.multiplier[0] ;
 wire \mult_add_u0.mult0.multiplier[1] ;
 wire \mult_add_u0.mult0.multiplier[2] ;
 wire \mult_add_u0.mult0.multiplier[3] ;
 wire \mult_add_u0.mult0.multiplier[4] ;
 wire \mult_add_u0.mult0.multiplier[5] ;
 wire \mult_add_u0.mult0.multiplier[6] ;
 wire \mult_add_u0.mult0.product[3] ;
 wire \mult_add_u0.mult0.product[4] ;
 wire \mult_add_u0.mult0.product[5] ;
 wire \mult_add_u0.mult0.product[6] ;
 wire \mult_add_u0.mult0.q0[1] ;
 wire \mult_add_u0.mult0.q0[2] ;
 wire \mult_add_u0.mult0.q0[3] ;
 wire \mult_add_u0.mult0.q0[4] ;
 wire \mult_add_u0.mult0.q0[5] ;
 wire \mult_add_u0.mult0.q0[6] ;
 wire \mult_add_u0.mult0.q0_s1 ;
 wire \mult_add_u0.mult0.q0_s2 ;
 wire \mult_add_u0.mult0.q0_s3 ;
 wire \mult_add_u0.mult0.q0_s4 ;
 wire \mult_add_u0.mult0.q0_s5 ;
 wire \mult_add_u0.mult0.q0_s6 ;
 wire \mult_add_u0.mult0.step1._00_ ;
 wire \mult_add_u0.mult0.step1._01_ ;
 wire \mult_add_u0.mult0.step1._02_ ;
 wire \mult_add_u0.mult0.step1._03_ ;
 wire \mult_add_u0.mult0.step1._04_ ;
 wire \mult_add_u0.mult0.step1._05_ ;
 wire \mult_add_u0.mult0.step1._06_ ;
 wire \mult_add_u0.mult0.step1._07_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.int_ip[0] ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.int_ip[1] ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.int_ip[2] ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.int_ip[3] ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.int_ip[4] ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.int_ip[5] ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.int_ip[6] ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.S[1] ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.S[2] ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.S[3] ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.S[4] ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.S[5] ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.S[6] ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.cg21 ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.cg43 ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.cg54 ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.cg[0] ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.cg[1] ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.cg[2] ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.cg[3] ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.cg[4] ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.cg[5] ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.cp21 ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.cp43 ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.cp54 ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d1_0.a2._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d1_0.a2.in0 ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d1_0.a2.out ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d1_0.g1 ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d1_0.o2._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d2_0.a2._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d2_0.a2.out ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d2_0.g1 ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d2_0.o2._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d3_0.a1._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d3_0.a2._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d3_0.a2.out ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d3_0.g1 ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d3_0.o2._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d3_1.a2._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d3_1.a2.out ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d3_1.o2._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d4_0.a2._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d4_0.a2.in0 ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d4_0.a2.out ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d4_0.g1 ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d4_0.o2._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d5_0.a1._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d5_0.a1.in0 ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d5_0.a2._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d5_0.a2.out ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d5_0.g1 ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d5_0.o2._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d5_1.a2._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d5_1.a2.out ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d5_1.o2._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d6_0.a1._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d6_0.a1.in0 ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d6_0.a2._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d6_0.a2.out ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d6_0.g1 ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d6_0.o2._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d6_1.a2._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d6_1.a2.out ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d6_1.o2._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_0.a._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_0.o._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_1.a._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_1.o._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_2.a._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_2.o._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_3.a._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_3.o._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_4.a._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_4.o._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_5.a._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_5.o._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s1.temp ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s1.xor2_0._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s1.xor2_1._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s2.temp ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s2.xor2_0._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s2.xor2_1._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s3.temp ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s3.xor2_0._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s3.xor2_1._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s4.temp ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s4.xor2_0._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s4.xor2_1._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s5.temp ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s5.xor2_0._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s5.xor2_1._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s6.temp ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s6.xor2_0._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s6.xor2_1._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.x0._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.x1._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.x2._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.x3._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.x4._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.x5._0_ ;
 wire \mult_add_u0.mult0.step1.add_sub4_u0.x6._0_ ;
 wire \mult_add_u0.mult0.step2._00_ ;
 wire \mult_add_u0.mult0.step2._01_ ;
 wire \mult_add_u0.mult0.step2._02_ ;
 wire \mult_add_u0.mult0.step2._03_ ;
 wire \mult_add_u0.mult0.step2._04_ ;
 wire \mult_add_u0.mult0.step2._05_ ;
 wire \mult_add_u0.mult0.step2._06_ ;
 wire \mult_add_u0.mult0.step2._07_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.int_ip[0] ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.int_ip[1] ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.int_ip[2] ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.int_ip[3] ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.int_ip[4] ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.int_ip[5] ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.int_ip[6] ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.S[1] ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.S[2] ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.S[3] ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.S[4] ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.S[5] ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.S[6] ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.cg21 ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.cg43 ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.cg54 ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.cg[0] ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.cg[1] ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.cg[2] ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.cg[3] ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.cg[4] ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.cg[5] ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.cp21 ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.cp43 ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.cp54 ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d1_0.a2._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d1_0.a2.in0 ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d1_0.a2.out ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d1_0.g1 ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d1_0.o2._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d2_0.a2._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d2_0.a2.out ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d2_0.g1 ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d2_0.o2._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d3_0.a1._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d3_0.a2._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d3_0.a2.out ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d3_0.g1 ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d3_0.o2._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d3_1.a2._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d3_1.a2.out ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d3_1.o2._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d4_0.a2._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d4_0.a2.in0 ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d4_0.a2.out ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d4_0.g1 ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d4_0.o2._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d5_0.a1._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d5_0.a1.in0 ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d5_0.a2._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d5_0.a2.out ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d5_0.g1 ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d5_0.o2._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d5_1.a2._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d5_1.a2.out ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d5_1.o2._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d6_0.a1._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d6_0.a1.in0 ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d6_0.a2._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d6_0.a2.out ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d6_0.g1 ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d6_0.o2._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d6_1.a2._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d6_1.a2.out ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d6_1.o2._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_0.a._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_0.o._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_1.a._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_1.o._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_2.a._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_2.o._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_3.a._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_3.o._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_4.a._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_4.o._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_5.a._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_5.o._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s1.temp ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s1.xor2_0._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s1.xor2_1._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s2.temp ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s2.xor2_0._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s2.xor2_1._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s3.temp ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s3.xor2_0._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s3.xor2_1._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s4.temp ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s4.xor2_0._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s4.xor2_1._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s5.temp ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s5.xor2_0._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s5.xor2_1._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s6.temp ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s6.xor2_0._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s6.xor2_1._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.x0._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.x1._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.x2._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.x3._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.x4._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.x5._0_ ;
 wire \mult_add_u0.mult0.step2.add_sub4_u0.x6._0_ ;
 wire \mult_add_u0.mult0.step3._00_ ;
 wire \mult_add_u0.mult0.step3._01_ ;
 wire \mult_add_u0.mult0.step3._02_ ;
 wire \mult_add_u0.mult0.step3._03_ ;
 wire \mult_add_u0.mult0.step3._04_ ;
 wire \mult_add_u0.mult0.step3._05_ ;
 wire \mult_add_u0.mult0.step3._06_ ;
 wire \mult_add_u0.mult0.step3._07_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.int_ip[0] ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.int_ip[1] ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.int_ip[2] ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.int_ip[3] ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.int_ip[4] ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.int_ip[5] ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.int_ip[6] ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.S[1] ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.S[2] ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.S[3] ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.S[4] ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.S[5] ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.S[6] ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.cg21 ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.cg43 ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.cg54 ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.cg[0] ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.cg[1] ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.cg[2] ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.cg[3] ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.cg[4] ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.cg[5] ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.cp21 ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.cp43 ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.cp54 ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d1_0.a2._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d1_0.a2.in0 ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d1_0.a2.out ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d1_0.g1 ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d1_0.o2._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d2_0.a2._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d2_0.a2.out ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d2_0.g1 ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d2_0.o2._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d3_0.a1._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d3_0.a2._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d3_0.a2.out ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d3_0.g1 ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d3_0.o2._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d3_1.a2._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d3_1.a2.out ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d3_1.o2._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d4_0.a2._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d4_0.a2.in0 ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d4_0.a2.out ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d4_0.g1 ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d4_0.o2._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d5_0.a1._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d5_0.a1.in0 ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d5_0.a2._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d5_0.a2.out ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d5_0.g1 ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d5_0.o2._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d5_1.a2._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d5_1.a2.out ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d5_1.o2._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d6_0.a1._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d6_0.a1.in0 ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d6_0.a2._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d6_0.a2.out ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d6_0.g1 ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d6_0.o2._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d6_1.a2._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d6_1.a2.out ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d6_1.o2._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_0.a._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_0.o._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_1.a._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_1.o._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_2.a._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_2.o._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_3.a._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_3.o._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_4.a._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_4.o._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_5.a._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_5.o._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s1.temp ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s1.xor2_0._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s1.xor2_1._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s2.temp ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s2.xor2_0._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s2.xor2_1._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s3.temp ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s3.xor2_0._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s3.xor2_1._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s4.temp ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s4.xor2_0._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s4.xor2_1._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s5.temp ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s5.xor2_0._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s5.xor2_1._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s6.temp ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s6.xor2_0._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s6.xor2_1._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.x0._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.x1._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.x2._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.x3._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.x4._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.x5._0_ ;
 wire \mult_add_u0.mult0.step3.add_sub4_u0.x6._0_ ;
 wire \mult_add_u0.mult0.step4._00_ ;
 wire \mult_add_u0.mult0.step4._01_ ;
 wire \mult_add_u0.mult0.step4._02_ ;
 wire \mult_add_u0.mult0.step4._03_ ;
 wire \mult_add_u0.mult0.step4._04_ ;
 wire \mult_add_u0.mult0.step4._05_ ;
 wire \mult_add_u0.mult0.step4._06_ ;
 wire \mult_add_u0.mult0.step4._07_ ;
 wire \mult_add_u0.mult0.step4._08_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.int_ip[0] ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.int_ip[1] ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.int_ip[2] ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.int_ip[3] ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.int_ip[4] ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.int_ip[5] ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.int_ip[6] ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.S[0] ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.S[1] ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.S[2] ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.S[3] ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.S[4] ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.S[5] ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.S[6] ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.cg21 ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.cg43 ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.cg54 ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.cg[0] ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.cg[1] ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.cg[2] ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.cg[3] ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.cg[4] ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.cg[5] ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.cp21 ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.cp43 ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.cp54 ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d1_0.a2._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d1_0.a2.in0 ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d1_0.a2.out ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d1_0.g1 ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d1_0.o2._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d2_0.a2._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d2_0.a2.out ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d2_0.g1 ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d2_0.o2._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d3_0.a1._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d3_0.a2._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d3_0.a2.out ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d3_0.g1 ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d3_0.o2._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d3_1.a2._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d3_1.a2.out ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d3_1.o2._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d4_0.a2._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d4_0.a2.in0 ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d4_0.a2.out ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d4_0.g1 ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d4_0.o2._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d5_0.a1._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d5_0.a1.in0 ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d5_0.a2._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d5_0.a2.out ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d5_0.g1 ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d5_0.o2._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d5_1.a2._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d5_1.a2.out ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d5_1.o2._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d6_0.a1._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d6_0.a1.in0 ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d6_0.a2._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d6_0.a2.out ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d6_0.g1 ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d6_0.o2._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d6_1.a2._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d6_1.a2.out ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d6_1.o2._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_0.a._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_0.o._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_1.a._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_1.o._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_2.a._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_2.o._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_3.a._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_3.o._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_4.a._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_4.o._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_5.a._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_5.o._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s0.temp ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s0.xor2_0._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s0.xor2_1._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s1.temp ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s1.xor2_0._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s1.xor2_1._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s2.temp ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s2.xor2_0._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s2.xor2_1._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s3.temp ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s3.xor2_0._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s3.xor2_1._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s4.temp ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s4.xor2_0._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s4.xor2_1._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s5.temp ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s5.xor2_0._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s5.xor2_1._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s6.temp ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s6.xor2_0._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s6.xor2_1._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.x0._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.x1._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.x2._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.x3._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.x4._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.x5._0_ ;
 wire \mult_add_u0.mult0.step4.add_sub4_u0.x6._0_ ;
 wire \mult_add_u0.mult0.step5._00_ ;
 wire \mult_add_u0.mult0.step5._01_ ;
 wire \mult_add_u0.mult0.step5._03_ ;
 wire \mult_add_u0.mult0.step5._04_ ;
 wire \mult_add_u0.mult0.step5._05_ ;
 wire \mult_add_u0.mult0.step5._06_ ;
 wire \mult_add_u0.mult0.step5._07_ ;
 wire \mult_add_u0.mult0.step5._08_ ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.int_ip[0] ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.int_ip[1] ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.int_ip[2] ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.int_ip[3] ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.int_ip[4] ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.int_ip[5] ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.S[0] ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.S[1] ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.S[2] ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.S[3] ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.S[4] ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.S[5] ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.cg21 ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.cg43 ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.cg[0] ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.cg[1] ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.cg[2] ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.cg[3] ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.cg[4] ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.cp21 ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.cp43 ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d1_0.a2._0_ ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d1_0.a2.in0 ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d1_0.a2.out ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d1_0.g1 ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d1_0.o2._0_ ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d2_0.a2._0_ ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d2_0.a2.out ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d2_0.g1 ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d2_0.o2._0_ ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d3_0.a1._0_ ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d3_0.a2._0_ ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d3_0.a2.out ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d3_0.g1 ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d3_0.o2._0_ ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d3_1.a2._0_ ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d3_1.a2.out ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d3_1.o2._0_ ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d4_0.a2._0_ ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d4_0.a2.in0 ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d4_0.a2.out ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d4_0.g1 ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d4_0.o2._0_ ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d5_0.a1._0_ ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d5_0.a1.in0 ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d5_0.a2._0_ ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d5_0.a2.out ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d5_0.g1 ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d5_0.o2._0_ ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d5_1.a2._0_ ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d5_1.a2.out ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d5_1.o2._0_ ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_0.a._0_ ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_0.o._0_ ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_1.a._0_ ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_1.o._0_ ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_2.a._0_ ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_2.o._0_ ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_3.a._0_ ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_3.o._0_ ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_4.a._0_ ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_4.o._0_ ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s0.temp ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s0.xor2_0._0_ ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s0.xor2_1._0_ ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s1.temp ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s1.xor2_0._0_ ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s1.xor2_1._0_ ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s2.temp ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s2.xor2_0._0_ ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s2.xor2_1._0_ ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s3.temp ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s3.xor2_0._0_ ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s3.xor2_1._0_ ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s4.temp ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s4.xor2_0._0_ ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s4.xor2_1._0_ ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s5.temp ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s5.xor2_0._0_ ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s5.xor2_1._0_ ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.x0._0_ ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.x1._0_ ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.x2._0_ ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.x3._0_ ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.x4._0_ ;
 wire \mult_add_u0.mult0.step5.add_sub4_u0.x5._0_ ;
 wire \mult_add_u0.mult0.step6._00_ ;
 wire \mult_add_u0.mult0.step6._01_ ;
 wire \mult_add_u0.mult0.step6._03_ ;
 wire \mult_add_u0.mult0.step6._04_ ;
 wire \mult_add_u0.mult0.step6._05_ ;
 wire \mult_add_u0.mult0.step6._06_ ;
 wire \mult_add_u0.mult0.step6._08_ ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.int_ip[0] ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.int_ip[1] ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.int_ip[2] ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.int_ip[3] ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.int_ip[4] ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.S[0] ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.S[1] ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.S[2] ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.S[3] ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.S[4] ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.cg21 ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.cg[0] ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.cg[1] ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.cg[2] ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.cg[3] ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.cp21 ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d1_0.a2._0_ ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d1_0.a2.in0 ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d1_0.a2.out ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d1_0.g1 ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d1_0.o2._0_ ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d2_0.a2._0_ ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d2_0.a2.out ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d2_0.g1 ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d2_0.o2._0_ ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d3_0.a1._0_ ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d3_0.a2._0_ ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d3_0.a2.out ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d3_0.g1 ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d3_0.o2._0_ ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d3_1.a2._0_ ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d3_1.a2.out ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d3_1.o2._0_ ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d4_0.a2._0_ ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d4_0.a2.in0 ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d4_0.a2.out ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d4_0.g1 ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d4_0.o2._0_ ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.p_0.a._0_ ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.p_0.o._0_ ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.p_1.a._0_ ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.p_1.o._0_ ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.p_2.a._0_ ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.p_2.o._0_ ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.p_3.a._0_ ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.p_3.o._0_ ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s0.temp ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s0.xor2_0._0_ ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s0.xor2_1._0_ ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s1.temp ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s1.xor2_0._0_ ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s1.xor2_1._0_ ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s2.temp ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s2.xor2_0._0_ ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s2.xor2_1._0_ ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s3.temp ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s3.xor2_0._0_ ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s3.xor2_1._0_ ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s4.temp ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s4.xor2_0._0_ ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s4.xor2_1._0_ ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.x0._0_ ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.x1._0_ ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.x2._0_ ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.x3._0_ ;
 wire \mult_add_u0.mult0.step6.add_sub4_u0.x4._0_ ;
 wire \mult_add_u0.mult0.step7._00_ ;
 wire \mult_add_u0.mult0.step7._01_ ;
 wire \mult_add_u0.mult0.step7._03_ ;
 wire \mult_add_u0.mult0.step7._04_ ;
 wire \mult_add_u0.mult0.step7._05_ ;
 wire \mult_add_u0.mult0.step7._08_ ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.int_ip[0] ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.int_ip[1] ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.int_ip[2] ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.int_ip[3] ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.S[0] ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.S[1] ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.S[2] ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.S[3] ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.cg21 ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.cg[0] ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.cg[1] ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.cg[2] ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.cp21 ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d1_0.a2._0_ ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d1_0.a2.in0 ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d1_0.a2.out ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d1_0.g1 ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d1_0.o2._0_ ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d2_0.a2._0_ ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d2_0.a2.out ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d2_0.g1 ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d2_0.o2._0_ ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d3_0.a1._0_ ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d3_0.a2._0_ ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d3_0.a2.out ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d3_0.g1 ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d3_0.o2._0_ ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d3_1.a2._0_ ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d3_1.a2.out ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d3_1.o2._0_ ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.p_0.a._0_ ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.p_0.o._0_ ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.p_1.a._0_ ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.p_1.o._0_ ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.p_2.a._0_ ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.p_2.o._0_ ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s0.temp ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s0.xor2_0._0_ ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s0.xor2_1._0_ ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s1.temp ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s1.xor2_0._0_ ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s1.xor2_1._0_ ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s2.temp ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s2.xor2_0._0_ ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s2.xor2_1._0_ ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s3.temp ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s3.xor2_0._0_ ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s3.xor2_1._0_ ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.x0._0_ ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.x1._0_ ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.x2._0_ ;
 wire \mult_add_u0.mult0.step7.add_sub4_u0.x3._0_ ;
 wire \mult_add_u0.mult0.step7.next_acc[0] ;
 wire \mult_add_u0.mult0.step7.next_acc[1] ;
 wire \mult_add_u0.mult0.step7.next_acc[2] ;
 wire \mult_add_u0.mult0.x_sign._0_ ;
 wire \mult_add_u0.out[0] ;
 wire \mult_add_u0.out[1] ;
 wire \mult_add_u0.out[2] ;
 wire \mult_add_u0.out[3] ;
 wire \mult_add_u0.out[4] ;
 wire \mult_add_u0.out[5] ;
 wire \mult_add_u0.out[6] ;
 wire \mult_add_u0.out[7] ;
 wire \mult_u0.Q[0][0] ;
 wire \mult_u0.Q[0][1] ;
 wire \mult_u0.Q[0][2] ;
 wire \mult_u0.Q[0][3] ;
 wire \mult_u0.Q[0][4] ;
 wire \mult_u0.Q[0][5] ;
 wire \mult_u0.Q[1][0] ;
 wire \mult_u0.Q[1][1] ;
 wire \mult_u0.Q[1][2] ;
 wire \mult_u0.Q[1][3] ;
 wire \mult_u0.Q[1][4] ;
 wire \mult_u0.Q[2][0] ;
 wire \mult_u0.Q[2][1] ;
 wire \mult_u0.Q[2][2] ;
 wire \mult_u0.Q[2][3] ;
 wire \mult_u0.Q[3][0] ;
 wire \mult_u0.Q[3][1] ;
 wire \mult_u0.Q[3][2] ;
 wire \mult_u0.Q[3][6] ;
 wire \mult_u0.Q[4][0] ;
 wire \mult_u0.Q[4][1] ;
 wire \mult_u0.Q[4][5] ;
 wire \mult_u0.Q[4][6] ;
 wire \mult_u0.Q[5][0] ;
 wire \mult_u0.Q[5][4] ;
 wire \mult_u0.Q[5][5] ;
 wire \mult_u0.Q[5][6] ;
 wire \mult_u0.Q_s1[0] ;
 wire \mult_u0.Q_s1[1] ;
 wire \mult_u0.Q_s1[2] ;
 wire \mult_u0.Q_s1[3] ;
 wire \mult_u0.Q_s1[4] ;
 wire \mult_u0.Q_s1[5] ;
 wire \mult_u0.Q_s2[0] ;
 wire \mult_u0.Q_s2[1] ;
 wire \mult_u0.Q_s2[2] ;
 wire \mult_u0.Q_s2[3] ;
 wire \mult_u0.Q_s2[4] ;
 wire \mult_u0.Q_s3[0] ;
 wire \mult_u0.Q_s3[1] ;
 wire \mult_u0.Q_s3[2] ;
 wire \mult_u0.Q_s3[3] ;
 wire \mult_u0.Q_s4[0] ;
 wire \mult_u0.Q_s4[1] ;
 wire \mult_u0.Q_s4[2] ;
 wire \mult_u0.Q_s4[6] ;
 wire \mult_u0.Q_s5[0] ;
 wire \mult_u0.Q_s5[1] ;
 wire \mult_u0.Q_s5[5] ;
 wire \mult_u0.Q_s5[6] ;
 wire \mult_u0.Q_s6[0] ;
 wire \mult_u0.Q_s6[4] ;
 wire \mult_u0.Q_s6[5] ;
 wire \mult_u0.Q_s6[6] ;
 wire \mult_u0._000_ ;
 wire \mult_u0._001_ ;
 wire \mult_u0._002_ ;
 wire \mult_u0._003_ ;
 wire \mult_u0._004_ ;
 wire \mult_u0._005_ ;
 wire \mult_u0._006_ ;
 wire \mult_u0._007_ ;
 wire \mult_u0._008_ ;
 wire \mult_u0._009_ ;
 wire \mult_u0._010_ ;
 wire \mult_u0._011_ ;
 wire \mult_u0._012_ ;
 wire \mult_u0._013_ ;
 wire \mult_u0._014_ ;
 wire \mult_u0._015_ ;
 wire \mult_u0._016_ ;
 wire \mult_u0.acc[1][0] ;
 wire \mult_u0.acc[1][1] ;
 wire \mult_u0.acc[1][2] ;
 wire \mult_u0.acc[1][3] ;
 wire \mult_u0.acc[1][4] ;
 wire \mult_u0.acc[1][5] ;
 wire \mult_u0.acc[1][6] ;
 wire \mult_u0.acc[2][0] ;
 wire \mult_u0.acc[2][1] ;
 wire \mult_u0.acc[2][2] ;
 wire \mult_u0.acc[2][3] ;
 wire \mult_u0.acc[2][4] ;
 wire \mult_u0.acc[2][5] ;
 wire \mult_u0.acc[2][6] ;
 wire \mult_u0.acc[3][0] ;
 wire \mult_u0.acc[3][1] ;
 wire \mult_u0.acc[3][2] ;
 wire \mult_u0.acc[3][3] ;
 wire \mult_u0.acc[3][4] ;
 wire \mult_u0.acc[3][5] ;
 wire \mult_u0.acc[3][6] ;
 wire \mult_u0.acc[4][0] ;
 wire \mult_u0.acc[4][1] ;
 wire \mult_u0.acc[4][2] ;
 wire \mult_u0.acc[4][3] ;
 wire \mult_u0.acc[4][4] ;
 wire \mult_u0.acc[4][5] ;
 wire \mult_u0.acc[4][6] ;
 wire \mult_u0.acc[5][0] ;
 wire \mult_u0.acc[5][1] ;
 wire \mult_u0.acc[5][2] ;
 wire \mult_u0.acc[5][3] ;
 wire \mult_u0.acc[5][4] ;
 wire \mult_u0.acc[6][0] ;
 wire \mult_u0.acc[6][1] ;
 wire \mult_u0.acc[6][2] ;
 wire \mult_u0.acc[6][3] ;
 wire \mult_u0.acc_s1[0] ;
 wire \mult_u0.acc_s1[1] ;
 wire \mult_u0.acc_s1[2] ;
 wire \mult_u0.acc_s1[3] ;
 wire \mult_u0.acc_s1[4] ;
 wire \mult_u0.acc_s1[5] ;
 wire \mult_u0.acc_s1[6] ;
 wire \mult_u0.acc_s2[0] ;
 wire \mult_u0.acc_s2[1] ;
 wire \mult_u0.acc_s2[2] ;
 wire \mult_u0.acc_s2[3] ;
 wire \mult_u0.acc_s2[4] ;
 wire \mult_u0.acc_s2[5] ;
 wire \mult_u0.acc_s2[6] ;
 wire \mult_u0.acc_s3[0] ;
 wire \mult_u0.acc_s3[1] ;
 wire \mult_u0.acc_s3[2] ;
 wire \mult_u0.acc_s3[3] ;
 wire \mult_u0.acc_s3[4] ;
 wire \mult_u0.acc_s3[5] ;
 wire \mult_u0.acc_s3[6] ;
 wire \mult_u0.acc_s4[0] ;
 wire \mult_u0.acc_s4[1] ;
 wire \mult_u0.acc_s4[2] ;
 wire \mult_u0.acc_s4[3] ;
 wire \mult_u0.acc_s4[4] ;
 wire \mult_u0.acc_s4[5] ;
 wire \mult_u0.acc_s5[0] ;
 wire \mult_u0.acc_s5[1] ;
 wire \mult_u0.acc_s5[2] ;
 wire \mult_u0.acc_s5[3] ;
 wire \mult_u0.acc_s5[4] ;
 wire \mult_u0.acc_s6[0] ;
 wire \mult_u0.acc_s6[1] ;
 wire \mult_u0.acc_s6[2] ;
 wire \mult_u0.acc_s6[3] ;
 wire \mult_u0.mul_sign ;
 wire \mult_u0.mul_sign_s1 ;
 wire \mult_u0.mul_sign_s2 ;
 wire \mult_u0.mul_sign_s3 ;
 wire \mult_u0.mul_sign_s4 ;
 wire \mult_u0.mul_sign_s5 ;
 wire \mult_u0.mul_sign_s6 ;
 wire \mult_u0.multiplicand[0] ;
 wire \mult_u0.multiplicand[1] ;
 wire \mult_u0.multiplicand[2] ;
 wire \mult_u0.multiplicand[3] ;
 wire \mult_u0.multiplicand[4] ;
 wire \mult_u0.multiplicand[5] ;
 wire \mult_u0.multiplicand[6] ;
 wire \mult_u0.multiplicand_s1[0] ;
 wire \mult_u0.multiplicand_s1[1] ;
 wire \mult_u0.multiplicand_s1[2] ;
 wire \mult_u0.multiplicand_s1[3] ;
 wire \mult_u0.multiplicand_s1[4] ;
 wire \mult_u0.multiplicand_s1[5] ;
 wire \mult_u0.multiplicand_s1[6] ;
 wire \mult_u0.multiplicand_s2[0] ;
 wire \mult_u0.multiplicand_s2[1] ;
 wire \mult_u0.multiplicand_s2[2] ;
 wire \mult_u0.multiplicand_s2[3] ;
 wire \mult_u0.multiplicand_s2[4] ;
 wire \mult_u0.multiplicand_s2[5] ;
 wire \mult_u0.multiplicand_s2[6] ;
 wire \mult_u0.multiplicand_s3[0] ;
 wire \mult_u0.multiplicand_s3[1] ;
 wire \mult_u0.multiplicand_s3[2] ;
 wire \mult_u0.multiplicand_s3[3] ;
 wire \mult_u0.multiplicand_s3[4] ;
 wire \mult_u0.multiplicand_s3[5] ;
 wire \mult_u0.multiplicand_s3[6] ;
 wire \mult_u0.multiplicand_s4[0] ;
 wire \mult_u0.multiplicand_s4[1] ;
 wire \mult_u0.multiplicand_s4[2] ;
 wire \mult_u0.multiplicand_s4[3] ;
 wire \mult_u0.multiplicand_s4[4] ;
 wire \mult_u0.multiplicand_s4[5] ;
 wire \mult_u0.multiplicand_s5[0] ;
 wire \mult_u0.multiplicand_s5[1] ;
 wire \mult_u0.multiplicand_s5[2] ;
 wire \mult_u0.multiplicand_s5[3] ;
 wire \mult_u0.multiplicand_s5[4] ;
 wire \mult_u0.multiplicand_s6[0] ;
 wire \mult_u0.multiplicand_s6[1] ;
 wire \mult_u0.multiplicand_s6[2] ;
 wire \mult_u0.multiplicand_s6[3] ;
 wire \mult_u0.multiplier[0] ;
 wire \mult_u0.multiplier[1] ;
 wire \mult_u0.multiplier[2] ;
 wire \mult_u0.multiplier[3] ;
 wire \mult_u0.multiplier[4] ;
 wire \mult_u0.multiplier[5] ;
 wire \mult_u0.multiplier[6] ;
 wire \mult_u0.product[3] ;
 wire \mult_u0.product[4] ;
 wire \mult_u0.product[5] ;
 wire \mult_u0.product[6] ;
 wire \mult_u0.product_r[0] ;
 wire \mult_u0.product_r[1] ;
 wire \mult_u0.product_r[2] ;
 wire \mult_u0.product_r[3] ;
 wire \mult_u0.product_r[4] ;
 wire \mult_u0.product_r[5] ;
 wire \mult_u0.product_r[6] ;
 wire \mult_u0.product_r[7] ;
 wire \mult_u0.q0[1] ;
 wire \mult_u0.q0[2] ;
 wire \mult_u0.q0[3] ;
 wire \mult_u0.q0[4] ;
 wire \mult_u0.q0[5] ;
 wire \mult_u0.q0[6] ;
 wire \mult_u0.q0_s1 ;
 wire \mult_u0.q0_s2 ;
 wire \mult_u0.q0_s3 ;
 wire \mult_u0.q0_s4 ;
 wire \mult_u0.q0_s5 ;
 wire \mult_u0.q0_s6 ;
 wire \mult_u0.step1._00_ ;
 wire \mult_u0.step1._01_ ;
 wire \mult_u0.step1._02_ ;
 wire \mult_u0.step1._03_ ;
 wire \mult_u0.step1._04_ ;
 wire \mult_u0.step1._05_ ;
 wire \mult_u0.step1._06_ ;
 wire \mult_u0.step1._07_ ;
 wire \mult_u0.step1.add_sub4_u0.int_ip[0] ;
 wire \mult_u0.step1.add_sub4_u0.int_ip[1] ;
 wire \mult_u0.step1.add_sub4_u0.int_ip[2] ;
 wire \mult_u0.step1.add_sub4_u0.int_ip[3] ;
 wire \mult_u0.step1.add_sub4_u0.int_ip[4] ;
 wire \mult_u0.step1.add_sub4_u0.int_ip[5] ;
 wire \mult_u0.step1.add_sub4_u0.int_ip[6] ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.S[1] ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.S[2] ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.S[3] ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.S[4] ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.S[5] ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.S[6] ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.cg21 ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.cg43 ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.cg54 ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.cg[0] ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.cg[1] ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.cg[2] ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.cg[3] ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.cg[4] ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.cg[5] ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.cp21 ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.cp43 ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.cp54 ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.d1_0.a2._0_ ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.d1_0.a2.in0 ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.d1_0.a2.out ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.d1_0.g1 ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.d1_0.o2._0_ ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.d2_0.a2._0_ ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.d2_0.a2.out ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.d2_0.g1 ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.d2_0.o2._0_ ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.d3_0.a1._0_ ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.d3_0.a2._0_ ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.d3_0.a2.out ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.d3_0.g1 ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.d3_0.o2._0_ ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.d3_1.a2._0_ ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.d3_1.a2.out ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.d3_1.o2._0_ ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.d4_0.a2._0_ ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.d4_0.a2.in0 ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.d4_0.a2.out ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.d4_0.g1 ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.d4_0.o2._0_ ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.d5_0.a1._0_ ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.d5_0.a1.in0 ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.d5_0.a2._0_ ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.d5_0.a2.out ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.d5_0.g1 ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.d5_0.o2._0_ ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.d5_1.a2._0_ ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.d5_1.a2.out ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.d5_1.o2._0_ ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.d6_0.a1._0_ ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.d6_0.a1.in0 ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.d6_0.a2._0_ ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.d6_0.a2.out ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.d6_0.g1 ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.d6_0.o2._0_ ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.d6_1.a2._0_ ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.d6_1.a2.out ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.d6_1.o2._0_ ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.p_0.a._0_ ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.p_0.o._0_ ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.p_1.a._0_ ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.p_1.o._0_ ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.p_2.a._0_ ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.p_2.o._0_ ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.p_3.a._0_ ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.p_3.o._0_ ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.p_4.a._0_ ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.p_4.o._0_ ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.p_5.a._0_ ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.p_5.o._0_ ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.s1.temp ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.s1.xor2_0._0_ ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.s1.xor2_1._0_ ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.s2.temp ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.s2.xor2_0._0_ ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.s2.xor2_1._0_ ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.s3.temp ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.s3.xor2_0._0_ ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.s3.xor2_1._0_ ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.s4.temp ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.s4.xor2_0._0_ ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.s4.xor2_1._0_ ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.s5.temp ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.s5.xor2_0._0_ ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.s5.xor2_1._0_ ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.s6.temp ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.s6.xor2_0._0_ ;
 wire \mult_u0.step1.add_sub4_u0.ppa8_u0.s6.xor2_1._0_ ;
 wire \mult_u0.step1.add_sub4_u0.x0._0_ ;
 wire \mult_u0.step1.add_sub4_u0.x1._0_ ;
 wire \mult_u0.step1.add_sub4_u0.x2._0_ ;
 wire \mult_u0.step1.add_sub4_u0.x3._0_ ;
 wire \mult_u0.step1.add_sub4_u0.x4._0_ ;
 wire \mult_u0.step1.add_sub4_u0.x5._0_ ;
 wire \mult_u0.step1.add_sub4_u0.x6._0_ ;
 wire \mult_u0.step2._00_ ;
 wire \mult_u0.step2._01_ ;
 wire \mult_u0.step2._02_ ;
 wire \mult_u0.step2._03_ ;
 wire \mult_u0.step2._04_ ;
 wire \mult_u0.step2._05_ ;
 wire \mult_u0.step2._06_ ;
 wire \mult_u0.step2._07_ ;
 wire \mult_u0.step2.add_sub4_u0.int_ip[0] ;
 wire \mult_u0.step2.add_sub4_u0.int_ip[1] ;
 wire \mult_u0.step2.add_sub4_u0.int_ip[2] ;
 wire \mult_u0.step2.add_sub4_u0.int_ip[3] ;
 wire \mult_u0.step2.add_sub4_u0.int_ip[4] ;
 wire \mult_u0.step2.add_sub4_u0.int_ip[5] ;
 wire \mult_u0.step2.add_sub4_u0.int_ip[6] ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.S[1] ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.S[2] ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.S[3] ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.S[4] ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.S[5] ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.S[6] ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.cg21 ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.cg43 ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.cg54 ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.cg[0] ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.cg[1] ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.cg[2] ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.cg[3] ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.cg[4] ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.cg[5] ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.cp21 ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.cp43 ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.cp54 ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.d1_0.a2._0_ ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.d1_0.a2.in0 ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.d1_0.a2.out ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.d1_0.g1 ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.d1_0.o2._0_ ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.d2_0.a2._0_ ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.d2_0.a2.out ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.d2_0.g1 ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.d2_0.o2._0_ ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.d3_0.a1._0_ ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.d3_0.a2._0_ ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.d3_0.a2.out ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.d3_0.g1 ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.d3_0.o2._0_ ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.d3_1.a2._0_ ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.d3_1.a2.out ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.d3_1.o2._0_ ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.d4_0.a2._0_ ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.d4_0.a2.in0 ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.d4_0.a2.out ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.d4_0.g1 ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.d4_0.o2._0_ ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.d5_0.a1._0_ ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.d5_0.a1.in0 ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.d5_0.a2._0_ ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.d5_0.a2.out ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.d5_0.g1 ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.d5_0.o2._0_ ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.d5_1.a2._0_ ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.d5_1.a2.out ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.d5_1.o2._0_ ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.d6_0.a1._0_ ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.d6_0.a1.in0 ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.d6_0.a2._0_ ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.d6_0.a2.out ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.d6_0.g1 ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.d6_0.o2._0_ ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.d6_1.a2._0_ ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.d6_1.a2.out ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.d6_1.o2._0_ ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.p_0.a._0_ ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.p_0.o._0_ ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.p_1.a._0_ ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.p_1.o._0_ ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.p_2.a._0_ ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.p_2.o._0_ ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.p_3.a._0_ ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.p_3.o._0_ ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.p_4.a._0_ ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.p_4.o._0_ ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.p_5.a._0_ ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.p_5.o._0_ ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.s1.temp ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.s1.xor2_0._0_ ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.s1.xor2_1._0_ ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.s2.temp ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.s2.xor2_0._0_ ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.s2.xor2_1._0_ ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.s3.temp ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.s3.xor2_0._0_ ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.s3.xor2_1._0_ ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.s4.temp ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.s4.xor2_0._0_ ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.s4.xor2_1._0_ ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.s5.temp ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.s5.xor2_0._0_ ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.s5.xor2_1._0_ ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.s6.temp ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.s6.xor2_0._0_ ;
 wire \mult_u0.step2.add_sub4_u0.ppa8_u0.s6.xor2_1._0_ ;
 wire \mult_u0.step2.add_sub4_u0.x0._0_ ;
 wire \mult_u0.step2.add_sub4_u0.x1._0_ ;
 wire \mult_u0.step2.add_sub4_u0.x2._0_ ;
 wire \mult_u0.step2.add_sub4_u0.x3._0_ ;
 wire \mult_u0.step2.add_sub4_u0.x4._0_ ;
 wire \mult_u0.step2.add_sub4_u0.x5._0_ ;
 wire \mult_u0.step2.add_sub4_u0.x6._0_ ;
 wire \mult_u0.step3._00_ ;
 wire \mult_u0.step3._01_ ;
 wire \mult_u0.step3._02_ ;
 wire \mult_u0.step3._03_ ;
 wire \mult_u0.step3._04_ ;
 wire \mult_u0.step3._05_ ;
 wire \mult_u0.step3._06_ ;
 wire \mult_u0.step3._07_ ;
 wire \mult_u0.step3.add_sub4_u0.int_ip[0] ;
 wire \mult_u0.step3.add_sub4_u0.int_ip[1] ;
 wire \mult_u0.step3.add_sub4_u0.int_ip[2] ;
 wire \mult_u0.step3.add_sub4_u0.int_ip[3] ;
 wire \mult_u0.step3.add_sub4_u0.int_ip[4] ;
 wire \mult_u0.step3.add_sub4_u0.int_ip[5] ;
 wire \mult_u0.step3.add_sub4_u0.int_ip[6] ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.S[1] ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.S[2] ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.S[3] ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.S[4] ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.S[5] ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.S[6] ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.cg21 ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.cg43 ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.cg54 ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.cg[0] ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.cg[1] ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.cg[2] ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.cg[3] ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.cg[4] ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.cg[5] ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.cp21 ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.cp43 ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.cp54 ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.d1_0.a2._0_ ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.d1_0.a2.in0 ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.d1_0.a2.out ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.d1_0.g1 ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.d1_0.o2._0_ ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.d2_0.a2._0_ ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.d2_0.a2.out ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.d2_0.g1 ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.d2_0.o2._0_ ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.d3_0.a1._0_ ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.d3_0.a2._0_ ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.d3_0.a2.out ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.d3_0.g1 ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.d3_0.o2._0_ ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.d3_1.a2._0_ ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.d3_1.a2.out ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.d3_1.o2._0_ ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.d4_0.a2._0_ ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.d4_0.a2.in0 ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.d4_0.a2.out ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.d4_0.g1 ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.d4_0.o2._0_ ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.d5_0.a1._0_ ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.d5_0.a1.in0 ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.d5_0.a2._0_ ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.d5_0.a2.out ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.d5_0.g1 ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.d5_0.o2._0_ ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.d5_1.a2._0_ ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.d5_1.a2.out ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.d5_1.o2._0_ ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.d6_0.a1._0_ ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.d6_0.a1.in0 ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.d6_0.a2._0_ ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.d6_0.a2.out ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.d6_0.g1 ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.d6_0.o2._0_ ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.d6_1.a2._0_ ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.d6_1.a2.out ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.d6_1.o2._0_ ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.p_0.a._0_ ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.p_0.o._0_ ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.p_1.a._0_ ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.p_1.o._0_ ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.p_2.a._0_ ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.p_2.o._0_ ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.p_3.a._0_ ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.p_3.o._0_ ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.p_4.a._0_ ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.p_4.o._0_ ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.p_5.a._0_ ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.p_5.o._0_ ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.s1.temp ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.s1.xor2_0._0_ ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.s1.xor2_1._0_ ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.s2.temp ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.s2.xor2_0._0_ ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.s2.xor2_1._0_ ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.s3.temp ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.s3.xor2_0._0_ ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.s3.xor2_1._0_ ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.s4.temp ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.s4.xor2_0._0_ ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.s4.xor2_1._0_ ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.s5.temp ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.s5.xor2_0._0_ ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.s5.xor2_1._0_ ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.s6.temp ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.s6.xor2_0._0_ ;
 wire \mult_u0.step3.add_sub4_u0.ppa8_u0.s6.xor2_1._0_ ;
 wire \mult_u0.step3.add_sub4_u0.x0._0_ ;
 wire \mult_u0.step3.add_sub4_u0.x1._0_ ;
 wire \mult_u0.step3.add_sub4_u0.x2._0_ ;
 wire \mult_u0.step3.add_sub4_u0.x3._0_ ;
 wire \mult_u0.step3.add_sub4_u0.x4._0_ ;
 wire \mult_u0.step3.add_sub4_u0.x5._0_ ;
 wire \mult_u0.step3.add_sub4_u0.x6._0_ ;
 wire \mult_u0.step4._00_ ;
 wire \mult_u0.step4._01_ ;
 wire \mult_u0.step4._02_ ;
 wire \mult_u0.step4._03_ ;
 wire \mult_u0.step4._04_ ;
 wire \mult_u0.step4._05_ ;
 wire \mult_u0.step4._06_ ;
 wire \mult_u0.step4._07_ ;
 wire \mult_u0.step4._08_ ;
 wire \mult_u0.step4.add_sub4_u0.int_ip[0] ;
 wire \mult_u0.step4.add_sub4_u0.int_ip[1] ;
 wire \mult_u0.step4.add_sub4_u0.int_ip[2] ;
 wire \mult_u0.step4.add_sub4_u0.int_ip[3] ;
 wire \mult_u0.step4.add_sub4_u0.int_ip[4] ;
 wire \mult_u0.step4.add_sub4_u0.int_ip[5] ;
 wire \mult_u0.step4.add_sub4_u0.int_ip[6] ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.S[0] ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.S[1] ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.S[2] ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.S[3] ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.S[4] ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.S[5] ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.S[6] ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.cg21 ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.cg43 ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.cg54 ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.cg[0] ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.cg[1] ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.cg[2] ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.cg[3] ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.cg[4] ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.cg[5] ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.cp21 ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.cp43 ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.cp54 ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.d1_0.a2._0_ ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.d1_0.a2.in0 ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.d1_0.a2.out ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.d1_0.g1 ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.d1_0.o2._0_ ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.d2_0.a2._0_ ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.d2_0.a2.out ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.d2_0.g1 ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.d2_0.o2._0_ ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.d3_0.a1._0_ ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.d3_0.a2._0_ ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.d3_0.a2.out ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.d3_0.g1 ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.d3_0.o2._0_ ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.d3_1.a2._0_ ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.d3_1.a2.out ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.d3_1.o2._0_ ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.d4_0.a2._0_ ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.d4_0.a2.in0 ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.d4_0.a2.out ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.d4_0.g1 ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.d4_0.o2._0_ ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.d5_0.a1._0_ ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.d5_0.a1.in0 ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.d5_0.a2._0_ ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.d5_0.a2.out ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.d5_0.g1 ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.d5_0.o2._0_ ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.d5_1.a2._0_ ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.d5_1.a2.out ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.d5_1.o2._0_ ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.d6_0.a1._0_ ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.d6_0.a1.in0 ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.d6_0.a2._0_ ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.d6_0.a2.out ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.d6_0.g1 ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.d6_0.o2._0_ ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.d6_1.a2._0_ ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.d6_1.a2.out ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.d6_1.o2._0_ ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.p_0.a._0_ ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.p_0.o._0_ ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.p_1.a._0_ ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.p_1.o._0_ ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.p_2.a._0_ ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.p_2.o._0_ ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.p_3.a._0_ ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.p_3.o._0_ ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.p_4.a._0_ ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.p_4.o._0_ ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.p_5.a._0_ ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.p_5.o._0_ ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.s0.temp ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.s0.xor2_0._0_ ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.s0.xor2_1._0_ ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.s1.temp ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.s1.xor2_0._0_ ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.s1.xor2_1._0_ ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.s2.temp ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.s2.xor2_0._0_ ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.s2.xor2_1._0_ ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.s3.temp ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.s3.xor2_0._0_ ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.s3.xor2_1._0_ ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.s4.temp ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.s4.xor2_0._0_ ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.s4.xor2_1._0_ ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.s5.temp ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.s5.xor2_0._0_ ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.s5.xor2_1._0_ ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.s6.temp ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.s6.xor2_0._0_ ;
 wire \mult_u0.step4.add_sub4_u0.ppa8_u0.s6.xor2_1._0_ ;
 wire \mult_u0.step4.add_sub4_u0.x0._0_ ;
 wire \mult_u0.step4.add_sub4_u0.x1._0_ ;
 wire \mult_u0.step4.add_sub4_u0.x2._0_ ;
 wire \mult_u0.step4.add_sub4_u0.x3._0_ ;
 wire \mult_u0.step4.add_sub4_u0.x4._0_ ;
 wire \mult_u0.step4.add_sub4_u0.x5._0_ ;
 wire \mult_u0.step4.add_sub4_u0.x6._0_ ;
 wire \mult_u0.step5._00_ ;
 wire \mult_u0.step5._01_ ;
 wire \mult_u0.step5._03_ ;
 wire \mult_u0.step5._04_ ;
 wire \mult_u0.step5._05_ ;
 wire \mult_u0.step5._06_ ;
 wire \mult_u0.step5._07_ ;
 wire \mult_u0.step5._08_ ;
 wire \mult_u0.step5.add_sub4_u0.int_ip[0] ;
 wire \mult_u0.step5.add_sub4_u0.int_ip[1] ;
 wire \mult_u0.step5.add_sub4_u0.int_ip[2] ;
 wire \mult_u0.step5.add_sub4_u0.int_ip[3] ;
 wire \mult_u0.step5.add_sub4_u0.int_ip[4] ;
 wire \mult_u0.step5.add_sub4_u0.int_ip[5] ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.S[0] ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.S[1] ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.S[2] ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.S[3] ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.S[4] ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.S[5] ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.cg21 ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.cg43 ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.cg[0] ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.cg[1] ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.cg[2] ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.cg[3] ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.cg[4] ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.cp21 ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.cp43 ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.d1_0.a2._0_ ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.d1_0.a2.in0 ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.d1_0.a2.out ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.d1_0.g1 ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.d1_0.o2._0_ ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.d2_0.a2._0_ ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.d2_0.a2.out ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.d2_0.g1 ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.d2_0.o2._0_ ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.d3_0.a1._0_ ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.d3_0.a2._0_ ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.d3_0.a2.out ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.d3_0.g1 ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.d3_0.o2._0_ ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.d3_1.a2._0_ ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.d3_1.a2.out ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.d3_1.o2._0_ ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.d4_0.a2._0_ ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.d4_0.a2.in0 ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.d4_0.a2.out ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.d4_0.g1 ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.d4_0.o2._0_ ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.d5_0.a1._0_ ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.d5_0.a1.in0 ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.d5_0.a2._0_ ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.d5_0.a2.out ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.d5_0.g1 ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.d5_0.o2._0_ ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.d5_1.a2._0_ ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.d5_1.a2.out ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.d5_1.o2._0_ ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.p_0.a._0_ ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.p_0.o._0_ ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.p_1.a._0_ ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.p_1.o._0_ ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.p_2.a._0_ ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.p_2.o._0_ ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.p_3.a._0_ ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.p_3.o._0_ ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.p_4.a._0_ ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.p_4.o._0_ ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.s0.temp ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.s0.xor2_0._0_ ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.s0.xor2_1._0_ ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.s1.temp ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.s1.xor2_0._0_ ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.s1.xor2_1._0_ ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.s2.temp ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.s2.xor2_0._0_ ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.s2.xor2_1._0_ ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.s3.temp ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.s3.xor2_0._0_ ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.s3.xor2_1._0_ ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.s4.temp ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.s4.xor2_0._0_ ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.s4.xor2_1._0_ ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.s5.temp ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.s5.xor2_0._0_ ;
 wire \mult_u0.step5.add_sub4_u0.ppa8_u0.s5.xor2_1._0_ ;
 wire \mult_u0.step5.add_sub4_u0.x0._0_ ;
 wire \mult_u0.step5.add_sub4_u0.x1._0_ ;
 wire \mult_u0.step5.add_sub4_u0.x2._0_ ;
 wire \mult_u0.step5.add_sub4_u0.x3._0_ ;
 wire \mult_u0.step5.add_sub4_u0.x4._0_ ;
 wire \mult_u0.step5.add_sub4_u0.x5._0_ ;
 wire \mult_u0.step6._00_ ;
 wire \mult_u0.step6._01_ ;
 wire \mult_u0.step6._03_ ;
 wire \mult_u0.step6._04_ ;
 wire \mult_u0.step6._05_ ;
 wire \mult_u0.step6._06_ ;
 wire \mult_u0.step6._08_ ;
 wire \mult_u0.step6.add_sub4_u0.int_ip[0] ;
 wire \mult_u0.step6.add_sub4_u0.int_ip[1] ;
 wire \mult_u0.step6.add_sub4_u0.int_ip[2] ;
 wire \mult_u0.step6.add_sub4_u0.int_ip[3] ;
 wire \mult_u0.step6.add_sub4_u0.int_ip[4] ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.S[0] ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.S[1] ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.S[2] ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.S[3] ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.S[4] ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.cg21 ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.cg[0] ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.cg[1] ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.cg[2] ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.cg[3] ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.cp21 ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.d1_0.a2._0_ ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.d1_0.a2.in0 ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.d1_0.a2.out ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.d1_0.g1 ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.d1_0.o2._0_ ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.d2_0.a2._0_ ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.d2_0.a2.out ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.d2_0.g1 ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.d2_0.o2._0_ ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.d3_0.a1._0_ ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.d3_0.a2._0_ ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.d3_0.a2.out ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.d3_0.g1 ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.d3_0.o2._0_ ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.d3_1.a2._0_ ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.d3_1.a2.out ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.d3_1.o2._0_ ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.d4_0.a2._0_ ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.d4_0.a2.in0 ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.d4_0.a2.out ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.d4_0.g1 ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.d4_0.o2._0_ ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.p_0.a._0_ ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.p_0.o._0_ ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.p_1.a._0_ ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.p_1.o._0_ ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.p_2.a._0_ ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.p_2.o._0_ ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.p_3.a._0_ ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.p_3.o._0_ ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.s0.temp ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.s0.xor2_0._0_ ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.s0.xor2_1._0_ ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.s1.temp ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.s1.xor2_0._0_ ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.s1.xor2_1._0_ ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.s2.temp ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.s2.xor2_0._0_ ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.s2.xor2_1._0_ ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.s3.temp ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.s3.xor2_0._0_ ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.s3.xor2_1._0_ ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.s4.temp ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.s4.xor2_0._0_ ;
 wire \mult_u0.step6.add_sub4_u0.ppa8_u0.s4.xor2_1._0_ ;
 wire \mult_u0.step6.add_sub4_u0.x0._0_ ;
 wire \mult_u0.step6.add_sub4_u0.x1._0_ ;
 wire \mult_u0.step6.add_sub4_u0.x2._0_ ;
 wire \mult_u0.step6.add_sub4_u0.x3._0_ ;
 wire \mult_u0.step6.add_sub4_u0.x4._0_ ;
 wire \mult_u0.step7._00_ ;
 wire \mult_u0.step7._01_ ;
 wire \mult_u0.step7._03_ ;
 wire \mult_u0.step7._04_ ;
 wire \mult_u0.step7._05_ ;
 wire \mult_u0.step7._08_ ;
 wire \mult_u0.step7.add_sub4_u0.int_ip[0] ;
 wire \mult_u0.step7.add_sub4_u0.int_ip[1] ;
 wire \mult_u0.step7.add_sub4_u0.int_ip[2] ;
 wire \mult_u0.step7.add_sub4_u0.int_ip[3] ;
 wire \mult_u0.step7.add_sub4_u0.ppa8_u0.S[0] ;
 wire \mult_u0.step7.add_sub4_u0.ppa8_u0.S[1] ;
 wire \mult_u0.step7.add_sub4_u0.ppa8_u0.S[2] ;
 wire \mult_u0.step7.add_sub4_u0.ppa8_u0.S[3] ;
 wire \mult_u0.step7.add_sub4_u0.ppa8_u0.cg21 ;
 wire \mult_u0.step7.add_sub4_u0.ppa8_u0.cg[0] ;
 wire \mult_u0.step7.add_sub4_u0.ppa8_u0.cg[1] ;
 wire \mult_u0.step7.add_sub4_u0.ppa8_u0.cg[2] ;
 wire \mult_u0.step7.add_sub4_u0.ppa8_u0.cp21 ;
 wire \mult_u0.step7.add_sub4_u0.ppa8_u0.d1_0.a2._0_ ;
 wire \mult_u0.step7.add_sub4_u0.ppa8_u0.d1_0.a2.in0 ;
 wire \mult_u0.step7.add_sub4_u0.ppa8_u0.d1_0.a2.out ;
 wire \mult_u0.step7.add_sub4_u0.ppa8_u0.d1_0.g1 ;
 wire \mult_u0.step7.add_sub4_u0.ppa8_u0.d1_0.o2._0_ ;
 wire \mult_u0.step7.add_sub4_u0.ppa8_u0.d2_0.a2._0_ ;
 wire \mult_u0.step7.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ;
 wire \mult_u0.step7.add_sub4_u0.ppa8_u0.d2_0.a2.out ;
 wire \mult_u0.step7.add_sub4_u0.ppa8_u0.d2_0.g1 ;
 wire \mult_u0.step7.add_sub4_u0.ppa8_u0.d2_0.o2._0_ ;
 wire \mult_u0.step7.add_sub4_u0.ppa8_u0.d3_0.a1._0_ ;
 wire \mult_u0.step7.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ;
 wire \mult_u0.step7.add_sub4_u0.ppa8_u0.d3_0.a2._0_ ;
 wire \mult_u0.step7.add_sub4_u0.ppa8_u0.d3_0.a2.out ;
 wire \mult_u0.step7.add_sub4_u0.ppa8_u0.d3_0.g1 ;
 wire \mult_u0.step7.add_sub4_u0.ppa8_u0.d3_0.o2._0_ ;
 wire \mult_u0.step7.add_sub4_u0.ppa8_u0.d3_1.a2._0_ ;
 wire \mult_u0.step7.add_sub4_u0.ppa8_u0.d3_1.a2.out ;
 wire \mult_u0.step7.add_sub4_u0.ppa8_u0.d3_1.o2._0_ ;
 wire \mult_u0.step7.add_sub4_u0.ppa8_u0.p_0.a._0_ ;
 wire \mult_u0.step7.add_sub4_u0.ppa8_u0.p_0.o._0_ ;
 wire \mult_u0.step7.add_sub4_u0.ppa8_u0.p_1.a._0_ ;
 wire \mult_u0.step7.add_sub4_u0.ppa8_u0.p_1.o._0_ ;
 wire \mult_u0.step7.add_sub4_u0.ppa8_u0.p_2.a._0_ ;
 wire \mult_u0.step7.add_sub4_u0.ppa8_u0.p_2.o._0_ ;
 wire \mult_u0.step7.add_sub4_u0.ppa8_u0.s0.temp ;
 wire \mult_u0.step7.add_sub4_u0.ppa8_u0.s0.xor2_0._0_ ;
 wire \mult_u0.step7.add_sub4_u0.ppa8_u0.s0.xor2_1._0_ ;
 wire \mult_u0.step7.add_sub4_u0.ppa8_u0.s1.temp ;
 wire \mult_u0.step7.add_sub4_u0.ppa8_u0.s1.xor2_0._0_ ;
 wire \mult_u0.step7.add_sub4_u0.ppa8_u0.s1.xor2_1._0_ ;
 wire \mult_u0.step7.add_sub4_u0.ppa8_u0.s2.temp ;
 wire \mult_u0.step7.add_sub4_u0.ppa8_u0.s2.xor2_0._0_ ;
 wire \mult_u0.step7.add_sub4_u0.ppa8_u0.s2.xor2_1._0_ ;
 wire \mult_u0.step7.add_sub4_u0.ppa8_u0.s3.temp ;
 wire \mult_u0.step7.add_sub4_u0.ppa8_u0.s3.xor2_0._0_ ;
 wire \mult_u0.step7.add_sub4_u0.ppa8_u0.s3.xor2_1._0_ ;
 wire \mult_u0.step7.add_sub4_u0.x0._0_ ;
 wire \mult_u0.step7.add_sub4_u0.x1._0_ ;
 wire \mult_u0.step7.add_sub4_u0.x2._0_ ;
 wire \mult_u0.step7.add_sub4_u0.x3._0_ ;
 wire \mult_u0.step7.next_acc[0] ;
 wire \mult_u0.step7.next_acc[1] ;
 wire \mult_u0.step7.next_acc[2] ;
 wire \mult_u0.x_sign._0_ ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \out[0] ;
 wire \out[1] ;
 wire \out[2] ;
 wire \out[3] ;
 wire \out[4] ;
 wire \out[5] ;
 wire \out[6] ;
 wire \out[7] ;
 wire \sel[0] ;
 wire \sel[1] ;
 wire \sel_d0[0] ;
 wire \sel_d0[1] ;
 wire \sel_d1[0] ;
 wire \sel_d1[1] ;
 wire \sel_d2[0] ;
 wire \sel_d2[1] ;
 wire \sel_d3[0] ;
 wire \sel_d3[1] ;
 wire \sel_d4[0] ;
 wire \sel_d4[1] ;
 wire \sel_d5[0] ;
 wire \sel_d5[1] ;
 wire \sel_d6[0] ;
 wire \sel_d6[1] ;
 wire \sel_d7[0] ;
 wire \sel_d7[1] ;
 wire \sel_d8[0] ;
 wire \sel_d8[1] ;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__174__I (.I(net62),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__175__I (.I(_043_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__190__A2 (.I(_052_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__190__A3 (.I(_055_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__192__A1 (.I(_044_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__192__A2 (.I(_045_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__192__A3 (.I(_060_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__202__A1 (.I(_067_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__204__A2 (.I(_067_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__204__B (.I(_044_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__205__A1 (.I(_070_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__207__A1 (.I(_067_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__209__A2 (.I(_067_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__209__B (.I(_044_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__210__A1 (.I(_074_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__212__A1 (.I(_067_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__214__A1 (.I(\out[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__214__A2 (.I(_067_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__214__B (.I(_044_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__217__A1 (.I(_067_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__219__A2 (.I(_067_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__219__B (.I(_044_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__222__A1 (.I(_067_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__224__A2 (.I(_067_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__224__B (.I(_044_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__227__A1 (.I(_067_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__229__A2 (.I(_067_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__229__B (.I(_044_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__230__A1 (.I(_090_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__232__A1 (.I(_067_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__234__A2 (.I(_067_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__234__B (.I(_044_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__237__A1 (.I(_067_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__239__A2 (.I(_067_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__239__B (.I(_044_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__240__A1 (.I(_098_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__242__A1 (.I(_045_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__242__A2 (.I(_060_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__245__I (.I(_045_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__246__I (.I(_060_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__247__A1 (.I(_104_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__247__A2 (.I(_105_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__247__B (.I(\add_u0.a[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__248__I (.I(_043_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__249__A2 (.I(_103_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__249__C (.I(_107_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__251__A1 (.I(_104_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__251__A2 (.I(_105_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__251__B (.I(\add_u0.a[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__252__A2 (.I(_103_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__252__C (.I(_107_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__254__A1 (.I(_104_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__254__A2 (.I(_105_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__254__B (.I(\add_u0.a[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__255__A2 (.I(_103_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__255__C (.I(_107_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__257__A1 (.I(_104_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__257__A2 (.I(_105_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__258__A2 (.I(_103_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__258__C (.I(_107_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__260__A1 (.I(_104_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__260__A2 (.I(_105_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__260__B (.I(\add_u0.a[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__261__A2 (.I(_103_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__261__C (.I(_107_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__263__A1 (.I(_104_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__263__A2 (.I(_105_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__263__B (.I(\add_u0.a[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__264__A2 (.I(_103_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__264__C (.I(_107_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__266__A1 (.I(_104_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__266__A2 (.I(_105_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__266__B (.I(\add_u0.a[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__267__A2 (.I(_103_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__267__C (.I(_107_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__269__A1 (.I(_104_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__269__A2 (.I(_105_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__270__A2 (.I(_103_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__270__C (.I(_107_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__272__A1 (.I(_104_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__272__A2 (.I(_105_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__272__B (.I(\add_u0.b[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__273__A2 (.I(_103_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__273__C (.I(_107_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__275__A1 (.I(_104_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__275__A2 (.I(_105_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__275__B (.I(\add_u0.b[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__276__A2 (.I(_103_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__276__C (.I(_107_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__278__A1 (.I(_104_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__278__A2 (.I(_105_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__278__B (.I(\add_u0.b[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__279__A2 (.I(_103_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__279__C (.I(_107_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__281__A1 (.I(_104_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__281__A2 (.I(_060_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__281__B (.I(\add_u0.b[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__282__A2 (.I(_103_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__282__C (.I(_107_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__284__A1 (.I(_104_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__284__A2 (.I(_060_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__284__B (.I(\add_u0.b[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__285__A2 (.I(_103_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__285__C (.I(_043_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__287__A1 (.I(_104_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__287__A2 (.I(_060_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__287__B (.I(\add_u0.b[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__288__A2 (.I(_103_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__288__C (.I(_043_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__290__A1 (.I(_104_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__290__A2 (.I(_060_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__290__B (.I(\add_u0.b[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__291__A2 (.I(_103_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__291__C (.I(_043_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__293__A1 (.I(_104_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__293__A2 (.I(_060_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__293__B (.I(\add_u0.b[7] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__294__A2 (.I(_103_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__294__C (.I(_043_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__296__A1 (.I(_104_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__296__A2 (.I(_060_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__297__A2 (.I(_103_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__297__C (.I(_043_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__299__A1 (.I(_104_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__299__A2 (.I(_060_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__300__A2 (.I(_103_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__300__C (.I(_043_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__302__A1 (.I(_104_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__302__A2 (.I(_060_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__303__A2 (.I(_103_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__303__C (.I(_043_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__305__A1 (.I(_104_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__305__A2 (.I(_060_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__306__A2 (.I(_103_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__306__C (.I(_043_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__308__A1 (.I(_045_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__308__A2 (.I(_060_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__309__C (.I(_043_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__311__A1 (.I(_045_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__311__A2 (.I(_060_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__312__C (.I(_043_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__314__A1 (.I(_045_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__314__A2 (.I(_060_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__315__C (.I(_043_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__317__A1 (.I(_045_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__317__A2 (.I(_060_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__317__B (.I(\mult_add_u0.m[7] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__318__C (.I(_043_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__319__A2 (.I(_044_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__319__A3 (.I(_105_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__323__A2 (.I(_156_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__325__A2 (.I(_105_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__325__A3 (.I(_158_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__326__B (.I(_107_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__327__A2 (.I(_156_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__328__A2 (.I(_105_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__328__A3 (.I(_158_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__329__B (.I(_107_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__330__A2 (.I(_156_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__331__A1 (.I(\out[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__331__A2 (.I(_105_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__331__A3 (.I(_158_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__332__B (.I(_107_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__333__A2 (.I(_156_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__334__A2 (.I(_105_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__334__A3 (.I(_158_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__335__B (.I(_107_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__336__A2 (.I(_156_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__337__A2 (.I(_105_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__337__A3 (.I(_158_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__338__B (.I(_107_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__339__A2 (.I(_156_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__340__A2 (.I(_105_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__340__A3 (.I(_158_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__341__B (.I(_107_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__342__A2 (.I(_156_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__343__A2 (.I(_105_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__343__A3 (.I(_158_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__344__B (.I(_107_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__345__A2 (.I(_156_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__346__A2 (.I(_105_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__346__A3 (.I(_158_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__347__B (.I(_107_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__368__D (.I(\sel_d4[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__371__D (.I(\sel_d5[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__476__CLK (.I(clknet_3_2__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._053__A1  (.I(\add_u0.b[7] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._055__I  (.I(\add_u0.b[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._056__I  (.I(\add_u0.b[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._057__A2  (.I(\add_u0.a[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._057__B2  (.I(\add_u0.a[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._059__I  (.I(\add_u0.a[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._060__A1  (.I(\add_u0.b[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._060__B1  (.I(\add_u0.b[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._061__I  (.I(\add_u0.b[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._062__A1  (.I(\add_u0.a[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._063__I  (.I(\add_u0.a[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._064__A1  (.I(\add_u0.b[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._065__I  (.I(\add_u0.a[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._066__A1  (.I(\add_u0.b[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._066__B1  (.I(\add_u0.b[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._067__A1  (.I(\add_u0.b[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._069__I  (.I(\add_u0.a[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._070__A1  (.I(\add_u0.a[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._070__A2  (.I(\add_u0.b[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._072__A1  (.I(\add_u0.a[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._072__A2  (.I(\add_u0.b[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._073__A1  (.I(\add_u0.b[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._074__I  (.I(\add_u0.b[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._075__A2  (.I(\add_u0.a[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._076__I  (.I(\add_u0.a[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._077__I  (.I(\add_u0.b[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._078__A1  (.I(\add_u0.b[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._078__B1  (.I(\add_u0.b[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._078__C2  (.I(\add_u0.a[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._081__I  (.I(\add_u0.b[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._082__A2  (.I(\add_u0.a[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._085__A1  (.I(\add_u0.a[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._088__I0  (.I(\add_u0.a[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._088__I1  (.I(\add_u0.b[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._088__S  (.I(\add_u0._033_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._089__A1  (.I(\add_u0.c_in ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._091__I0  (.I(\add_u0.a[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._091__I1  (.I(\add_u0.b[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._091__S  (.I(\add_u0._033_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._092__A1  (.I(\add_u0.c_in ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._094__I0  (.I(\add_u0.a[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._094__I1  (.I(\add_u0.b[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._094__S  (.I(\add_u0._033_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._095__A1  (.I(\add_u0.c_in ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._097__I1  (.I(\add_u0.b[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._097__S  (.I(\add_u0._033_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._098__A1  (.I(\add_u0.c_in ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._100__I0  (.I(\add_u0.a[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._100__I1  (.I(\add_u0.b[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._100__S  (.I(\add_u0._033_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._101__A1  (.I(\add_u0.c_in ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._103__I0  (.I(\add_u0.a[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._103__I1  (.I(\add_u0.b[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._103__S  (.I(\add_u0._033_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._104__A1  (.I(\add_u0.c_in ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._106__A1  (.I(\add_u0.c_in ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._108__I0  (.I(\add_u0.b[7] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._108__S  (.I(\add_u0._033_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._110__A1  (.I(\add_u0.a[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._110__A2  (.I(\add_u0._033_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._111__A2  (.I(\add_u0._033_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._112__A1  (.I(\add_u0.a[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._112__A2  (.I(\add_u0._033_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._113__A2  (.I(\add_u0._033_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._114__A1  (.I(\add_u0.b[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._114__A2  (.I(\add_u0._033_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._115__A2  (.I(\add_u0._033_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._116__A2  (.I(\add_u0._033_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._117__A2  (.I(\add_u0._033_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._118__A1  (.I(\add_u0.a[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._118__A2  (.I(\add_u0._033_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._119__A2  (.I(\add_u0._033_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._120__A1  (.I(\add_u0.a[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._120__A2  (.I(\add_u0._033_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0._121__A2  (.I(\add_u0._033_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0.ppa_u0.d1_0.a2._1__A1  (.I(\add_u0.c_in ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_add_u0.ppa_u0.s0.xor2_1._1__A2  (.I(\add_u0.c_in ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_clk_I (.I(net114),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_0__f_clk_I (.I(clknet_0_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_1__f_clk_I (.I(clknet_0_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_2__f_clk_I (.I(clknet_0_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_3__f_clk_I (.I(clknet_0_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_4__f_clk_I (.I(clknet_0_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_5__f_clk_I (.I(clknet_0_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_6__f_clk_I (.I(clknet_0_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_7__f_clk_I (.I(clknet_0_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_0_clk_I (.I(clknet_3_0__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_10_clk_I (.I(clknet_3_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_11_clk_I (.I(clknet_3_3__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_12_clk_I (.I(clknet_3_3__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_13_clk_I (.I(clknet_3_3__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_14_clk_I (.I(clknet_3_3__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_15_clk_I (.I(clknet_3_3__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_16_clk_I (.I(clknet_3_2__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_17_clk_I (.I(clknet_3_2__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_18_clk_I (.I(clknet_3_2__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_1_clk_I (.I(clknet_3_0__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_20_clk_I (.I(clknet_3_2__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_21_clk_I (.I(clknet_3_2__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_22_clk_I (.I(clknet_3_2__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_23_clk_I (.I(clknet_3_2__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_24_clk_I (.I(clknet_3_2__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_25_clk_I (.I(clknet_3_2__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_26_clk_I (.I(clknet_3_2__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_27_clk_I (.I(clknet_3_3__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_28_clk_I (.I(clknet_3_3__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_29_clk_I (.I(clknet_3_3__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_2_clk_I (.I(clknet_3_0__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_30_clk_I (.I(clknet_3_3__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_31_clk_I (.I(clknet_3_3__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_32_clk_I (.I(clknet_3_3__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_33_clk_I (.I(clknet_3_3__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_34_clk_I (.I(clknet_3_3__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_35_clk_I (.I(clknet_3_6__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_36_clk_I (.I(clknet_3_6__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_37_clk_I (.I(clknet_3_6__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_38_clk_I (.I(clknet_3_6__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_39_clk_I (.I(clknet_3_6__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_3_clk_I (.I(clknet_3_0__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_40_clk_I (.I(clknet_3_6__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_41_clk_I (.I(clknet_3_6__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_42_clk_I (.I(clknet_3_6__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_44_clk_I (.I(clknet_3_7__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_45_clk_I (.I(clknet_3_7__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_46_clk_I (.I(clknet_3_7__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_48_clk_I (.I(clknet_3_7__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_49_clk_I (.I(clknet_3_7__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_4_clk_I (.I(clknet_3_2__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_50_clk_I (.I(clknet_3_6__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_51_clk_I (.I(clknet_3_7__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_53_clk_I (.I(clknet_3_4__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_54_clk_I (.I(clknet_3_5__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_55_clk_I (.I(clknet_3_4__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_56_clk_I (.I(clknet_3_5__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_57_clk_I (.I(clknet_3_7__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_58_clk_I (.I(clknet_3_5__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_59_clk_I (.I(clknet_3_5__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_5_clk_I (.I(clknet_3_0__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_60_clk_I (.I(clknet_3_5__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_61_clk_I (.I(clknet_3_5__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_62_clk_I (.I(clknet_3_5__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_63_clk_I (.I(clknet_3_5__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_64_clk_I (.I(clknet_3_5__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_65_clk_I (.I(clknet_3_5__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_66_clk_I (.I(clknet_3_5__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_67_clk_I (.I(clknet_3_5__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_68_clk_I (.I(clknet_3_5__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_69_clk_I (.I(clknet_3_4__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_6_clk_I (.I(clknet_3_2__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_70_clk_I (.I(clknet_3_4__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_71_clk_I (.I(clknet_3_4__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_72_clk_I (.I(clknet_3_4__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_73_clk_I (.I(clknet_3_4__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_75_clk_I (.I(clknet_3_4__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_76_clk_I (.I(clknet_3_4__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_77_clk_I (.I(clknet_3_4__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_78_clk_I (.I(clknet_3_4__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_79_clk_I (.I(clknet_3_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_7_clk_I (.I(clknet_3_0__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_80_clk_I (.I(clknet_3_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_81_clk_I (.I(clknet_3_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_82_clk_I (.I(clknet_3_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_83_clk_I (.I(clknet_3_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_84_clk_I (.I(clknet_3_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_86_clk_I (.I(clknet_3_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_87_clk_I (.I(clknet_3_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_88_clk_I (.I(clknet_3_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_89_clk_I (.I(clknet_3_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_8_clk_I (.I(clknet_3_0__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_90_clk_I (.I(clknet_3_0__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_91_clk_I (.I(clknet_3_0__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_92_clk_I (.I(clknet_3_0__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_93_clk_I (.I(clknet_3_0__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_94_clk_I (.I(clknet_3_0__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_95_clk_I (.I(clknet_3_0__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_96_clk_I (.I(clknet_3_0__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_9_clk_I (.I(clknet_3_0__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(i_wb_addr[18]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(i_wb_addr[19]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(i_wb_addr[1]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(i_wb_addr[20]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(i_wb_addr[21]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(i_wb_addr[22]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(i_wb_addr[23]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(i_wb_addr[24]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(i_wb_addr[25]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(i_wb_addr[26]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(i_wb_addr[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(i_wb_addr[27]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(i_wb_addr[28]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(i_wb_addr[29]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(i_wb_addr[2]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(i_wb_addr[30]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(i_wb_addr[31]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(i_wb_addr[3]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(i_wb_addr[4]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(i_wb_addr[5]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(i_wb_addr[6]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(i_wb_addr[10]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(i_wb_addr[7]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(i_wb_addr[8]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(i_wb_addr[9]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(i_wb_cyc),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input34_I (.I(i_wb_data[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input35_I (.I(i_wb_data[10]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input36_I (.I(i_wb_data[11]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input37_I (.I(i_wb_data[12]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input38_I (.I(i_wb_data[13]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input39_I (.I(i_wb_data[14]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(i_wb_addr[11]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input40_I (.I(i_wb_data[15]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input41_I (.I(i_wb_data[16]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input42_I (.I(i_wb_data[17]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input43_I (.I(i_wb_data[18]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input44_I (.I(i_wb_data[19]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input45_I (.I(i_wb_data[1]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input46_I (.I(i_wb_data[20]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input47_I (.I(i_wb_data[21]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input48_I (.I(i_wb_data[22]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input49_I (.I(i_wb_data[23]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(i_wb_addr[12]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input50_I (.I(i_wb_data[24]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input51_I (.I(i_wb_data[25]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input52_I (.I(i_wb_data[2]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input53_I (.I(i_wb_data[3]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input54_I (.I(i_wb_data[4]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input55_I (.I(i_wb_data[5]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input56_I (.I(i_wb_data[6]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input57_I (.I(i_wb_data[7]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input58_I (.I(i_wb_data[8]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input59_I (.I(i_wb_data[9]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(i_wb_addr[13]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input60_I (.I(i_wb_stb),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input61_I (.I(i_wb_we),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input62_I (.I(reset),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(i_wb_addr[14]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(i_wb_addr[15]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(i_wb_addr[16]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(i_wb_addr[17]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0._018__I  (.I(net62),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0._034__D  (.I(\add_u0.b[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0._035__D  (.I(\add_u0.b[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0._036__D  (.I(\add_u0.b[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0._037__D  (.I(\add_u0.b[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0._038__D  (.I(\add_u0.b[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0._039__D  (.I(\add_u0.b[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0._040__D  (.I(\add_u0.b[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0._041__D  (.I(\add_u0.b[7] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0._073__CLK  (.I(clknet_3_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0._093__CLK  (.I(clknet_3_6__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.add0._056__I  (.I(\mult_add_u0.add0.b[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.add0._078__A1  (.I(\mult_add_u0.add0.b[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.add0._088__S  (.I(\mult_add_u0.add0._033_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.add0._091__S  (.I(\mult_add_u0.add0._033_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.add0._094__S  (.I(\mult_add_u0.add0._033_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.add0._097__S  (.I(\mult_add_u0.add0._033_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.add0._100__I1  (.I(\mult_add_u0.add0.b[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.add0._100__S  (.I(\mult_add_u0.add0._033_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.add0._103__S  (.I(\mult_add_u0.add0._033_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.add0._108__S  (.I(\mult_add_u0.add0._033_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.add0._110__A2  (.I(\mult_add_u0.add0._033_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.add0._111__A2  (.I(\mult_add_u0.add0._033_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.add0._112__A2  (.I(\mult_add_u0.add0._033_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.add0._113__A2  (.I(\mult_add_u0.add0._033_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.add0._114__A2  (.I(\mult_add_u0.add0._033_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.add0._115__A2  (.I(\mult_add_u0.add0._033_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.add0._116__A2  (.I(\mult_add_u0.add0._033_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.add0._117__A2  (.I(\mult_add_u0.add0._033_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.add0._118__A2  (.I(\mult_add_u0.add0._033_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.add0._119__A2  (.I(\mult_add_u0.add0._033_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.add0._120__A2  (.I(\mult_add_u0.add0._033_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.add0._121__A2  (.I(\mult_add_u0.add0._033_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0._026__I  (.I(net62),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0._027__A2  (.I(\mult_add_u0.mult0._009_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0._029__A1  (.I(\mult_add_u0.mult0._009_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0._031__A1  (.I(\mult_add_u0.mult0._009_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0._033__A1  (.I(\mult_add_u0.mult0._009_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0._035__A1  (.I(\mult_add_u0.mult0._009_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0._037__A1  (.I(\mult_add_u0.mult0._009_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0._039__A1  (.I(\mult_add_u0.mult0._009_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0._041__A1  (.I(\mult_add_u0.mult0._009_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0._053__CLK  (.I(clknet_3_4__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0._100__D  (.I(\mult_add_u0.mult0.Q[3][1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0._108__CLK  (.I(clknet_3_7__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0._122__CLK  (.I(clknet_3_7__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0._141__D  (.I(\mult_add_u0.mult0.multiplicand[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0._142__D  (.I(\mult_add_u0.mult0.multiplicand[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0._143__D  (.I(\mult_add_u0.mult0.multiplicand[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0._144__D  (.I(\mult_add_u0.mult0.multiplicand[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0._145__D  (.I(\mult_add_u0.mult0.multiplicand[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0._146__D  (.I(\mult_add_u0.mult0.multiplicand[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0._163__D  (.I(\mult_add_u0.mult0.multiplicand_s3[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0._182__D  (.I(\add_u0.a[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0._183__D  (.I(\add_u0.a[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0._184__D  (.I(\add_u0.a[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0._186__D  (.I(\add_u0.a[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0._187__D  (.I(\add_u0.a[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0._188__D  (.I(\add_u0.a[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step1._09__A2  (.I(\mult_add_u0.mult0.multiplier[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step1._11__S  (.I(\mult_add_u0.mult0.step1._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step1._13__S  (.I(\mult_add_u0.mult0.step1._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step1._15__S  (.I(\mult_add_u0.mult0.step1._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step1._17__S  (.I(\mult_add_u0.mult0.step1._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step1._19__S  (.I(\mult_add_u0.mult0.step1._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step1._21__S  (.I(\mult_add_u0.mult0.step1._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step1._32__I  (.I(\mult_add_u0.mult0.multiplier[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d1_0.a2._1__A1  (.I(\mult_add_u0.mult0.multiplier[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step1.add_sub4_u0.x0._1__A1  (.I(\mult_add_u0.mult0.multiplier[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step1.add_sub4_u0.x1._1__A1  (.I(\mult_add_u0.mult0.multiplier[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step1.add_sub4_u0.x1._1__A2  (.I(\mult_add_u0.mult0.multiplicand[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step1.add_sub4_u0.x2._1__A1  (.I(\mult_add_u0.mult0.multiplier[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step1.add_sub4_u0.x2._1__A2  (.I(\mult_add_u0.mult0.multiplicand[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step1.add_sub4_u0.x3._1__A1  (.I(\mult_add_u0.mult0.multiplier[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step1.add_sub4_u0.x3._1__A2  (.I(\mult_add_u0.mult0.multiplicand[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step1.add_sub4_u0.x4._1__A1  (.I(\mult_add_u0.mult0.multiplier[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step1.add_sub4_u0.x4._1__A2  (.I(\mult_add_u0.mult0.multiplicand[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step1.add_sub4_u0.x5._1__A1  (.I(\mult_add_u0.mult0.multiplier[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step1.add_sub4_u0.x5._1__A2  (.I(\mult_add_u0.mult0.multiplicand[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step1.add_sub4_u0.x6._1__A1  (.I(\mult_add_u0.mult0.multiplier[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step1.add_sub4_u0.x6._1__A2  (.I(\mult_add_u0.mult0.multiplicand[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step2._09__A2  (.I(\mult_add_u0.mult0.Q_s1[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step2._11__S  (.I(\mult_add_u0.mult0.step2._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step2._13__S  (.I(\mult_add_u0.mult0.step2._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step2._15__S  (.I(\mult_add_u0.mult0.step2._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step2._17__S  (.I(\mult_add_u0.mult0.step2._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step2._19__S  (.I(\mult_add_u0.mult0.step2._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step2._21__S  (.I(\mult_add_u0.mult0.step2._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step2._32__I  (.I(\mult_add_u0.mult0.Q_s1[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d1_0.a2._1__A1  (.I(\mult_add_u0.mult0.Q_s1[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step2.add_sub4_u0.x0._1__A1  (.I(\mult_add_u0.mult0.Q_s1[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step2.add_sub4_u0.x1._1__A1  (.I(\mult_add_u0.mult0.Q_s1[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step2.add_sub4_u0.x2._1__A1  (.I(\mult_add_u0.mult0.Q_s1[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step2.add_sub4_u0.x3._1__A1  (.I(\mult_add_u0.mult0.Q_s1[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step2.add_sub4_u0.x4._1__A1  (.I(\mult_add_u0.mult0.Q_s1[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step2.add_sub4_u0.x5._1__A1  (.I(\mult_add_u0.mult0.Q_s1[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step2.add_sub4_u0.x6._1__A1  (.I(\mult_add_u0.mult0.Q_s1[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step3._09__A2  (.I(\mult_add_u0.mult0.Q_s2[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step3._11__S  (.I(\mult_add_u0.mult0.step3._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step3._13__S  (.I(\mult_add_u0.mult0.step3._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step3._15__S  (.I(\mult_add_u0.mult0.step3._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step3._17__S  (.I(\mult_add_u0.mult0.step3._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step3._19__S  (.I(\mult_add_u0.mult0.step3._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step3._21__S  (.I(\mult_add_u0.mult0.step3._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step3._32__I  (.I(\mult_add_u0.mult0.Q_s2[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d1_0.a2._1__A1  (.I(\mult_add_u0.mult0.Q_s2[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step3.add_sub4_u0.x0._1__A1  (.I(\mult_add_u0.mult0.Q_s2[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step3.add_sub4_u0.x1._1__A1  (.I(\mult_add_u0.mult0.Q_s2[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step3.add_sub4_u0.x2._1__A1  (.I(\mult_add_u0.mult0.Q_s2[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step3.add_sub4_u0.x3._1__A1  (.I(\mult_add_u0.mult0.Q_s2[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step3.add_sub4_u0.x4._1__A1  (.I(\mult_add_u0.mult0.Q_s2[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step3.add_sub4_u0.x5._1__A1  (.I(\mult_add_u0.mult0.Q_s2[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step3.add_sub4_u0.x6._1__A1  (.I(\mult_add_u0.mult0.Q_s2[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step4._09__A2  (.I(\mult_add_u0.mult0.Q_s3[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step4._11__S  (.I(\mult_add_u0.mult0.step4._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step4._13__S  (.I(\mult_add_u0.mult0.step4._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step4._15__S  (.I(\mult_add_u0.mult0.step4._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step4._17__S  (.I(\mult_add_u0.mult0.step4._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step4._19__S  (.I(\mult_add_u0.mult0.step4._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step4._21__S  (.I(\mult_add_u0.mult0.step4._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step4._23__S  (.I(\mult_add_u0.mult0.step4._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step4._32__I  (.I(\mult_add_u0.mult0.Q_s3[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d1_0.a2._1__A1  (.I(\mult_add_u0.mult0.Q_s3[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s0.xor2_1._1__A2  (.I(\mult_add_u0.mult0.Q_s3[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step4.add_sub4_u0.x0._1__A1  (.I(\mult_add_u0.mult0.Q_s3[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step4.add_sub4_u0.x1._1__A1  (.I(\mult_add_u0.mult0.Q_s3[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step4.add_sub4_u0.x2._1__A1  (.I(\mult_add_u0.mult0.Q_s3[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step4.add_sub4_u0.x2._1__A2  (.I(\mult_add_u0.mult0.multiplicand_s3[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step4.add_sub4_u0.x3._1__A1  (.I(\mult_add_u0.mult0.Q_s3[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step4.add_sub4_u0.x4._1__A1  (.I(\mult_add_u0.mult0.Q_s3[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step4.add_sub4_u0.x5._1__A1  (.I(\mult_add_u0.mult0.Q_s3[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step4.add_sub4_u0.x6._1__A1  (.I(\mult_add_u0.mult0.Q_s3[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step5._09__A2  (.I(\mult_add_u0.mult0.Q_s4[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step5._13__S  (.I(\mult_add_u0.mult0.step5._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step5._15__S  (.I(\mult_add_u0.mult0.step5._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step5._17__S  (.I(\mult_add_u0.mult0.step5._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step5._19__S  (.I(\mult_add_u0.mult0.step5._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step5._21__S  (.I(\mult_add_u0.mult0.step5._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step5._23__S  (.I(\mult_add_u0.mult0.step5._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step5._26__I  (.I(\mult_add_u0.mult0.Q_s4[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step5._32__I  (.I(\mult_add_u0.mult0.Q_s4[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d1_0.a2._1__A1  (.I(\mult_add_u0.mult0.Q_s4[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s0.xor2_1._1__A2  (.I(\mult_add_u0.mult0.Q_s4[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step5.add_sub4_u0.x0._1__A1  (.I(\mult_add_u0.mult0.Q_s4[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step5.add_sub4_u0.x1._1__A1  (.I(\mult_add_u0.mult0.Q_s4[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step5.add_sub4_u0.x2._1__A1  (.I(\mult_add_u0.mult0.Q_s4[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step5.add_sub4_u0.x3._1__A1  (.I(\mult_add_u0.mult0.Q_s4[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step5.add_sub4_u0.x4._1__A1  (.I(\mult_add_u0.mult0.Q_s4[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step5.add_sub4_u0.x5._1__A1  (.I(\mult_add_u0.mult0.Q_s4[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step6._09__A2  (.I(\mult_add_u0.mult0.Q_s5[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step6._13__S  (.I(\mult_add_u0.mult0.step6._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step6._15__S  (.I(\mult_add_u0.mult0.step6._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step6._17__S  (.I(\mult_add_u0.mult0.step6._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step6._19__S  (.I(\mult_add_u0.mult0.step6._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step6._23__S  (.I(\mult_add_u0.mult0.step6._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step6._32__I  (.I(\mult_add_u0.mult0.Q_s5[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d1_0.a2._1__A1  (.I(\mult_add_u0.mult0.Q_s5[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s0.xor2_1._1__A2  (.I(\mult_add_u0.mult0.Q_s5[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step6.add_sub4_u0.x0._1__A1  (.I(\mult_add_u0.mult0.Q_s5[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step6.add_sub4_u0.x1._1__A1  (.I(\mult_add_u0.mult0.Q_s5[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step6.add_sub4_u0.x2._1__A1  (.I(\mult_add_u0.mult0.Q_s5[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step6.add_sub4_u0.x3._1__A1  (.I(\mult_add_u0.mult0.Q_s5[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step6.add_sub4_u0.x4._1__A1  (.I(\mult_add_u0.mult0.Q_s5[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step7._09__A2  (.I(\mult_add_u0.mult0.Q_s6[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d1_0.a2._1__A1  (.I(\mult_add_u0.mult0.Q_s6[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s0.xor2_1._1__A2  (.I(\mult_add_u0.mult0.Q_s6[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step7.add_sub4_u0.x0._1__A1  (.I(\mult_add_u0.mult0.Q_s6[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step7.add_sub4_u0.x1._1__A1  (.I(\mult_add_u0.mult0.Q_s6[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step7.add_sub4_u0.x2._1__A1  (.I(\mult_add_u0.mult0.Q_s6[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.step7.add_sub4_u0.x3._1__A1  (.I(\mult_add_u0.mult0.Q_s6[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_add_u0.mult0.x_sign._1__A2  (.I(\mult_add_u0.m[7] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0._026__I  (.I(net62),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0._027__A2  (.I(\mult_u0._009_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0._029__A1  (.I(\mult_u0._009_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0._031__A1  (.I(\mult_u0._009_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0._033__A1  (.I(\mult_u0._009_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0._034__I  (.I(\mult_u0.step7.next_acc[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0._035__A1  (.I(\mult_u0._009_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0._036__I  (.I(\mult_u0.step7.next_acc[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0._037__A1  (.I(\mult_u0._009_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0._038__I  (.I(\mult_u0.step7.next_acc[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0._039__A1  (.I(\mult_u0._009_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0._041__A1  (.I(\mult_u0._009_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0._073__D  (.I(\mult_u0.Q[1][2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0._143__D  (.I(\mult_u0.multiplicand[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0._146__D  (.I(\mult_u0.multiplicand[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0._182__D  (.I(\add_u0.b[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0._183__D  (.I(\add_u0.b[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0._184__D  (.I(\add_u0.b[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0._185__D  (.I(\add_u0.b[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0._186__D  (.I(\add_u0.b[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0._187__D  (.I(\add_u0.b[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0._188__D  (.I(\add_u0.b[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0._189__D  (.I(\add_u0.a[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0._190__D  (.I(\add_u0.a[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0._191__D  (.I(\add_u0.a[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0._193__D  (.I(\add_u0.a[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0._194__D  (.I(\add_u0.a[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0._195__D  (.I(\add_u0.a[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step1._09__A2  (.I(\mult_u0.multiplier[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step1._11__S  (.I(\mult_u0.step1._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step1._13__S  (.I(\mult_u0.step1._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step1._15__S  (.I(\mult_u0.step1._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step1._17__S  (.I(\mult_u0.step1._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step1._19__S  (.I(\mult_u0.step1._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step1._21__S  (.I(\mult_u0.step1._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step1._32__I  (.I(\mult_u0.multiplier[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step1.add_sub4_u0.ppa8_u0.d1_0.a2._1__A1  (.I(\mult_u0.multiplier[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step1.add_sub4_u0.x0._1__A1  (.I(\mult_u0.multiplier[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step1.add_sub4_u0.x1._1__A1  (.I(\mult_u0.multiplier[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step1.add_sub4_u0.x2._1__A1  (.I(\mult_u0.multiplier[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step1.add_sub4_u0.x3._1__A1  (.I(\mult_u0.multiplier[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step1.add_sub4_u0.x3._1__A2  (.I(\mult_u0.multiplicand[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step1.add_sub4_u0.x4._1__A1  (.I(\mult_u0.multiplier[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step1.add_sub4_u0.x5._1__A1  (.I(\mult_u0.multiplier[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step1.add_sub4_u0.x6._1__A1  (.I(\mult_u0.multiplier[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step1.add_sub4_u0.x6._1__A2  (.I(\mult_u0.multiplicand[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step2._09__A2  (.I(\mult_u0.Q_s1[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step2._11__S  (.I(\mult_u0.step2._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step2._13__S  (.I(\mult_u0.step2._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step2._15__S  (.I(\mult_u0.step2._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step2._17__S  (.I(\mult_u0.step2._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step2._19__S  (.I(\mult_u0.step2._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step2._21__S  (.I(\mult_u0.step2._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step2._26__I  (.I(\mult_u0.Q_s1[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step2._32__I  (.I(\mult_u0.Q_s1[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step2.add_sub4_u0.ppa8_u0.d1_0.a2._1__A1  (.I(\mult_u0.Q_s1[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step2.add_sub4_u0.x0._1__A1  (.I(\mult_u0.Q_s1[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step2.add_sub4_u0.x1._1__A1  (.I(\mult_u0.Q_s1[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step2.add_sub4_u0.x2._1__A1  (.I(\mult_u0.Q_s1[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step2.add_sub4_u0.x3._1__A1  (.I(\mult_u0.Q_s1[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step2.add_sub4_u0.x4._1__A1  (.I(\mult_u0.Q_s1[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step2.add_sub4_u0.x5._1__A1  (.I(\mult_u0.Q_s1[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step2.add_sub4_u0.x6._1__A1  (.I(\mult_u0.Q_s1[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step3._09__A2  (.I(\mult_u0.Q_s2[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step3._11__S  (.I(\mult_u0.step3._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step3._13__S  (.I(\mult_u0.step3._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step3._15__S  (.I(\mult_u0.step3._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step3._17__S  (.I(\mult_u0.step3._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step3._19__S  (.I(\mult_u0.step3._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step3._21__S  (.I(\mult_u0.step3._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step3._27__I  (.I(\mult_u0.Q_s2[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step3._32__I  (.I(\mult_u0.Q_s2[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step3.add_sub4_u0.ppa8_u0.d1_0.a2._1__A1  (.I(\mult_u0.Q_s2[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step3.add_sub4_u0.x0._1__A1  (.I(\mult_u0.Q_s2[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step3.add_sub4_u0.x1._1__A1  (.I(\mult_u0.Q_s2[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step3.add_sub4_u0.x2._1__A1  (.I(\mult_u0.Q_s2[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step3.add_sub4_u0.x3._1__A1  (.I(\mult_u0.Q_s2[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step3.add_sub4_u0.x4._1__A1  (.I(\mult_u0.Q_s2[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step3.add_sub4_u0.x5._1__A1  (.I(\mult_u0.Q_s2[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step3.add_sub4_u0.x6._1__A1  (.I(\mult_u0.Q_s2[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step4._09__A2  (.I(\mult_u0.Q_s3[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step4._11__S  (.I(\mult_u0.step4._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step4._13__S  (.I(\mult_u0.step4._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step4._15__S  (.I(\mult_u0.step4._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step4._17__S  (.I(\mult_u0.step4._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step4._19__S  (.I(\mult_u0.step4._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step4._21__S  (.I(\mult_u0.step4._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step4._23__S  (.I(\mult_u0.step4._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step4._27__I  (.I(\mult_u0.Q_s3[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step4._32__I  (.I(\mult_u0.Q_s3[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step4.add_sub4_u0.ppa8_u0.d1_0.a2._1__A1  (.I(\mult_u0.Q_s3[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step4.add_sub4_u0.ppa8_u0.s0.xor2_1._1__A2  (.I(\mult_u0.Q_s3[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step4.add_sub4_u0.x0._1__A1  (.I(\mult_u0.Q_s3[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step4.add_sub4_u0.x1._1__A1  (.I(\mult_u0.Q_s3[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step4.add_sub4_u0.x2._1__A1  (.I(\mult_u0.Q_s3[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step4.add_sub4_u0.x3._1__A1  (.I(\mult_u0.Q_s3[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step4.add_sub4_u0.x4._1__A1  (.I(\mult_u0.Q_s3[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step4.add_sub4_u0.x5._1__A1  (.I(\mult_u0.Q_s3[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step4.add_sub4_u0.x6._1__A1  (.I(\mult_u0.Q_s3[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step5._09__A2  (.I(\mult_u0.Q_s4[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step5._13__S  (.I(\mult_u0.step5._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step5._15__S  (.I(\mult_u0.step5._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step5._17__S  (.I(\mult_u0.step5._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step5._19__S  (.I(\mult_u0.step5._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step5._21__S  (.I(\mult_u0.step5._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step5._23__S  (.I(\mult_u0.step5._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step5._32__I  (.I(\mult_u0.Q_s4[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step5.add_sub4_u0.ppa8_u0.d1_0.a2._1__A1  (.I(\mult_u0.Q_s4[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step5.add_sub4_u0.ppa8_u0.s0.xor2_1._1__A2  (.I(\mult_u0.Q_s4[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step5.add_sub4_u0.x0._1__A1  (.I(\mult_u0.Q_s4[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step5.add_sub4_u0.x1._1__A1  (.I(\mult_u0.Q_s4[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step5.add_sub4_u0.x2._1__A1  (.I(\mult_u0.Q_s4[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step5.add_sub4_u0.x3._1__A1  (.I(\mult_u0.Q_s4[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step5.add_sub4_u0.x4._1__A1  (.I(\mult_u0.Q_s4[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step5.add_sub4_u0.x5._1__A1  (.I(\mult_u0.Q_s4[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step6._09__A2  (.I(\mult_u0.Q_s5[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step6._13__S  (.I(\mult_u0.step6._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step6._15__S  (.I(\mult_u0.step6._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step6._17__S  (.I(\mult_u0.step6._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step6._19__S  (.I(\mult_u0.step6._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step6._23__S  (.I(\mult_u0.step6._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step6._32__I  (.I(\mult_u0.Q_s5[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step6.add_sub4_u0.ppa8_u0.d1_0.a2._1__A1  (.I(\mult_u0.Q_s5[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step6.add_sub4_u0.ppa8_u0.s0.xor2_1._1__A2  (.I(\mult_u0.Q_s5[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step6.add_sub4_u0.x0._1__A1  (.I(\mult_u0.Q_s5[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step6.add_sub4_u0.x1._1__A1  (.I(\mult_u0.Q_s5[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step6.add_sub4_u0.x2._1__A1  (.I(\mult_u0.Q_s5[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step6.add_sub4_u0.x3._1__A1  (.I(\mult_u0.Q_s5[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step6.add_sub4_u0.x4._1__A1  (.I(\mult_u0.Q_s5[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step7._09__A2  (.I(\mult_u0.Q_s6[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step7._14__I  (.I(\mult_u0.step7._03_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step7._16__I  (.I(\mult_u0.step7._04_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step7._18__I  (.I(\mult_u0.step7._05_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step7._24__I  (.I(\mult_u0.step7._08_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step7.add_sub4_u0.ppa8_u0.d1_0.a2._1__A1  (.I(\mult_u0.Q_s6[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step7.add_sub4_u0.ppa8_u0.s0.xor2_1._1__A2  (.I(\mult_u0.Q_s6[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step7.add_sub4_u0.x0._1__A1  (.I(\mult_u0.Q_s6[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step7.add_sub4_u0.x1._1__A1  (.I(\mult_u0.Q_s6[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step7.add_sub4_u0.x2._1__A1  (.I(\mult_u0.Q_s6[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.step7.add_sub4_u0.x3._1__A1  (.I(\mult_u0.Q_s6[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_mult_u0.x_sign._1__A1  (.I(\add_u0.b[7] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire1_I (.I(clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_161 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_163 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_181 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_201 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_203 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_214 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_22 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_231 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_240 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_251 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_26 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_261 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_271 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_281 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_30 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_372 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_382 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_391 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_42 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_434 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_44 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_441 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_444 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_461 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_471 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_475 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_484 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_491 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_506 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_541 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_543 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_55 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_552 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_580 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_582 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_614 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_616 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_677 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_679 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_682 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_684 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_135 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_141 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_161 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_165 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_169 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_181 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_211 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_213 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_280 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_288 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_370 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_372 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_395 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_397 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_41 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_448 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_452 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_454 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_473 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_481 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_485 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_487 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_523 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_585 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_613 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_621 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_654 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_662 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_671 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_678 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_686 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_92 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_216 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_232 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_26 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_264 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_272 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_347 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_356 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_360 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_362 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_371 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_405 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_409 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_430 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_460 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_476 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_484 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_488 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_534 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_542 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_570 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_574 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_576 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_593 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_62 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_623 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_627 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_629 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_648 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_650 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_686 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_84 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_86 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_94 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_98 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_102 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_109 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_134 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_204 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_24 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_253 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_257 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_265 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_305 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_309 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_344 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_353 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_382 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_399 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_428 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_444 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_452 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_454 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_465 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_469 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_52 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_535 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_543 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_551 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_553 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_560 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_564 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_634 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_65 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_673 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_681 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_685 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_74 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_90 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_98 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_100 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_109 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_127 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_131 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_135 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_208 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_22 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_220 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_322 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_326 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_334 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_347 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_360 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_362 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_369 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_38 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_385 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_394 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_404 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_42 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_432 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_44 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_440 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_444 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_454 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_456 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_524 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_528 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_530 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_612 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_616 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_624 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_644 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_65 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_650 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_98 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_131 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_135 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_143 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_185 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_189 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_308 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_31 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_319 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_342 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_358 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_362 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_372 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_376 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_403 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_407 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_415 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_425 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_49 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_498 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_506 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_51 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_510 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_517 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_543 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_551 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_573 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_58 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_589 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_593 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_599 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_612 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_620 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_662 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_671 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_678 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_686 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_74 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_94 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_96 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_99 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_134 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_196 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_204 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_208 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_245 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_249 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_288 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_327 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_358 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_36 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_390 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_406 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_414 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_418 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_43 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_455 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_459 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_475 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_483 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_51 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_537 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_545 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_582 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_590 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_594 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_614 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_622 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_76 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_79 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_83 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_87 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_91 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_185 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_265 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_301 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_309 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_372 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_380 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_391 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_406 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_438 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_454 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_489 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_522 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_524 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_541 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_550 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_554 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_581 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_59 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_618 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_630 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_662 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_673 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_681 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_685 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_73 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_77 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_91 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_93 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_99 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_102 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_106 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_114 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_119 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_12 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_127 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_131 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_228 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_230 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_260 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_268 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_272 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_315 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_331 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_339 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_341 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_360 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_364 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_369 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_414 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_418 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_432 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_470 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_474 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_483 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_524 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_540 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_557 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_559 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_587 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_607 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_629 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_648 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_656 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_658 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_671 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_68 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_76 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_97 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_99 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_102 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_109 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_127 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_131 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_141 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_22 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_231 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_239 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_243 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_255 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_259 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_26 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_351 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_438 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_442 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_450 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_452 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_489 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_493 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_533 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_580 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_588 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_592 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_594 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_613 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_617 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_647 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_663 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_675 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_108 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_128 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_132 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_178 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_180 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_228 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_261 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_265 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_273 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_298 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_306 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_308 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_334 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_338 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_347 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_358 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_36 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_374 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_407 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_426 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_44 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_458 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_462 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_488 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_498 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_502 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_510 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_514 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_544 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_552 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_57 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_570 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_601 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_609 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_613 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_615 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_639 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_647 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_651 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_653 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_666 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_674 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_678 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_89 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_91 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_105 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_133 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_153 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_201 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_216 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_220 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_223 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_239 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_255 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_26 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_292 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_30 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_337 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_347 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_374 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_385 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_417 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_430 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_449 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_453 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_461 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_465 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_469 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_487 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_489 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_494 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_538 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_559 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_577 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_62 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_648 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_650 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_146 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_170 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_230 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_238 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_267 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_269 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_299 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_369 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_371 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_374 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_382 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_395 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_403 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_435 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_465 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_469 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_471 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_489 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_505 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_509 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_511 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_518 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_52 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_522 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_524 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_533 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_549 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_557 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_560 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_576 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_578 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_581 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_589 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_593 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_606 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_610 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_614 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_630 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_638 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_642 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_660 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_662 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_114 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_135 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_148 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_152 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_184 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_200 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_208 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_28 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_298 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_306 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_401 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_417 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_426 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_428 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_443 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_460 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_482 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_51 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_55 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_558 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_62 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_640 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_654 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_656 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_685 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_76 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_92 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_113 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_208 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_22 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_24 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_27 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_285 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_292 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_296 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_300 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_302 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_337 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_359 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_366 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_379 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_403 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_417 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_453 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_469 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_477 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_487 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_495 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_531 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_573 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_593 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_74 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_131 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_135 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_195 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_203 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_220 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_224 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_254 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_266 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_342 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_356 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_388 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_396 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_430 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_432 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_447 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_466 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_482 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_537 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_545 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_590 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_648 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_652 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_654 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_684 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_132 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_140 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_146 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_208 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_224 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_238 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_301 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_308 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_334 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_365 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_399 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_403 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_41 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_472 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_476 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_484 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_488 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_512 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_519 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_529 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_580 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_627 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_635 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_643 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_662 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_673 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_677 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_685 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_131 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_194 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_198 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_220 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_224 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_226 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_306 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_310 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_316 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_323 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_364 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_376 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_380 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_415 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_428 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_432 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_436 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_548 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_550 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_557 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_559 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_589 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_613 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_629 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_653 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_684 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_170 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_181 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_255 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_259 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_261 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_303 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_327 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_33 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_334 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_364 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_372 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_382 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_389 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_414 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_418 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_438 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_440 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_447 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_502 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_510 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_537 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_549 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_585 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_589 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_593 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_629 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_633 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_635 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_638 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_652 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_660 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_673 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_681 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_685 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_105 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_109 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_196 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_204 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_208 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_22 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_267 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_271 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_273 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_298 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_336 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_344 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_356 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_358 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_415 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_428 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_430 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_445 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_453 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_455 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_462 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_478 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_505 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_52 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_551 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_553 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_576 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_580 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_582 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_612 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_628 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_68 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_214 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_284 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_31 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_310 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_367 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_393 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_401 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_432 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_448 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_452 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_454 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_461 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_465 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_468 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_476 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_547 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_549 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_579 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_603 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_611 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_642 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_658 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_662 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_679 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_12 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_191 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_237 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_294 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_385 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_389 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_453 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_466 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_474 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_510 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_536 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_554 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_558 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_570 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_623 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_627 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_629 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_63 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_669 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_682 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_686 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_26 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_28 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_465 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_523 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_593 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_63 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_631 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_633 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_679 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_102 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_115 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_166 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_170 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_197 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_199 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_229 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_299 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_303 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_31 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_327 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_382 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_403 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_481 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_483 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_499 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_503 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_517 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_542 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_546 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_587 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_601 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_681 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_685 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_74 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_90 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_98 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_108 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_14 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_315 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_414 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_418 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_473 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_475 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_482 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_568 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_576 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_580 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_616 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_646 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_654 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_658 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_660 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_684 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_102 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_181 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_234 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_271 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_301 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_309 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_350 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_420 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_428 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_438 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_454 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_469 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_477 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_481 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_489 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_497 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_501 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_514 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_518 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_522 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_524 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_533 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_541 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_543 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_594 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_601 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_605 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_607 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_610 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_614 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_618 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_634 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_638 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_654 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_662 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_685 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_98 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_175 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_220 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_250 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_266 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_345 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_426 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_430 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_436 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_452 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_456 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_550 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_558 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_578 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_586 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_590 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_598 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_636 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_666 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_678 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_686 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_74 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_113 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_14 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_23 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_234 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_27 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_302 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_310 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_367 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_391 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_465 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_469 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_57 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_572 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_576 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_592 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_594 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_617 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_649 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_653 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_87 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_105 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_113 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_196 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_204 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_208 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_248 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_343 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_347 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_372 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_374 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_38 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_404 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_438 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_442 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_473 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_489 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_510 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_513 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_545 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_553 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_557 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_559 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_578 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_586 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_590 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_623 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_627 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_629 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_648 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_652 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_662 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_666 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_127 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_157 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_208 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_28 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_287 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_289 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_337 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_391 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_41 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_454 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_489 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_49 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_511 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_524 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_535 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_537 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_546 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_554 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_569 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_585 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_612 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_628 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_646 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_663 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_685 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_131 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_178 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_180 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_267 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_271 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_273 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_342 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_360 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_364 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_424 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_454 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_470 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_478 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_482 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_512 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_516 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_525 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_529 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_589 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_593 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_601 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_609 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_613 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_622 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_22 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_26 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_28 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_39 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_420 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_522 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_524 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_529 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_548 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_552 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_583 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_593 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_663 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_85 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_117 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_133 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_197 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_218 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_266 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_299 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_38 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_426 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_434 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_465 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_48 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_481 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_485 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_487 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_519 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_52 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_523 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_525 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_547 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_551 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_572 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_576 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_58 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_605 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_62 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_627 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_629 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_646 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_684 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_84 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_135 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_14 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_16 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_222 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_234 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_266 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_270 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_292 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_356 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_359 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_361 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_459 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_52 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_523 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_559 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_568 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_58 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_62 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_74 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_77 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_81 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_141 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_218 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_234 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_252 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_301 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_305 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_309 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_31 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_362 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_366 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_374 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_382 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_41 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_435 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_443 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_447 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_465 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_467 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_47 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_50 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_509 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_513 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_539 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_547 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_551 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_555 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_583 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_631 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_682 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_686 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_124 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_128 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_150 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_243 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_270 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_344 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_356 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_38 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_391 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_404 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_42 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_438 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_46 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_482 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_499 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_507 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_538 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_540 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_553 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_564 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_583 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_599 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_603 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_605 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_62 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_638 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_654 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_658 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_92 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_94 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_119 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_126 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_134 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_167 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_216 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_220 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_236 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_251 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_268 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_353 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_406 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_41 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_48 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_507 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_511 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_519 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_52 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_523 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_535 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_541 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_55 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_557 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_582 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_586 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_59 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_594 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_605 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_609 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_61 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_611 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_627 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_631 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_647 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_663 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_685 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_150 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_178 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_182 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_184 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_191 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_292 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_299 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_307 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_316 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_323 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_339 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_347 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_38 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_385 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_40 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_410 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_483 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_487 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_489 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_542 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_546 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_570 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_574 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_576 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_606 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_616 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_624 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_628 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_648 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_678 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_682 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_686 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_84 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_102 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_113 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_16 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_181 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_197 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_20 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_214 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_24 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_270 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_302 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_337 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_347 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_409 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_425 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_429 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_445 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_453 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_473 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_480 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_512 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_516 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_518 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_55 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_572 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_580 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_588 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_592 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_594 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_599 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_85 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_87 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_94 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_11 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_220 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_257 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_320 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_360 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_362 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_369 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_385 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_437 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_441 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_445 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_453 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_460 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_522 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_542 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_546 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_550 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_558 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_566 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_644 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_65 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_119 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_186 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_190 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_324 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_362 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_4 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_413 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_415 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_444 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_448 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_452 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_454 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_459 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_466 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_47 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_470 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_472 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_477 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_479 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_502 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_506 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_51 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_553 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_585 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_593 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_605 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_609 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_640 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_646 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_662 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_130 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_148 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_156 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_160 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_198 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_245 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_288 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_354 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_375 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_412 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_446 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_479 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_487 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_489 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_50 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_512 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_548 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_594 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_598 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_600 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_634 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_645 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_149 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_165 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_23 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_243 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_252 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_27 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_289 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_293 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_301 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_309 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_31 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_323 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_336 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_340 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_379 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_41 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_447 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_461 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_463 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_472 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_488 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_496 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_503 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_511 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_519 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_523 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_531 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_533 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_536 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_544 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_546 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_553 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_585 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_593 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_91 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_95 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_99 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_121 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_150 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_156 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_186 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_243 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_246 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_270 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_288 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_294 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_326 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_330 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_339 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_38 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_406 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_414 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_418 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_42 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_442 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_450 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_454 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_485 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_489 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_537 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_541 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_549 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_558 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_568 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_572 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_58 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_581 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_595 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_627 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_629 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_668 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_676 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_684 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_84 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_92 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_102 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_140 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_152 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_156 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_167 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_187 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_203 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_237 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_26 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_288 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_30 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_306 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_327 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_369 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_373 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_377 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_395 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_407 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_411 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_420 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_434 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_438 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_440 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_47 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_49 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_52 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_56 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_583 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_585 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_592 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_594 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_60 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_64 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_68 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_76 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_84 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_100 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_115 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_128 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_132 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_183 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_191 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_237 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_283 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_288 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_296 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_300 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_343 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_403 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_405 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_412 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_423 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_425 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_465 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_469 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_471 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_505 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_539 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_561 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_593 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_613 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_629 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_637 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_647 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_651 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_653 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_660 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_675 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_89 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_91 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_121 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_14 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_200 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_216 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_218 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_223 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_227 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_260 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_292 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_308 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_310 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_323 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_339 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_347 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_374 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_376 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_399 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_403 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_417 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_435 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_441 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_445 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_46 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_477 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_485 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_489 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_498 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_514 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_568 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_583 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_585 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_592 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_600 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_604 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_606 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_62 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_625 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_629 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_677 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_685 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_84 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_100 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_121 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_125 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_129 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_131 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_161 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_169 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_187 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_251 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_259 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_266 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_270 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_298 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_305 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_335 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_367 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_395 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_437 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_439 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_449 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_453 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_47 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_473 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_475 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_484 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_522 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_524 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_548 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_558 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_566 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_573 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_593 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_605 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_609 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_663 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_681 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_685 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_77 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_81 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_83 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_127 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_135 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_27 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_270 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_338 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_360 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_370 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_386 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_390 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_404 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_408 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_460 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_47 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_494 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_51 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_545 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_547 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_554 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_558 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_566 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_587 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_603 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_616 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_629 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_650 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_652 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_685 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_96 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_127 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_131 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_166 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_168 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_181 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_301 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_309 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_342 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_358 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_374 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_382 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_426 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_429 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_439 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_441 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_452 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_454 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_474 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_494 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_524 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_605 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_624 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_628 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_644 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_85 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_93 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_97 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_128 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_132 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_150 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_156 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_198 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_202 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_288 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_292 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_300 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_304 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_323 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_341 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_343 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_39 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_390 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_394 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_401 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_403 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_410 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_418 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_430 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_469 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_485 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_489 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_525 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_533 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_549 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_55 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_553 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_587 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_623 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_627 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_629 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_63 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_636 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_638 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_684 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_119 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_191 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_195 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_228 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_232 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_240 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_251 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_255 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_259 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_267 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_30 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_305 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_319 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_328 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_354 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_361 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_378 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_407 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_414 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_424 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_452 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_454 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_471 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_49 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_502 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_518 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_522 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_524 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_535 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_578 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_582 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_586 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_594 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_601 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_609 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_625 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_633 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_673 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_681 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_685 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_90 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_94 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_96 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_127 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_135 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_202 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_261 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_265 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_273 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_298 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_302 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_345 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_360 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_364 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_372 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_376 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_403 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_468 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_476 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_478 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_487 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_489 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_543 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_551 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_553 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_613 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_620 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_624 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_628 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_76 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_92 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_94 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_109 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_130 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_146 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_181 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_211 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_215 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_26 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_284 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_323 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_331 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_376 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_378 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_403 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_407 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_420 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_424 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_462 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_466 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_470 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_49 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_501 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_51 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_517 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_533 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_549 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_557 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_559 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_589 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_655 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_663 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_671 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_678 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_686 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_87 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_91 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_99 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_130 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_166 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_181 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_197 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_268 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_272 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_284 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_337 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_345 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_388 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_407 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_415 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_43 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_430 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_434 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_453 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_473 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_477 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_51 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_539 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_543 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_551 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_555 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_557 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_612 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_628 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_636 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_125 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_129 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_132 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_150 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_156 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_218 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_222 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_226 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_230 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_234 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_238 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_25 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_257 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_275 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_296 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_336 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_342 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_356 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_360 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_364 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_372 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_41 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_410 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_414 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_418 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_426 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_465 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_469 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_475 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_485 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_489 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_496 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_515 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_519 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_523 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_55 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_57 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_610 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_614 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_618 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_665 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_681 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_685 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_87 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_91 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_109 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_118 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_129 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_161 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_169 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_183 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_199 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_235 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_239 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_243 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_265 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_295 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_435 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_439 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_441 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_444 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_452 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_454 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_465 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_498 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_514 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_518 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_547 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_551 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_555 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_559 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_561 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_628 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_645 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_649 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_653 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_655 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_662 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_679 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_135 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_14 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_148 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_156 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_182 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_198 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_22 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_230 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_246 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_250 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_341 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_372 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_402 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_418 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_467 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_473 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_489 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_523 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_54 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_559 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_578 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_604 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_608 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_624 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_628 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_640 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_644 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_119 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_121 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_189 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_251 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_253 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_289 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_293 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_295 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_298 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_350 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_447 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_465 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_498 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_514 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_518 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_545 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_557 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_589 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_593 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_615 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_625 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_657 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_679 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_78 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_82 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_84 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_128 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_130 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_202 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_249 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_275 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_330 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_418 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_426 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_434 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_438 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_47 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_489 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_496 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_55 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_558 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_57 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_580 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_582 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_589 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_598 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_625 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_629 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_648 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_656 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_76 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_114 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_146 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_196 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_200 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_208 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_261 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_265 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_301 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_309 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_31 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_324 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_361 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_377 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_41 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_421 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_507 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_523 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_535 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_539 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_561 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_57 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_590 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_594 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_603 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_640 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_644 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_685 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_87 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_91 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_99 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_126 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_130 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_220 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_228 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_29 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_372 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_403 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_430 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_434 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_464 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_480 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_488 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_525 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_541 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_545 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_547 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_577 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_581 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_585 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_592 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_596 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_61 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_627 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_629 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_92 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_94 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_12 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_166 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_197 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_229 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_239 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_243 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_280 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_284 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_288 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_304 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_319 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_395 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_397 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_41 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_452 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_454 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_46 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_494 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_499 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_507 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_517 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_539 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_54 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_543 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_575 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_58 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_631 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_635 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_644 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_660 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_671 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_685 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_92 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_96 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_98 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_105 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_146 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_156 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_159 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_163 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_187 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_203 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_216 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_232 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_240 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_246 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_253 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_26 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_269 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_288 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_304 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_316 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_318 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_410 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_412 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_482 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_496 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_54 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_594 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_610 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_612 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_615 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_623 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_627 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_629 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_656 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_679 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_76 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_84 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_97 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_157 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_181 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_194 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_198 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_200 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_23 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_230 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_238 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_259 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_267 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_303 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_307 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_359 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_375 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_453 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_461 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_465 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_520 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_524 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_539 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_555 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_571 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_575 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_579 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_592 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_594 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_601 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_609 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_61 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_611 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_641 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_643 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_646 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_654 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_656 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_685 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_118 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_133 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_150 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_169 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_198 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_216 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_223 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_227 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_229 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_271 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_29 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_324 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_328 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_344 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_360 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_362 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_405 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_413 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_417 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_42 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_424 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_44 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_454 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_458 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_462 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_483 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_487 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_489 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_504 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_506 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_540 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_609 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_613 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_629 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_64 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_644 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_68 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_109 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_112 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_14 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_181 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_183 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_186 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_190 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_21 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_251 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_259 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_267 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_269 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_301 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_305 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_308 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_327 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_330 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_334 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_338 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_342 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_356 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_372 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_375 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_391 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_393 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_423 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_427 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_431 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_435 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_439 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_443 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_447 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_451 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_494 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_498 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_502 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_506 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_51 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_510 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_514 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_518 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_524 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_535 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_603 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_639 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_643 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_653 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_99 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_127 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_129 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_159 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_261 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_285 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_289 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_363 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_379 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_403 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_407 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_409 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_41 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_439 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_496 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_512 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_535 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_539 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_572 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_580 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_584 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_586 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_63 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_685 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_95 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_105 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_12 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_124 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_131 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_181 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_185 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_189 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_228 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_230 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_233 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_235 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_270 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_298 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_300 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_33 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_334 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_338 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_356 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_395 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_409 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_413 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_417 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_429 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_445 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_449 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_485 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_489 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_502 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_509 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_513 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_536 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_540 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_570 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_574 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_619 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_627 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_629 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_638 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_642 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_646 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_65 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_675 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_130 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_134 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_166 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_168 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_273 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_30 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_305 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_360 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_376 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_395 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_399 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_401 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_408 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_440 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_448 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_452 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_454 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_465 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_469 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_471 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_506 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_514 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_518 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_529 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_544 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_548 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_550 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_557 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_589 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_593 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_640 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_656 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_673 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_681 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_685 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_96 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_98 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_114 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_127 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_131 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_133 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_183 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_27 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_31 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_327 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_341 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_360 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_372 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_374 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_389 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_393 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_415 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_438 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_471 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_475 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_477 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_480 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_488 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_500 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_516 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_52 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_524 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_543 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_559 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_56 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_570 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_586 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_590 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_592 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_599 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_607 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_611 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_640 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_650 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_682 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_686 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_84 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_92 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_169 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_189 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_222 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_230 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_234 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_238 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_266 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_298 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_323 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_330 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_332 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_391 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_429 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_445 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_453 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_47 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_489 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_499 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_515 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_523 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_54 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_547 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_549 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_558 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_570 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_572 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_579 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_58 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_583 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_592 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_594 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_60 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_605 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_609 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_611 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_624 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_628 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_660 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_96 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_102 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_106 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_119 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_135 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_203 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_220 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_224 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_239 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_251 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_260 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_273 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_284 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_291 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_307 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_358 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_395 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_430 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_434 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_471 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_516 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_532 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_566 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_575 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_608 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_616 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_624 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_628 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_78 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_94 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_12 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_121 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_153 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_169 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_267 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_321 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_323 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_326 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_330 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_380 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_395 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_397 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_404 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_406 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_409 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_413 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_415 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_432 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_449 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_453 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_519 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_523 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_535 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_539 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_547 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_551 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_594 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_619 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_651 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_659 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_663 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_73 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_77 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_93 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_124 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_126 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_133 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_148 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_156 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_160 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_228 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_246 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_248 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_255 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_26 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_269 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_336 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_358 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_390 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_398 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_452 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_46 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_482 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_50 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_512 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_516 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_54 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_548 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_56 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_608 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_624 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_628 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_63 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_168 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_185 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_189 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_208 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_238 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_267 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_269 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_361 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_377 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_39 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_443 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_447 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_46 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_48 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_490 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_494 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_496 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_523 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_559 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_567 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_571 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_579 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_78 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_82 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_84 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_121 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_146 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_166 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_168 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_189 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_354 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_361 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_365 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_367 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_374 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_382 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_413 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_417 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_440 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_472 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_488 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_500 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_504 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_559 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_115 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_117 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_120 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_124 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_128 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_132 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_148 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_216 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_220 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_224 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_24 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_26 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_292 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_296 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_300 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_310 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_316 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_319 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_323 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_339 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_347 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_372 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_374 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_379 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_411 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_47 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_484 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_488 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_496 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_500 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_504 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_51 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_536 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_544 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_548 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_558 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_56 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_566 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_596 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_62 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_668 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_684 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_84 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_86 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_115 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_156 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_164 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_166 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_200 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_232 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_240 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_251 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_259 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_295 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_368 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_393 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_425 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_427 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_440 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_448 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_452 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_454 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_464 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_496 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_500 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_502 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_509 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_85 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_100 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_102 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_109 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_125 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_133 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_204 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_208 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_219 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_273 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_294 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_327 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_366 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_370 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_374 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_376 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_406 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_414 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_418 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_456 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_460 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_476 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_484 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_488 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_538 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_554 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_558 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_96 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_121 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_153 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_189 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_191 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_198 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_200 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_259 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_298 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_302 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_310 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_337 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_350 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_361 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_377 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_403 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_423 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_453 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_472 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_501 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_514 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_523 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_533 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_565 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_581 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_589 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_593 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_85 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_89 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_128 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_132 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_176 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_178 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_201 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_216 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_218 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_275 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_358 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_390 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_406 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_426 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_439 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_482 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_516 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_531 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_547 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_555 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_559 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_135 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_165 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_199 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_203 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_235 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_243 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_281 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_283 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_306 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_333 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_337 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_345 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_357 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_365 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_373 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_377 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_416 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_424 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_488 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_508 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_516 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_524 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_85 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_89 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_148 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_186 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_203 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_260 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_294 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_301 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_305 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_336 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_370 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_400 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_406 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_414 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_418 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_426 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_435 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_473 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_481 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_483 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_50 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_504 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_536 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_54 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_552 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_56 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_63 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_84 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_86 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_141 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_215 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_251 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_255 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_309 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_380 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_391 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_418 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_426 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_430 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_438 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_450 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_454 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_461 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_512 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_516 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_524 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_57 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_92 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_105 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_118 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_128 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_132 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_197 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_218 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_267 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_269 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_284 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_305 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_309 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_316 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_376 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_388 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_390 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_453 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_471 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_498 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_50 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_530 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_546 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_554 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_558 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_58 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_68 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_102 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_228 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_255 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_265 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_273 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_275 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_306 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_357 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_365 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_381 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_437 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_447 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_465 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_495 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_511 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_519 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_523 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_57 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_87 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_89 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_120 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_148 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_152 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_159 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_175 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_191 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_216 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_288 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_378 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_410 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_434 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_470 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_486 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_102 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_115 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_118 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_131 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_135 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_143 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_183 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_187 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_191 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_195 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_199 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_203 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_236 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_240 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_255 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_319 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_326 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_339 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_355 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_363 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_403 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_407 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_444 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_452 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_461 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_499 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_515 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_523 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_531 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_539 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_543 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_545 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_575 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_585 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_589 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_61 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_647 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_65 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_663 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_674 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_682 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_686 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_76 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_79 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_83 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_95 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_184 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_188 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_195 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_197 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_90_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_90_210 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_283 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_299 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_307 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_90_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_90_387 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_423 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_431 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_433 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_90_487 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_519 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_523 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_73 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_75 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_146 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_166 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_168 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_181 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_185 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_189 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_218 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_234 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_322 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_337 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_345 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_356 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_389 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_397 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_415 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_480 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_484 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_488 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_84 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_143 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_145 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_194 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_210 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_259 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_272 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_293 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_309 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_323 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_331 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_335 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_337 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_344 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_348 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_350 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_365 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_367 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_399 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_415 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_423 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_427 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_150 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_202 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_216 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_267 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_293 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_335 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_343 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_347 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_428 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_432 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_469 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_485 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_489 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_168 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_189 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_196 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_204 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_237 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_249 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_271 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_284 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_299 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_303 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_305 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_373 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_380 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_384 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_399 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_430 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_166 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_199 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_203 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_364 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_366 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_394 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_401 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_417 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_424 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_437 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_439 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_95_458 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_626 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_95_632 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_664 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_680 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_226 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_253 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_266 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_280 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_288 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_292 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_300 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_308 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_349 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_357 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_361 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_363 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_370 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_374 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_376 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_379 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_383 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_393 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_425 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_433 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_443 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_445 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_452 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_454 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_457 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_521 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_527 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_591 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_597 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_661 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_667 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_683 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_687 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_240 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_248 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_250 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_253 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_269 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_271 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_308 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_342 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_36 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_376 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_410 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_444 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_478 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_512 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_546 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_580 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_614 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_648 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_682 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_686 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_125 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_127 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_156 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_160 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_164 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_168 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_170 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_200 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_204 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_208 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_21 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_220 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_222 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_225 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_227 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_257 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_273 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_346 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_352 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_356 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_39 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_395 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_399 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_403 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_419 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_422 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_426 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_43 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_456 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_460 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_492 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_496 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_50 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_503 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_511 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_513 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_550 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_556 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_562 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_58 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_588 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_620 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_83 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_98 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_99 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_131 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Left_143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Right_45 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Left_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Right_46 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Left_145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Right_47 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Left_146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Right_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Left_147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Right_49 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Left_148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Right_50 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Left_149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Right_51 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Left_150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Right_52 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Left_151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Right_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Left_152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Right_54 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Left_153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Right_55 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Left_154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Right_56 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Left_155 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Right_57 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Left_156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Right_58 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Left_157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Right_59 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Left_158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Right_60 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Left_159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Right_61 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Left_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Right_62 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Left_161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Right_63 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Left_162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Right_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Left_163 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Right_65 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Left_164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Right_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Left_165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Right_67 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Left_166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Right_68 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Left_167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Right_69 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Left_168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Right_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Left_169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Right_71 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Left_170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Right_72 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Left_171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Right_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Left_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Right_74 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Left_173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Right_75 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Left_174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Right_76 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Left_175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Right_77 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Left_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Right_78 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Left_177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Right_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Left_178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Right_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_Left_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_Right_81 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_Left_180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_Right_82 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Left_181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Right_83 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Left_182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Right_84 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Left_183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Right_85 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Left_184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Right_86 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_Left_185 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_Right_87 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_Left_186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_Right_88 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_Left_187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_Right_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_Left_188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_Right_90 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_Left_189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_Right_91 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_Left_190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_Right_92 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_Left_191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_Right_93 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_Left_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_Right_94 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_Left_193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_Right_95 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_Left_194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_Right_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_Left_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_Right_97 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_313 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_314 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_315 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_316 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_317 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_318 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_319 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_320 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_321 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_322 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_323 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_324 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_325 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_326 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_327 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_328 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_329 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_330 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_331 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_332 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_333 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_334 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_335 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_336 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_337 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_338 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_339 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_340 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_341 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_342 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_343 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_344 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_345 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_346 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_347 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_348 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_349 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_350 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_351 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_352 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_353 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_354 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_355 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_356 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_357 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_358 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_359 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_360 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_361 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_362 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_363 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_364 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_365 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_366 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_367 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_368 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_369 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_370 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_371 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_372 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_373 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_374 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_375 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_376 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_377 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_378 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_379 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_380 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_381 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_382 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_383 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_384 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_385 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_386 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_387 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_388 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_389 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_390 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_391 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_392 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_393 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_394 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_395 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_217 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_219 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_396 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_397 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_398 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_399 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_400 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_401 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_402 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_403 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_404 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_405 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_406 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_407 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_408 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_409 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_410 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_411 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_412 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_413 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_414 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_415 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_416 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_417 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_418 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_419 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_420 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_421 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_422 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_423 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_424 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_425 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_426 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_427 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_428 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_429 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_430 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_431 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_432 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_433 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_434 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_435 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_436 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_437 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_438 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_439 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_440 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_441 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_442 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_443 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_444 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_445 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_446 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_447 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_448 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_449 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_450 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_451 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_452 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_453 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_454 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_455 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_456 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_457 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_458 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_459 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_460 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_461 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_462 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_463 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_464 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_465 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_466 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_467 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_468 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_469 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_470 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_471 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_472 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_473 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_474 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_475 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_476 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_477 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_478 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_479 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_480 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_481 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_482 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_483 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_484 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_485 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_486 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_487 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_488 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_489 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_490 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_227 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_491 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_492 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_493 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_494 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_495 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_496 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_497 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_498 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_499 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_500 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_501 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_502 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_503 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_504 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_505 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_506 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_507 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_508 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_509 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_510 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_511 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_512 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_513 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_514 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_515 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_516 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_517 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_518 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_519 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_520 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_521 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_522 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_523 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_524 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_525 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_526 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_527 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_528 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_529 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_530 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_531 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_532 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_533 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_534 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_535 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_536 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_537 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_538 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_539 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_540 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_541 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_542 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_543 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_544 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_545 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_546 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_547 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_548 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_549 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_550 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_551 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_552 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_553 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_554 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_555 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_556 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_557 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_558 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_559 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_560 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_561 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_562 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_563 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_564 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_565 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_566 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_567 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_568 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_569 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_570 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_571 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_572 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_573 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_574 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_575 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_576 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_577 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_578 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_579 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_580 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_581 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_582 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_583 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_584 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_585 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_235 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_586 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_587 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_588 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_589 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_590 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_591 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_592 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_593 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_594 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_595 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_596 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_597 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_598 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_599 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_600 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_601 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_602 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_603 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_604 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_605 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_606 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_607 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_608 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_609 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_610 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_611 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_612 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_613 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_614 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_615 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_616 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_617 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_618 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_619 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_620 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_621 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_622 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_623 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_624 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_625 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_626 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_627 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_628 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_629 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_630 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_631 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_632 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_633 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_634 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_635 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_636 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_637 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_638 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_639 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_640 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_641 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_642 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_643 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_644 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_645 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_646 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_647 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_648 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_649 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_650 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_651 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_652 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_653 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_654 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_655 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_656 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_657 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_658 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_659 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_660 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_661 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_662 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_663 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_664 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_665 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_666 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_667 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_668 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_669 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_670 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_671 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_672 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_673 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_674 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_675 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_676 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_677 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_678 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_679 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_680 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_681 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_682 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_683 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_684 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_685 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_686 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_687 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_688 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_689 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_690 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_691 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_692 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_693 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_694 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_695 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_696 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_697 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_698 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_699 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_700 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_701 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_702 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_703 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_704 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_705 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_706 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_707 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_708 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_709 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_710 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_711 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_712 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_713 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_714 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_715 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_716 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_717 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_718 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_719 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_720 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_721 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_722 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_723 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_724 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_725 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_726 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_727 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_728 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_729 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_730 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_731 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_732 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_733 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_734 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_735 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_736 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_737 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_738 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_739 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_740 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_741 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_742 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_743 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_744 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_745 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_746 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_747 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_748 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_749 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_750 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_751 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_752 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_753 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_754 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_755 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_756 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_757 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_758 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_759 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_760 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_761 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_762 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_763 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_764 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_765 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_766 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_767 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_768 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_769 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_770 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_771 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_772 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_773 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_774 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_775 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_259 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_776 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_777 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_778 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_779 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_780 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_781 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_782 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_783 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_784 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_785 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_786 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_787 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_788 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_789 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_790 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_791 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_792 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_793 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_794 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_795 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_796 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_797 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_798 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_799 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_800 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_801 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_802 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_803 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_804 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_805 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_806 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_807 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_808 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_809 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_810 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_811 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_812 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_813 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_814 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_815 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_816 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_817 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_818 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_819 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_820 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_821 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_822 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_823 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_824 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_825 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_826 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_827 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_828 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_829 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_830 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_831 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_832 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_833 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_834 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_835 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_836 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_837 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_838 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_839 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_840 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_841 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_842 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_843 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_844 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_845 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_846 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_847 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_848 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_849 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_850 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_851 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_852 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_853 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_854 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_855 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_856 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_857 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_858 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_859 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_860 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_861 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_862 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_863 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_864 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_865 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_866 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_867 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_868 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_869 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_870 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_267 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_871 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_872 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_873 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_874 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_875 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_876 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_877 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_878 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_879 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_880 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_881 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_882 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_883 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_884 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_885 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_886 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_887 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_888 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_889 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_890 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_891 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_892 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_893 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_894 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_895 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_896 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_897 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_898 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_899 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_900 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_901 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_902 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_903 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_904 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_905 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_906 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_907 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_908 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_909 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_910 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_911 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_912 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_913 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_914 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_915 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_916 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_917 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_918 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_919 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_920 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_921 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_922 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_923 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_924 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_925 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_926 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_927 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_928 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_929 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_930 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_931 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_932 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_933 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_934 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_935 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_936 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_937 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_938 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_939 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_940 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_941 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_942 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_943 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_944 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_945 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_946 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_947 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_948 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_949 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_950 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_951 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_952 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_953 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_954 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_955 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_956 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_957 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_958 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_959 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_960 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_961 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_962 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_963 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_964 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_965 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_273 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_966 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_967 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_968 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_969 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_970 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_971 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_972 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_973 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_974 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_975 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_976 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_977 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_978 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_979 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_980 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_981 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_982 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_983 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_984 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_985 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_986 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_987 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_988 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_989 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_990 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_991 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_992 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_993 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_994 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1000 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1001 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1002 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_1003 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_995 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_996 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_997 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_998 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_999 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1004 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1005 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1006 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1007 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1008 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1009 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1010 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1011 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1012 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_1013 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1014 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1015 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1016 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1017 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1018 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1019 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1020 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1021 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_1022 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1023 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1024 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1025 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1026 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1027 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1028 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1029 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1030 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1031 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_1032 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1033 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1034 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1035 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1036 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1037 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1038 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1039 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1040 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_1041 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1042 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1043 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1044 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1045 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1046 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1047 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1048 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1049 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1050 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_1051 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1052 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1053 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1054 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1055 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1056 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1057 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1058 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1059 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_1060 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1061 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1062 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1063 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1064 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1065 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1066 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1067 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1068 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1069 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_1070 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1071 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1072 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1073 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1074 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1075 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1076 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1077 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1078 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_1079 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1080 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1081 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1082 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1083 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1084 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1085 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1086 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1087 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1088 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_1089 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1090 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1091 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1092 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1093 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1094 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1095 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1096 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1097 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_1098 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1099 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_1108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_1117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_1127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1131 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_1147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_299 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _174_ (.I(net62),
    .Z(_043_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _175_ (.I(_043_),
    .ZN(_044_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _176_ (.A1(net33),
    .A2(net60),
    .A3(net61),
    .Z(_045_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _177_ (.I(net9),
    .ZN(_046_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _178_ (.A1(net14),
    .A2(net13),
    .A3(net16),
    .A4(net15),
    .ZN(_047_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _179_ (.A1(net11),
    .A2(net10),
    .ZN(_048_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _180_ (.A1(_046_),
    .A2(net8),
    .A3(_047_),
    .A4(_048_),
    .ZN(_049_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _181_ (.A1(net25),
    .A2(net24),
    .ZN(_050_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _182_ (.A1(net18),
    .A2(net17),
    .A3(net20),
    .A4(net19),
    .ZN(_051_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _183_ (.A1(net22),
    .A2(net21),
    .A3(_050_),
    .A4(_051_),
    .ZN(_052_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _184_ (.A1(net28),
    .A2(net27),
    .A3(net30),
    .A4(net29),
    .ZN(_053_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _185_ (.A1(net12),
    .A2(net1),
    .A3(net23),
    .ZN(_054_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _186_ (.A1(net26),
    .A2(_053_),
    .A3(_054_),
    .ZN(_055_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _187_ (.A1(net32),
    .A2(net31),
    .A3(net3),
    .A4(net2),
    .ZN(_056_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _188_ (.A1(net5),
    .A2(net4),
    .A3(net7),
    .A4(net6),
    .ZN(_057_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _189_ (.A1(_056_),
    .A2(_057_),
    .ZN(_058_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _190_ (.A1(_049_),
    .A2(_052_),
    .A3(_055_),
    .A4(_058_),
    .ZN(_059_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _191_ (.I(_059_),
    .Z(_060_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _192_ (.A1(_044_),
    .A2(_045_),
    .A3(_060_),
    .ZN(_061_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _193_ (.I0(net50),
    .I1(\sel[0] ),
    .S(_061_),
    .Z(_062_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _194_ (.I(_062_),
    .Z(_000_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _195_ (.I0(net51),
    .I1(\sel[1] ),
    .S(_061_),
    .Z(_063_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _196_ (.I(_063_),
    .Z(_001_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _197_ (.I(\sel_d8[0] ),
    .Z(_064_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _198_ (.I(\sel_d8[1] ),
    .Z(_065_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_4 _199_ (.A1(_064_),
    .A2(_065_),
    .ZN(_066_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _200_ (.A1(_064_),
    .A2(_065_),
    .ZN(_067_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _201_ (.A1(_065_),
    .A2(\mult_add_u0.out[0] ),
    .ZN(_068_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _202_ (.A1(_067_),
    .A2(_068_),
    .ZN(_069_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _203_ (.A1(_064_),
    .A2(\mul_out_d0[0] ),
    .B1(\add_out_d7[0] ),
    .B2(_066_),
    .C(_069_),
    .ZN(_070_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _204_ (.A1(\out[0] ),
    .A2(_067_),
    .B(_044_),
    .ZN(_071_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _205_ (.A1(_070_),
    .A2(_071_),
    .ZN(_002_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _206_ (.A1(_065_),
    .A2(\mult_add_u0.out[1] ),
    .ZN(_072_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _207_ (.A1(_067_),
    .A2(_072_),
    .ZN(_073_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _208_ (.A1(_064_),
    .A2(\mul_out_d0[1] ),
    .B1(\add_out_d7[1] ),
    .B2(_066_),
    .C(_073_),
    .ZN(_074_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _209_ (.A1(\out[1] ),
    .A2(_067_),
    .B(_044_),
    .ZN(_075_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _210_ (.A1(_074_),
    .A2(_075_),
    .ZN(_003_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _211_ (.A1(_065_),
    .A2(\mult_add_u0.out[2] ),
    .ZN(_076_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _212_ (.A1(_067_),
    .A2(_076_),
    .ZN(_077_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _213_ (.A1(_064_),
    .A2(\mul_out_d0[2] ),
    .B1(\add_out_d7[2] ),
    .B2(_066_),
    .C(_077_),
    .ZN(_078_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _214_ (.A1(\out[2] ),
    .A2(_067_),
    .B(_044_),
    .ZN(_079_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _215_ (.A1(_078_),
    .A2(_079_),
    .ZN(_004_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _216_ (.A1(_065_),
    .A2(\mult_add_u0.out[3] ),
    .ZN(_080_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _217_ (.A1(_067_),
    .A2(_080_),
    .ZN(_081_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _218_ (.A1(_064_),
    .A2(\mul_out_d0[3] ),
    .B1(\add_out_d7[3] ),
    .B2(_066_),
    .C(_081_),
    .ZN(_082_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _219_ (.A1(\out[3] ),
    .A2(_067_),
    .B(_044_),
    .ZN(_083_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _220_ (.A1(_082_),
    .A2(_083_),
    .ZN(_005_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _221_ (.A1(_065_),
    .A2(\mult_add_u0.out[4] ),
    .ZN(_084_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _222_ (.A1(_067_),
    .A2(_084_),
    .ZN(_085_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _223_ (.A1(_064_),
    .A2(\mul_out_d0[4] ),
    .B1(\add_out_d7[4] ),
    .B2(_066_),
    .C(_085_),
    .ZN(_086_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _224_ (.A1(\out[4] ),
    .A2(_067_),
    .B(_044_),
    .ZN(_087_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _225_ (.A1(_086_),
    .A2(_087_),
    .ZN(_006_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _226_ (.A1(_065_),
    .A2(\mult_add_u0.out[5] ),
    .ZN(_088_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _227_ (.A1(_067_),
    .A2(_088_),
    .ZN(_089_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _228_ (.A1(_064_),
    .A2(\mul_out_d0[5] ),
    .B1(\add_out_d7[5] ),
    .B2(_066_),
    .C(_089_),
    .ZN(_090_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _229_ (.A1(\out[5] ),
    .A2(_067_),
    .B(_044_),
    .ZN(_091_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _230_ (.A1(_090_),
    .A2(_091_),
    .ZN(_007_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _231_ (.A1(_065_),
    .A2(\mult_add_u0.out[6] ),
    .ZN(_092_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _232_ (.A1(_067_),
    .A2(_092_),
    .ZN(_093_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _233_ (.A1(_064_),
    .A2(\mul_out_d0[6] ),
    .B1(\add_out_d7[6] ),
    .B2(_066_),
    .C(_093_),
    .ZN(_094_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _234_ (.A1(\out[6] ),
    .A2(_067_),
    .B(_044_),
    .ZN(_095_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _235_ (.A1(_094_),
    .A2(_095_),
    .ZN(_008_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _236_ (.A1(_065_),
    .A2(\mult_add_u0.out[7] ),
    .ZN(_096_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _237_ (.A1(_067_),
    .A2(_096_),
    .ZN(_097_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _238_ (.A1(_064_),
    .A2(\mul_out_d0[7] ),
    .B1(\add_out_d7[7] ),
    .B2(_066_),
    .C(_097_),
    .ZN(_098_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _239_ (.A1(\out[7] ),
    .A2(_067_),
    .B(_044_),
    .ZN(_099_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _240_ (.A1(_098_),
    .A2(_099_),
    .ZN(_009_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _241_ (.I(net34),
    .ZN(_100_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _242_ (.A1(_045_),
    .A2(_060_),
    .Z(_101_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _243_ (.I(_101_),
    .Z(_102_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _244_ (.I(_102_),
    .Z(_103_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _245_ (.I(_045_),
    .Z(_104_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 _246_ (.I(_060_),
    .Z(_105_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _247_ (.A1(_104_),
    .A2(_105_),
    .B(\add_u0.a[0] ),
    .ZN(_106_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _248_ (.I(_043_),
    .Z(_107_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _249_ (.A1(_100_),
    .A2(_103_),
    .B(_106_),
    .C(_107_),
    .ZN(_010_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _250_ (.I(net45),
    .ZN(_108_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _251_ (.A1(_104_),
    .A2(_105_),
    .B(\add_u0.a[1] ),
    .ZN(_109_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _252_ (.A1(_108_),
    .A2(_103_),
    .B(_109_),
    .C(_107_),
    .ZN(_011_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _253_ (.I(net52),
    .ZN(_110_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _254_ (.A1(_104_),
    .A2(_105_),
    .B(\add_u0.a[2] ),
    .ZN(_111_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _255_ (.A1(_110_),
    .A2(_103_),
    .B(_111_),
    .C(_107_),
    .ZN(_012_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _256_ (.I(net53),
    .ZN(_112_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _257_ (.A1(_104_),
    .A2(_105_),
    .B(\add_u0.a[3] ),
    .ZN(_113_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _258_ (.A1(_112_),
    .A2(_103_),
    .B(_113_),
    .C(_107_),
    .ZN(_013_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _259_ (.I(net54),
    .ZN(_114_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _260_ (.A1(_104_),
    .A2(_105_),
    .B(\add_u0.a[4] ),
    .ZN(_115_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _261_ (.A1(_114_),
    .A2(_103_),
    .B(_115_),
    .C(_107_),
    .ZN(_014_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _262_ (.I(net55),
    .ZN(_116_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _263_ (.A1(_104_),
    .A2(_105_),
    .B(\add_u0.a[5] ),
    .ZN(_117_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _264_ (.A1(_116_),
    .A2(_103_),
    .B(_117_),
    .C(_107_),
    .ZN(_015_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _265_ (.I(net56),
    .ZN(_118_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _266_ (.A1(_104_),
    .A2(_105_),
    .B(\add_u0.a[6] ),
    .ZN(_119_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _267_ (.A1(_118_),
    .A2(_103_),
    .B(_119_),
    .C(_107_),
    .ZN(_016_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _268_ (.I(net57),
    .ZN(_120_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _269_ (.A1(_104_),
    .A2(_105_),
    .B(\add_u0.a[7] ),
    .ZN(_121_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _270_ (.A1(_120_),
    .A2(_103_),
    .B(_121_),
    .C(_107_),
    .ZN(_017_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _271_ (.I(net58),
    .ZN(_122_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _272_ (.A1(_104_),
    .A2(_105_),
    .B(\add_u0.b[0] ),
    .ZN(_123_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _273_ (.A1(_122_),
    .A2(_103_),
    .B(_123_),
    .C(_107_),
    .ZN(_018_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _274_ (.I(net59),
    .ZN(_124_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _275_ (.A1(_104_),
    .A2(_105_),
    .B(\add_u0.b[1] ),
    .ZN(_125_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _276_ (.A1(_124_),
    .A2(_103_),
    .B(_125_),
    .C(_107_),
    .ZN(_019_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _277_ (.I(net35),
    .ZN(_126_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _278_ (.A1(_104_),
    .A2(_105_),
    .B(\add_u0.b[2] ),
    .ZN(_127_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _279_ (.A1(_126_),
    .A2(_103_),
    .B(_127_),
    .C(_107_),
    .ZN(_020_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _280_ (.I(net36),
    .ZN(_128_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _281_ (.A1(_104_),
    .A2(_060_),
    .B(\add_u0.b[3] ),
    .ZN(_129_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _282_ (.A1(_128_),
    .A2(_103_),
    .B(_129_),
    .C(_107_),
    .ZN(_021_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _283_ (.I(net37),
    .ZN(_130_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _284_ (.A1(_104_),
    .A2(_060_),
    .B(\add_u0.b[4] ),
    .ZN(_131_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _285_ (.A1(_130_),
    .A2(_103_),
    .B(_131_),
    .C(_043_),
    .ZN(_022_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _286_ (.I(net38),
    .ZN(_132_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _287_ (.A1(_104_),
    .A2(_060_),
    .B(\add_u0.b[5] ),
    .ZN(_133_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _288_ (.A1(_132_),
    .A2(_103_),
    .B(_133_),
    .C(_043_),
    .ZN(_023_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _289_ (.I(net39),
    .ZN(_134_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _290_ (.A1(_104_),
    .A2(_060_),
    .B(\add_u0.b[6] ),
    .ZN(_135_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _291_ (.A1(_134_),
    .A2(_103_),
    .B(_135_),
    .C(_043_),
    .ZN(_024_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _292_ (.I(net40),
    .ZN(_136_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _293_ (.A1(_104_),
    .A2(_060_),
    .B(\add_u0.b[7] ),
    .ZN(_137_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _294_ (.A1(_136_),
    .A2(_103_),
    .B(_137_),
    .C(_043_),
    .ZN(_025_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _295_ (.I(net41),
    .ZN(_138_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _296_ (.A1(_104_),
    .A2(_060_),
    .B(\mult_add_u0.m[0] ),
    .ZN(_139_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _297_ (.A1(_138_),
    .A2(_103_),
    .B(_139_),
    .C(_043_),
    .ZN(_026_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _298_ (.I(net42),
    .ZN(_140_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _299_ (.A1(_104_),
    .A2(_060_),
    .B(\mult_add_u0.m[1] ),
    .ZN(_141_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _300_ (.A1(_140_),
    .A2(_103_),
    .B(_141_),
    .C(_043_),
    .ZN(_027_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _301_ (.I(net43),
    .ZN(_142_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _302_ (.A1(_104_),
    .A2(_060_),
    .B(\mult_add_u0.m[2] ),
    .ZN(_143_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _303_ (.A1(_142_),
    .A2(_103_),
    .B(_143_),
    .C(_043_),
    .ZN(_028_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _304_ (.I(net44),
    .ZN(_144_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _305_ (.A1(_104_),
    .A2(_060_),
    .B(\mult_add_u0.m[3] ),
    .ZN(_145_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _306_ (.A1(_144_),
    .A2(_103_),
    .B(_145_),
    .C(_043_),
    .ZN(_029_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _307_ (.I(net46),
    .ZN(_146_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _308_ (.A1(_045_),
    .A2(_060_),
    .B(\mult_add_u0.m[4] ),
    .ZN(_147_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _309_ (.A1(_146_),
    .A2(_102_),
    .B(_147_),
    .C(_043_),
    .ZN(_030_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _310_ (.I(net47),
    .ZN(_148_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _311_ (.A1(_045_),
    .A2(_060_),
    .B(\mult_add_u0.m[5] ),
    .ZN(_149_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _312_ (.A1(_148_),
    .A2(_102_),
    .B(_149_),
    .C(_043_),
    .ZN(_031_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _313_ (.I(net48),
    .ZN(_150_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _314_ (.A1(_045_),
    .A2(_060_),
    .B(\mult_add_u0.m[6] ),
    .ZN(_151_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _315_ (.A1(_150_),
    .A2(_102_),
    .B(_151_),
    .C(_043_),
    .ZN(_032_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _316_ (.I(net49),
    .ZN(_152_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _317_ (.A1(_045_),
    .A2(_060_),
    .B(\mult_add_u0.m[7] ),
    .ZN(_153_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _318_ (.A1(_152_),
    .A2(_102_),
    .B(_153_),
    .C(_043_),
    .ZN(_033_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _319_ (.A1(net60),
    .A2(_044_),
    .A3(_105_),
    .Z(_154_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _320_ (.I(_154_),
    .Z(_034_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _321_ (.I(net61),
    .ZN(_155_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _322_ (.A1(net33),
    .A2(net60),
    .A3(_155_),
    .ZN(_156_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _323_ (.A1(o_wb_data[0]),
    .A2(_156_),
    .ZN(_157_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _324_ (.A1(net33),
    .A2(net60),
    .A3(_155_),
    .Z(_158_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _325_ (.A1(\out[0] ),
    .A2(_105_),
    .A3(_158_),
    .ZN(_159_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _326_ (.A1(_157_),
    .A2(_159_),
    .B(_107_),
    .ZN(_035_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _327_ (.A1(o_wb_data[1]),
    .A2(_156_),
    .ZN(_160_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _328_ (.A1(\out[1] ),
    .A2(_105_),
    .A3(_158_),
    .ZN(_161_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _329_ (.A1(_160_),
    .A2(_161_),
    .B(_107_),
    .ZN(_036_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _330_ (.A1(o_wb_data[2]),
    .A2(_156_),
    .ZN(_162_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _331_ (.A1(\out[2] ),
    .A2(_105_),
    .A3(_158_),
    .ZN(_163_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _332_ (.A1(_162_),
    .A2(_163_),
    .B(_107_),
    .ZN(_037_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _333_ (.A1(o_wb_data[3]),
    .A2(_156_),
    .ZN(_164_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _334_ (.A1(\out[3] ),
    .A2(_105_),
    .A3(_158_),
    .ZN(_165_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _335_ (.A1(_164_),
    .A2(_165_),
    .B(_107_),
    .ZN(_038_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _336_ (.A1(o_wb_data[4]),
    .A2(_156_),
    .ZN(_166_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _337_ (.A1(\out[4] ),
    .A2(_105_),
    .A3(_158_),
    .ZN(_167_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _338_ (.A1(_166_),
    .A2(_167_),
    .B(_107_),
    .ZN(_039_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _339_ (.A1(o_wb_data[5]),
    .A2(_156_),
    .ZN(_168_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _340_ (.A1(\out[5] ),
    .A2(_105_),
    .A3(_158_),
    .ZN(_169_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _341_ (.A1(_168_),
    .A2(_169_),
    .B(_107_),
    .ZN(_040_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _342_ (.A1(o_wb_data[6]),
    .A2(_156_),
    .ZN(_170_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _343_ (.A1(\out[6] ),
    .A2(_105_),
    .A3(_158_),
    .ZN(_171_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _344_ (.A1(_170_),
    .A2(_171_),
    .B(_107_),
    .ZN(_041_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _345_ (.A1(o_wb_data[7]),
    .A2(_156_),
    .ZN(_172_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _346_ (.A1(\out[7] ),
    .A2(_105_),
    .A3(_158_),
    .ZN(_173_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _347_ (.A1(_172_),
    .A2(_173_),
    .B(_107_),
    .ZN(_042_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _348_ (.D(_000_),
    .CLK(clknet_leaf_66_clk),
    .Q(\sel[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _349_ (.D(_001_),
    .CLK(clknet_leaf_66_clk),
    .Q(\sel[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _350_ (.D(_002_),
    .CLK(clknet_leaf_3_clk),
    .Q(\out[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _351_ (.D(_003_),
    .CLK(clknet_leaf_3_clk),
    .Q(\out[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _352_ (.D(_004_),
    .CLK(clknet_leaf_10_clk),
    .Q(\out[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _353_ (.D(_005_),
    .CLK(clknet_leaf_7_clk),
    .Q(\out[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _354_ (.D(_006_),
    .CLK(clknet_leaf_4_clk),
    .Q(\out[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _355_ (.D(_007_),
    .CLK(clknet_leaf_4_clk),
    .Q(\out[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _356_ (.D(_008_),
    .CLK(clknet_leaf_6_clk),
    .Q(\out[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _357_ (.D(_009_),
    .CLK(clknet_leaf_5_clk),
    .Q(\out[7] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _358_ (.D(\sel[0] ),
    .CLK(clknet_leaf_66_clk),
    .Q(\sel_d0[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _359_ (.D(\sel[1] ),
    .CLK(clknet_leaf_65_clk),
    .Q(\sel_d0[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _360_ (.D(net142),
    .CLK(clknet_leaf_65_clk),
    .Q(\sel_d1[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _361_ (.D(\sel_d0[1] ),
    .CLK(clknet_leaf_65_clk),
    .Q(\sel_d1[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _362_ (.D(\sel_d1[0] ),
    .CLK(clknet_leaf_71_clk),
    .Q(\sel_d2[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _363_ (.D(\sel_d1[1] ),
    .CLK(clknet_leaf_64_clk),
    .Q(\sel_d2[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _364_ (.D(\sel_d2[0] ),
    .CLK(clknet_leaf_71_clk),
    .Q(\sel_d3[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _365_ (.D(\sel_d2[1] ),
    .CLK(clknet_leaf_64_clk),
    .Q(\sel_d3[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _366_ (.D(\sel_d3[0] ),
    .CLK(clknet_leaf_69_clk),
    .Q(\sel_d4[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _367_ (.D(\sel_d3[1] ),
    .CLK(clknet_leaf_64_clk),
    .Q(\sel_d4[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _368_ (.D(\sel_d4[0] ),
    .CLK(clknet_leaf_89_clk),
    .Q(\sel_d5[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _369_ (.D(\sel_d4[1] ),
    .CLK(clknet_leaf_64_clk),
    .Q(\sel_d5[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _370_ (.D(\sel_d5[0] ),
    .CLK(clknet_leaf_89_clk),
    .Q(\sel_d6[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _371_ (.D(\sel_d5[1] ),
    .CLK(clknet_leaf_84_clk),
    .Q(\sel_d6[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _372_ (.D(\sel_d6[0] ),
    .CLK(clknet_leaf_84_clk),
    .Q(\sel_d7[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _373_ (.D(\sel_d6[1] ),
    .CLK(clknet_leaf_84_clk),
    .Q(\sel_d7[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _374_ (.D(\sel_d7[0] ),
    .CLK(clknet_leaf_84_clk),
    .Q(\sel_d8[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _375_ (.D(\sel_d7[1] ),
    .CLK(clknet_leaf_83_clk),
    .Q(\sel_d8[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _376_ (.D(\add_u0.ppa_u0.S[0] ),
    .CLK(clknet_leaf_95_clk),
    .Q(\add_out_d0[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _377_ (.D(\add_u0.ppa_u0.S[1] ),
    .CLK(clknet_leaf_2_clk),
    .Q(\add_out_d0[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _378_ (.D(\add_u0.ppa_u0.S[2] ),
    .CLK(clknet_leaf_3_clk),
    .Q(\add_out_d0[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _379_ (.D(\add_u0.ppa_u0.S[3] ),
    .CLK(clknet_leaf_2_clk),
    .Q(\add_out_d0[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _380_ (.D(\add_u0.ppa_u0.S[4] ),
    .CLK(clknet_leaf_94_clk),
    .Q(\add_out_d0[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _381_ (.D(\add_u0.ppa_u0.S[5] ),
    .CLK(clknet_leaf_95_clk),
    .Q(\add_out_d0[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _382_ (.D(\add_u0.ppa_u0.S[6] ),
    .CLK(clknet_leaf_95_clk),
    .Q(\add_out_d0[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _383_ (.D(\add_u0.sum[7] ),
    .CLK(clknet_leaf_91_clk),
    .Q(\add_out_d0[7] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _384_ (.D(net149),
    .CLK(clknet_leaf_96_clk),
    .Q(\add_out_d1[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _385_ (.D(net127),
    .CLK(clknet_leaf_1_clk),
    .Q(\add_out_d1[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _386_ (.D(\add_out_d0[2] ),
    .CLK(clknet_leaf_3_clk),
    .Q(\add_out_d1[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _387_ (.D(\add_out_d0[3] ),
    .CLK(clknet_leaf_2_clk),
    .Q(\add_out_d1[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _388_ (.D(\add_out_d0[4] ),
    .CLK(clknet_leaf_2_clk),
    .Q(\add_out_d1[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _389_ (.D(net125),
    .CLK(clknet_leaf_1_clk),
    .Q(\add_out_d1[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _390_ (.D(net135),
    .CLK(clknet_leaf_0_clk),
    .Q(\add_out_d1[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _391_ (.D(\add_out_d0[7] ),
    .CLK(clknet_leaf_91_clk),
    .Q(\add_out_d1[7] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _392_ (.D(net128),
    .CLK(clknet_leaf_90_clk),
    .Q(\add_out_d2[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _393_ (.D(\add_out_d1[1] ),
    .CLK(clknet_leaf_1_clk),
    .Q(\add_out_d2[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _394_ (.D(\add_out_d1[2] ),
    .CLK(clknet_leaf_3_clk),
    .Q(\add_out_d2[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _395_ (.D(\add_out_d1[3] ),
    .CLK(clknet_leaf_2_clk),
    .Q(\add_out_d2[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _396_ (.D(net126),
    .CLK(clknet_leaf_1_clk),
    .Q(\add_out_d2[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _397_ (.D(\add_out_d1[5] ),
    .CLK(clknet_leaf_1_clk),
    .Q(\add_out_d2[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _398_ (.D(\add_out_d1[6] ),
    .CLK(clknet_leaf_0_clk),
    .Q(\add_out_d2[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _399_ (.D(net134),
    .CLK(clknet_leaf_90_clk),
    .Q(\add_out_d2[7] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _400_ (.D(\add_out_d2[0] ),
    .CLK(clknet_leaf_90_clk),
    .Q(\add_out_d3[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _401_ (.D(\add_out_d2[1] ),
    .CLK(clknet_leaf_1_clk),
    .Q(\add_out_d3[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _402_ (.D(\add_out_d2[2] ),
    .CLK(clknet_leaf_8_clk),
    .Q(\add_out_d3[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _403_ (.D(net123),
    .CLK(clknet_leaf_3_clk),
    .Q(\add_out_d3[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _404_ (.D(\add_out_d2[4] ),
    .CLK(clknet_leaf_1_clk),
    .Q(\add_out_d3[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _405_ (.D(\add_out_d2[5] ),
    .CLK(clknet_leaf_0_clk),
    .Q(\add_out_d3[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _406_ (.D(\add_out_d2[6] ),
    .CLK(clknet_leaf_0_clk),
    .Q(\add_out_d3[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _407_ (.D(\add_out_d2[7] ),
    .CLK(clknet_leaf_90_clk),
    .Q(\add_out_d3[7] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _408_ (.D(\add_out_d3[0] ),
    .CLK(clknet_leaf_83_clk),
    .Q(\add_out_d4[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _409_ (.D(\add_out_d3[1] ),
    .CLK(clknet_leaf_0_clk),
    .Q(\add_out_d4[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _410_ (.D(\add_out_d3[2] ),
    .CLK(clknet_leaf_8_clk),
    .Q(\add_out_d4[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _411_ (.D(\add_out_d3[3] ),
    .CLK(clknet_leaf_3_clk),
    .Q(\add_out_d4[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _412_ (.D(\add_out_d3[4] ),
    .CLK(clknet_leaf_1_clk),
    .Q(\add_out_d4[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _413_ (.D(net140),
    .CLK(clknet_leaf_8_clk),
    .Q(\add_out_d4[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _414_ (.D(net138),
    .CLK(clknet_leaf_9_clk),
    .Q(\add_out_d4[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _415_ (.D(\add_out_d3[7] ),
    .CLK(clknet_leaf_90_clk),
    .Q(\add_out_d4[7] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _416_ (.D(\add_out_d4[0] ),
    .CLK(clknet_leaf_83_clk),
    .Q(\add_out_d5[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _417_ (.D(net145),
    .CLK(clknet_leaf_8_clk),
    .Q(\add_out_d5[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _418_ (.D(\add_out_d4[2] ),
    .CLK(clknet_leaf_7_clk),
    .Q(\add_out_d5[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _419_ (.D(\add_out_d4[3] ),
    .CLK(clknet_leaf_5_clk),
    .Q(\add_out_d5[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _420_ (.D(\add_out_d4[4] ),
    .CLK(clknet_leaf_8_clk),
    .Q(\add_out_d5[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _421_ (.D(\add_out_d4[5] ),
    .CLK(clknet_leaf_8_clk),
    .Q(\add_out_d5[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _422_ (.D(\add_out_d4[6] ),
    .CLK(clknet_leaf_9_clk),
    .Q(\add_out_d5[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _423_ (.D(\add_out_d4[7] ),
    .CLK(clknet_leaf_90_clk),
    .Q(\add_out_d5[7] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _424_ (.D(\add_out_d5[0] ),
    .CLK(clknet_leaf_83_clk),
    .Q(\add_out_d6[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _425_ (.D(\add_out_d5[1] ),
    .CLK(clknet_leaf_8_clk),
    .Q(\add_out_d6[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _426_ (.D(\add_out_d5[2] ),
    .CLK(clknet_leaf_7_clk),
    .Q(\add_out_d6[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _427_ (.D(\add_out_d5[3] ),
    .CLK(clknet_leaf_5_clk),
    .Q(\add_out_d6[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _428_ (.D(\add_out_d5[4] ),
    .CLK(clknet_leaf_8_clk),
    .Q(\add_out_d6[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _429_ (.D(net148),
    .CLK(clknet_leaf_9_clk),
    .Q(\add_out_d6[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _430_ (.D(\add_out_d5[6] ),
    .CLK(clknet_leaf_9_clk),
    .Q(\add_out_d6[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _431_ (.D(\add_out_d5[7] ),
    .CLK(clknet_leaf_83_clk),
    .Q(\add_out_d6[7] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _432_ (.D(\add_out_d6[0] ),
    .CLK(clknet_leaf_83_clk),
    .Q(\add_out_d7[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _433_ (.D(\add_out_d6[1] ),
    .CLK(clknet_leaf_9_clk),
    .Q(\add_out_d7[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _434_ (.D(\add_out_d6[2] ),
    .CLK(clknet_leaf_10_clk),
    .Q(\add_out_d7[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _435_ (.D(\add_out_d6[3] ),
    .CLK(clknet_leaf_7_clk),
    .Q(\add_out_d7[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _436_ (.D(\add_out_d6[4] ),
    .CLK(clknet_leaf_8_clk),
    .Q(\add_out_d7[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _437_ (.D(\add_out_d6[5] ),
    .CLK(clknet_leaf_9_clk),
    .Q(\add_out_d7[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _438_ (.D(\add_out_d6[6] ),
    .CLK(clknet_leaf_10_clk),
    .Q(\add_out_d7[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _439_ (.D(\add_out_d6[7] ),
    .CLK(clknet_leaf_83_clk),
    .Q(\add_out_d7[7] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _440_ (.D(\mult_u0.product_r[0] ),
    .CLK(clknet_leaf_10_clk),
    .Q(\mul_out_d0[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _441_ (.D(net146),
    .CLK(clknet_leaf_13_clk),
    .Q(\mul_out_d0[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _442_ (.D(\mult_u0.product_r[2] ),
    .CLK(clknet_leaf_14_clk),
    .Q(\mul_out_d0[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _443_ (.D(\mult_u0.product_r[3] ),
    .CLK(clknet_leaf_12_clk),
    .Q(\mul_out_d0[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _444_ (.D(\mult_u0.product_r[4] ),
    .CLK(clknet_leaf_11_clk),
    .Q(\mul_out_d0[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _445_ (.D(\mult_u0.product_r[5] ),
    .CLK(clknet_leaf_13_clk),
    .Q(\mul_out_d0[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _446_ (.D(\mult_u0.product_r[6] ),
    .CLK(clknet_leaf_13_clk),
    .Q(\mul_out_d0[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _447_ (.D(\mult_u0.product_r[7] ),
    .CLK(clknet_leaf_10_clk),
    .Q(\mul_out_d0[7] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _448_ (.D(_010_),
    .CLK(clknet_leaf_93_clk),
    .Q(\add_u0.a[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _449_ (.D(_011_),
    .CLK(clknet_leaf_93_clk),
    .Q(\add_u0.a[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _450_ (.D(_012_),
    .CLK(clknet_leaf_93_clk),
    .Q(\add_u0.a[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _451_ (.D(_013_),
    .CLK(clknet_leaf_92_clk),
    .Q(\add_u0.a[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _452_ (.D(_014_),
    .CLK(clknet_leaf_92_clk),
    .Q(\add_u0.a[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _453_ (.D(_015_),
    .CLK(clknet_leaf_92_clk),
    .Q(\add_u0.a[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _454_ (.D(_016_),
    .CLK(clknet_leaf_88_clk),
    .Q(\add_u0.a[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _455_ (.D(_017_),
    .CLK(clknet_leaf_88_clk),
    .Q(\add_u0.a[7] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _456_ (.D(_018_),
    .CLK(clknet_leaf_87_clk),
    .Q(\add_u0.b[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _457_ (.D(_019_),
    .CLK(clknet_leaf_86_clk),
    .Q(\add_u0.b[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _458_ (.D(_020_),
    .CLK(clknet_leaf_86_clk),
    .Q(\add_u0.b[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _459_ (.D(_021_),
    .CLK(clknet_leaf_86_clk),
    .Q(\add_u0.b[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _460_ (.D(_022_),
    .CLK(clknet_leaf_86_clk),
    .Q(\add_u0.b[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _461_ (.D(_023_),
    .CLK(clknet_leaf_86_clk),
    .Q(\add_u0.b[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _462_ (.D(_024_),
    .CLK(clknet_leaf_72_clk),
    .Q(\add_u0.b[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _463_ (.D(_025_),
    .CLK(clknet_leaf_72_clk),
    .Q(\add_u0.b[7] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _464_ (.D(_026_),
    .CLK(clknet_leaf_72_clk),
    .Q(\mult_add_u0.m[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _465_ (.D(_027_),
    .CLK(clknet_leaf_72_clk),
    .Q(\mult_add_u0.m[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _466_ (.D(_028_),
    .CLK(clknet_leaf_71_clk),
    .Q(\mult_add_u0.m[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _467_ (.D(_029_),
    .CLK(clknet_leaf_71_clk),
    .Q(\mult_add_u0.m[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _468_ (.D(_030_),
    .CLK(clknet_leaf_70_clk),
    .Q(\mult_add_u0.m[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _469_ (.D(_031_),
    .CLK(clknet_leaf_70_clk),
    .Q(\mult_add_u0.m[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _470_ (.D(_032_),
    .CLK(clknet_leaf_70_clk),
    .Q(\mult_add_u0.m[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _471_ (.D(_033_),
    .CLK(clknet_leaf_66_clk),
    .Q(\mult_add_u0.m[7] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _472_ (.D(_034_),
    .CLK(clknet_leaf_93_clk),
    .Q(o_wb_ack),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _473_ (.D(_035_),
    .CLK(clknet_leaf_94_clk),
    .Q(o_wb_data[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _474_ (.D(_036_),
    .CLK(clknet_leaf_3_clk),
    .Q(o_wb_data[1]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _475_ (.D(_037_),
    .CLK(clknet_leaf_3_clk),
    .Q(o_wb_data[2]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _476_ (.D(_038_),
    .CLK(clknet_3_2__leaf_clk),
    .Q(o_wb_data[3]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _477_ (.D(_039_),
    .CLK(clknet_leaf_4_clk),
    .Q(o_wb_data[4]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _478_ (.D(_040_),
    .CLK(clknet_leaf_4_clk),
    .Q(o_wb_data[5]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _479_ (.D(_041_),
    .CLK(clknet_leaf_3_clk),
    .Q(o_wb_data[6]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _480_ (.D(_042_),
    .CLK(clknet_leaf_3_clk),
    .Q(o_wb_data[7]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \add_u0._053_  (.A1(\add_u0.b[7] ),
    .A2(\add_u0.a[7] ),
    .Z(\add_u0._001_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 \add_u0._054_  (.I(\add_u0._001_ ),
    .Z(\add_u0.c_in ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \add_u0._055_  (.I(\add_u0.b[5] ),
    .ZN(\add_u0._002_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \add_u0._056_  (.I(\add_u0.b[4] ),
    .ZN(\add_u0._003_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 \add_u0._057_  (.A1(\add_u0._002_ ),
    .A2(\add_u0.a[5] ),
    .B1(\add_u0._003_ ),
    .B2(\add_u0.a[4] ),
    .ZN(\add_u0._004_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \add_u0._058_  (.I(\add_u0.a[3] ),
    .ZN(\add_u0._005_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \add_u0._059_  (.I(\add_u0.a[2] ),
    .ZN(\add_u0._006_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 \add_u0._060_  (.A1(\add_u0.b[3] ),
    .A2(\add_u0._005_ ),
    .B1(\add_u0.b[2] ),
    .B2(\add_u0._006_ ),
    .ZN(\add_u0._007_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \add_u0._061_  (.I(\add_u0.b[6] ),
    .ZN(\add_u0._008_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \add_u0._062_  (.A1(\add_u0.a[6] ),
    .A2(\add_u0._008_ ),
    .ZN(\add_u0._009_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \add_u0._063_  (.I(\add_u0.a[1] ),
    .ZN(\add_u0._010_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \add_u0._064_  (.A1(\add_u0.b[1] ),
    .A2(\add_u0._010_ ),
    .ZN(\add_u0._011_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \add_u0._065_  (.I(\add_u0.a[0] ),
    .ZN(\add_u0._012_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 \add_u0._066_  (.A1(\add_u0.b[1] ),
    .A2(\add_u0._010_ ),
    .B1(\add_u0.b[0] ),
    .B2(\add_u0._012_ ),
    .ZN(\add_u0._013_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \add_u0._067_  (.A1(\add_u0.b[2] ),
    .A2(\add_u0._006_ ),
    .ZN(\add_u0._014_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 \add_u0._068_  (.A1(\add_u0._011_ ),
    .A2(\add_u0._013_ ),
    .B(\add_u0._014_ ),
    .ZN(\add_u0._015_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \add_u0._069_  (.I(\add_u0.a[5] ),
    .ZN(\add_u0._016_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \add_u0._070_  (.A1(\add_u0.a[6] ),
    .A2(\add_u0.b[6] ),
    .Z(\add_u0._017_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0._071_  (.I(\add_u0._017_ ),
    .Z(\add_u0.a_in[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \add_u0._072_  (.A1(\add_u0.a[6] ),
    .A2(\add_u0.b[6] ),
    .ZN(\add_u0._018_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 \add_u0._073_  (.A1(\add_u0.b[5] ),
    .A2(\add_u0._016_ ),
    .B1(\add_u0.a_in[6] ),
    .B2(\add_u0._018_ ),
    .ZN(\add_u0._019_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \add_u0._074_  (.I(\add_u0.b[1] ),
    .ZN(\add_u0._020_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \add_u0._075_  (.A1(\add_u0._020_ ),
    .A2(\add_u0.a[1] ),
    .ZN(\add_u0._021_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \add_u0._076_  (.I(\add_u0.a[4] ),
    .ZN(\add_u0._022_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \add_u0._077_  (.I(\add_u0.b[0] ),
    .ZN(\add_u0._023_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 \add_u0._078_  (.A1(\add_u0.b[4] ),
    .A2(\add_u0._022_ ),
    .B1(\add_u0.b[3] ),
    .B2(\add_u0._005_ ),
    .C1(\add_u0._023_ ),
    .C2(\add_u0.a[0] ),
    .ZN(\add_u0._024_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 \add_u0._079_  (.A1(\add_u0._014_ ),
    .A2(\add_u0._021_ ),
    .A3(\add_u0._013_ ),
    .A4(\add_u0._024_ ),
    .Z(\add_u0._025_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 \add_u0._080_  (.A1(\add_u0._009_ ),
    .A2(\add_u0._015_ ),
    .B1(\add_u0._019_ ),
    .B2(\add_u0._025_ ),
    .ZN(\add_u0._026_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \add_u0._081_  (.I(\add_u0.b[3] ),
    .ZN(\add_u0._027_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 \add_u0._082_  (.A1(\add_u0._003_ ),
    .A2(\add_u0.a[4] ),
    .B1(\add_u0._027_ ),
    .B2(\add_u0.a[3] ),
    .ZN(\add_u0._028_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \add_u0._083_  (.A1(\add_u0._009_ ),
    .A2(\add_u0._028_ ),
    .ZN(\add_u0._029_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 \add_u0._084_  (.A1(\add_u0._007_ ),
    .A2(\add_u0._026_ ),
    .B(\add_u0._029_ ),
    .ZN(\add_u0._030_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \add_u0._085_  (.A1(\add_u0.a[6] ),
    .A2(\add_u0._008_ ),
    .B(\add_u0._019_ ),
    .ZN(\add_u0._031_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \add_u0._086_  (.A1(\add_u0._004_ ),
    .A2(\add_u0._030_ ),
    .B(\add_u0._031_ ),
    .ZN(\add_u0._032_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 \add_u0._087_  (.I(\add_u0._032_ ),
    .Z(\add_u0._033_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \add_u0._088_  (.I0(\add_u0.a[0] ),
    .I1(\add_u0.b[0] ),
    .S(\add_u0._033_ ),
    .Z(\add_u0._034_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \add_u0._089_  (.A1(\add_u0.c_in ),
    .A2(\add_u0._034_ ),
    .Z(\add_u0._035_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0._090_  (.I(\add_u0._035_ ),
    .Z(\add_u0.b_in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \add_u0._091_  (.I0(\add_u0.a[1] ),
    .I1(\add_u0.b[1] ),
    .S(\add_u0._033_ ),
    .Z(\add_u0._036_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \add_u0._092_  (.A1(\add_u0.c_in ),
    .A2(\add_u0._036_ ),
    .Z(\add_u0._037_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0._093_  (.I(\add_u0._037_ ),
    .Z(\add_u0.b_in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \add_u0._094_  (.I0(\add_u0.a[2] ),
    .I1(\add_u0.b[2] ),
    .S(\add_u0._033_ ),
    .Z(\add_u0._038_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \add_u0._095_  (.A1(\add_u0.c_in ),
    .A2(\add_u0._038_ ),
    .Z(\add_u0._039_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0._096_  (.I(\add_u0._039_ ),
    .Z(\add_u0.b_in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \add_u0._097_  (.I0(\add_u0.a[3] ),
    .I1(\add_u0.b[3] ),
    .S(\add_u0._033_ ),
    .Z(\add_u0._040_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \add_u0._098_  (.A1(\add_u0.c_in ),
    .A2(\add_u0._040_ ),
    .Z(\add_u0._041_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0._099_  (.I(\add_u0._041_ ),
    .Z(\add_u0.b_in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \add_u0._100_  (.I0(\add_u0.a[4] ),
    .I1(\add_u0.b[4] ),
    .S(\add_u0._033_ ),
    .Z(\add_u0._042_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \add_u0._101_  (.A1(\add_u0.c_in ),
    .A2(\add_u0._042_ ),
    .Z(\add_u0._043_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0._102_  (.I(\add_u0._043_ ),
    .Z(\add_u0.b_in[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \add_u0._103_  (.I0(\add_u0.a[5] ),
    .I1(\add_u0.b[5] ),
    .S(\add_u0._033_ ),
    .Z(\add_u0._044_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \add_u0._104_  (.A1(\add_u0.c_in ),
    .A2(\add_u0._044_ ),
    .Z(\add_u0._045_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0._105_  (.I(\add_u0._045_ ),
    .Z(\add_u0.b_in[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 \add_u0._106_  (.A1(\add_u0.c_in ),
    .A2(\add_u0._018_ ),
    .ZN(\add_u0._046_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0._107_  (.I(\add_u0._046_ ),
    .Z(\add_u0.b_in[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \add_u0._108_  (.I0(\add_u0.b[7] ),
    .I1(\add_u0.a[7] ),
    .S(\add_u0._033_ ),
    .Z(\add_u0._047_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0._109_  (.I(\add_u0._047_ ),
    .Z(\add_u0.sign ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \add_u0._110_  (.A1(\add_u0.a[0] ),
    .A2(\add_u0._033_ ),
    .ZN(\add_u0._048_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 \add_u0._111_  (.A1(\add_u0._023_ ),
    .A2(\add_u0._033_ ),
    .B(\add_u0._048_ ),
    .ZN(\add_u0.a_in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \add_u0._112_  (.A1(\add_u0.a[1] ),
    .A2(\add_u0._033_ ),
    .ZN(\add_u0._049_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 \add_u0._113_  (.A1(\add_u0._020_ ),
    .A2(\add_u0._033_ ),
    .B(\add_u0._049_ ),
    .ZN(\add_u0.a_in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \add_u0._114_  (.A1(\add_u0.b[2] ),
    .A2(\add_u0._033_ ),
    .ZN(\add_u0._050_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 \add_u0._115_  (.A1(\add_u0._006_ ),
    .A2(\add_u0._033_ ),
    .B(\add_u0._050_ ),
    .ZN(\add_u0.a_in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \add_u0._116_  (.A1(\add_u0.a[3] ),
    .A2(\add_u0._033_ ),
    .ZN(\add_u0._051_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 \add_u0._117_  (.A1(\add_u0._027_ ),
    .A2(\add_u0._033_ ),
    .B(\add_u0._051_ ),
    .ZN(\add_u0.a_in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \add_u0._118_  (.A1(\add_u0.a[4] ),
    .A2(\add_u0._033_ ),
    .ZN(\add_u0._052_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 \add_u0._119_  (.A1(\add_u0._003_ ),
    .A2(\add_u0._033_ ),
    .B(\add_u0._052_ ),
    .ZN(\add_u0.a_in[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \add_u0._120_  (.A1(\add_u0.a[5] ),
    .A2(\add_u0._033_ ),
    .ZN(\add_u0._000_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 \add_u0._121_  (.A1(\add_u0._002_ ),
    .A2(\add_u0._033_ ),
    .B(\add_u0._000_ ),
    .ZN(\add_u0.a_in[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0._122_  (.I(\add_u0.sign ),
    .Z(\add_u0.sum[7] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \add_u0.ppa_u0.d1_0.a2._1_  (.A1(\add_u0.c_in ),
    .A2(\add_u0.ppa_u0.d1_0.a2.in0 ),
    .Z(\add_u0.ppa_u0.d1_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.d1_0.a2._2_  (.I(\add_u0.ppa_u0.d1_0.a2._0_ ),
    .Z(\add_u0.ppa_u0.d1_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \add_u0.ppa_u0.d1_0.o2._1_  (.A1(\add_u0.ppa_u0.d1_0.g1 ),
    .A2(\add_u0.ppa_u0.d1_0.a2.out ),
    .Z(\add_u0.ppa_u0.d1_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.d1_0.o2._2_  (.I(\add_u0.ppa_u0.d1_0.o2._0_ ),
    .Z(\add_u0.ppa_u0.cg[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \add_u0.ppa_u0.d2_0.a2._1_  (.A1(\add_u0.ppa_u0.cg[0] ),
    .A2(\add_u0.ppa_u0.d2_0.a2.in0 ),
    .Z(\add_u0.ppa_u0.d2_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.d2_0.a2._2_  (.I(\add_u0.ppa_u0.d2_0.a2._0_ ),
    .Z(\add_u0.ppa_u0.d2_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \add_u0.ppa_u0.d2_0.o2._1_  (.A1(\add_u0.ppa_u0.d2_0.g1 ),
    .A2(\add_u0.ppa_u0.d2_0.a2.out ),
    .Z(\add_u0.ppa_u0.d2_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.d2_0.o2._2_  (.I(\add_u0.ppa_u0.d2_0.o2._0_ ),
    .Z(\add_u0.ppa_u0.cg[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \add_u0.ppa_u0.d3_0.a1._1_  (.A1(\add_u0.ppa_u0.d2_0.a2.in0 ),
    .A2(\add_u0.ppa_u0.d3_0.a1.in0 ),
    .Z(\add_u0.ppa_u0.d3_0.a1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.d3_0.a1._2_  (.I(\add_u0.ppa_u0.d3_0.a1._0_ ),
    .Z(\add_u0.ppa_u0.cp21 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \add_u0.ppa_u0.d3_0.a2._1_  (.A1(\add_u0.ppa_u0.d2_0.g1 ),
    .A2(\add_u0.ppa_u0.d3_0.a1.in0 ),
    .Z(\add_u0.ppa_u0.d3_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.d3_0.a2._2_  (.I(\add_u0.ppa_u0.d3_0.a2._0_ ),
    .Z(\add_u0.ppa_u0.d3_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \add_u0.ppa_u0.d3_0.o2._1_  (.A1(\add_u0.ppa_u0.d3_0.g1 ),
    .A2(\add_u0.ppa_u0.d3_0.a2.out ),
    .Z(\add_u0.ppa_u0.d3_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.d3_0.o2._2_  (.I(\add_u0.ppa_u0.d3_0.o2._0_ ),
    .Z(\add_u0.ppa_u0.cg21 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \add_u0.ppa_u0.d3_1.a2._1_  (.A1(\add_u0.ppa_u0.cg[0] ),
    .A2(\add_u0.ppa_u0.cp21 ),
    .Z(\add_u0.ppa_u0.d3_1.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.d3_1.a2._2_  (.I(\add_u0.ppa_u0.d3_1.a2._0_ ),
    .Z(\add_u0.ppa_u0.d3_1.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \add_u0.ppa_u0.d3_1.o2._1_  (.A1(\add_u0.ppa_u0.cg21 ),
    .A2(\add_u0.ppa_u0.d3_1.a2.out ),
    .Z(\add_u0.ppa_u0.d3_1.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.d3_1.o2._2_  (.I(\add_u0.ppa_u0.d3_1.o2._0_ ),
    .Z(\add_u0.ppa_u0.cg[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \add_u0.ppa_u0.d4_0.a2._1_  (.A1(\add_u0.ppa_u0.cg[2] ),
    .A2(\add_u0.ppa_u0.d4_0.a2.in0 ),
    .Z(\add_u0.ppa_u0.d4_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.d4_0.a2._2_  (.I(\add_u0.ppa_u0.d4_0.a2._0_ ),
    .Z(\add_u0.ppa_u0.d4_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \add_u0.ppa_u0.d4_0.o2._1_  (.A1(\add_u0.ppa_u0.d4_0.g1 ),
    .A2(\add_u0.ppa_u0.d4_0.a2.out ),
    .Z(\add_u0.ppa_u0.d4_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.d4_0.o2._2_  (.I(\add_u0.ppa_u0.d4_0.o2._0_ ),
    .Z(\add_u0.ppa_u0.cg[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \add_u0.ppa_u0.d5_0.a1._1_  (.A1(\add_u0.ppa_u0.d4_0.a2.in0 ),
    .A2(\add_u0.ppa_u0.d5_0.a1.in0 ),
    .Z(\add_u0.ppa_u0.d5_0.a1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.d5_0.a1._2_  (.I(\add_u0.ppa_u0.d5_0.a1._0_ ),
    .Z(\add_u0.ppa_u0.cp43 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \add_u0.ppa_u0.d5_0.a2._1_  (.A1(\add_u0.ppa_u0.d4_0.g1 ),
    .A2(\add_u0.ppa_u0.d5_0.a1.in0 ),
    .Z(\add_u0.ppa_u0.d5_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.d5_0.a2._2_  (.I(\add_u0.ppa_u0.d5_0.a2._0_ ),
    .Z(\add_u0.ppa_u0.d5_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \add_u0.ppa_u0.d5_0.o2._1_  (.A1(\add_u0.ppa_u0.d5_0.g1 ),
    .A2(\add_u0.ppa_u0.d5_0.a2.out ),
    .Z(\add_u0.ppa_u0.d5_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.d5_0.o2._2_  (.I(\add_u0.ppa_u0.d5_0.o2._0_ ),
    .Z(\add_u0.ppa_u0.cg43 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \add_u0.ppa_u0.d5_1.a2._1_  (.A1(\add_u0.ppa_u0.cg[2] ),
    .A2(\add_u0.ppa_u0.cp43 ),
    .Z(\add_u0.ppa_u0.d5_1.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.d5_1.a2._2_  (.I(\add_u0.ppa_u0.d5_1.a2._0_ ),
    .Z(\add_u0.ppa_u0.d5_1.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \add_u0.ppa_u0.d5_1.o2._1_  (.A1(\add_u0.ppa_u0.cg43 ),
    .A2(\add_u0.ppa_u0.d5_1.a2.out ),
    .Z(\add_u0.ppa_u0.d5_1.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.d5_1.o2._2_  (.I(\add_u0.ppa_u0.d5_1.o2._0_ ),
    .Z(\add_u0.ppa_u0.cg[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \add_u0.ppa_u0.d6_0.a1._1_  (.A1(\add_u0.ppa_u0.cp43 ),
    .A2(\add_u0.ppa_u0.d6_0.a1.in0 ),
    .Z(\add_u0.ppa_u0.d6_0.a1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.d6_0.a1._2_  (.I(\add_u0.ppa_u0.d6_0.a1._0_ ),
    .Z(\add_u0.ppa_u0.cp54 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \add_u0.ppa_u0.d6_0.a2._1_  (.A1(\add_u0.ppa_u0.cg43 ),
    .A2(\add_u0.ppa_u0.d6_0.a1.in0 ),
    .Z(\add_u0.ppa_u0.d6_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.d6_0.a2._2_  (.I(\add_u0.ppa_u0.d6_0.a2._0_ ),
    .Z(\add_u0.ppa_u0.d6_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \add_u0.ppa_u0.d6_0.o2._1_  (.A1(\add_u0.ppa_u0.d6_0.g1 ),
    .A2(\add_u0.ppa_u0.d6_0.a2.out ),
    .Z(\add_u0.ppa_u0.d6_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.d6_0.o2._2_  (.I(\add_u0.ppa_u0.d6_0.o2._0_ ),
    .Z(\add_u0.ppa_u0.cg54 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \add_u0.ppa_u0.d6_1.a2._1_  (.A1(\add_u0.ppa_u0.cg[2] ),
    .A2(\add_u0.ppa_u0.cp54 ),
    .Z(\add_u0.ppa_u0.d6_1.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.d6_1.a2._2_  (.I(\add_u0.ppa_u0.d6_1.a2._0_ ),
    .Z(\add_u0.ppa_u0.d6_1.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \add_u0.ppa_u0.d6_1.o2._1_  (.A1(\add_u0.ppa_u0.cg54 ),
    .A2(\add_u0.ppa_u0.d6_1.a2.out ),
    .Z(\add_u0.ppa_u0.d6_1.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.d6_1.o2._2_  (.I(\add_u0.ppa_u0.d6_1.o2._0_ ),
    .Z(\add_u0.ppa_u0.cg[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \add_u0.ppa_u0.p_0.a._1_  (.A1(\add_u0.b_in[0] ),
    .A2(\add_u0.a_in[0] ),
    .Z(\add_u0.ppa_u0.p_0.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.p_0.a._2_  (.I(\add_u0.ppa_u0.p_0.a._0_ ),
    .Z(\add_u0.ppa_u0.d1_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \add_u0.ppa_u0.p_0.o._1_  (.A1(\add_u0.b_in[0] ),
    .A2(\add_u0.a_in[0] ),
    .Z(\add_u0.ppa_u0.p_0.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.p_0.o._2_  (.I(\add_u0.ppa_u0.p_0.o._0_ ),
    .Z(\add_u0.ppa_u0.d1_0.a2.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \add_u0.ppa_u0.p_1.a._1_  (.A1(\add_u0.b_in[1] ),
    .A2(\add_u0.a_in[1] ),
    .Z(\add_u0.ppa_u0.p_1.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.p_1.a._2_  (.I(\add_u0.ppa_u0.p_1.a._0_ ),
    .Z(\add_u0.ppa_u0.d2_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \add_u0.ppa_u0.p_1.o._1_  (.A1(\add_u0.b_in[1] ),
    .A2(\add_u0.a_in[1] ),
    .Z(\add_u0.ppa_u0.p_1.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.p_1.o._2_  (.I(\add_u0.ppa_u0.p_1.o._0_ ),
    .Z(\add_u0.ppa_u0.d2_0.a2.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \add_u0.ppa_u0.p_2.a._1_  (.A1(\add_u0.b_in[2] ),
    .A2(\add_u0.a_in[2] ),
    .Z(\add_u0.ppa_u0.p_2.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.p_2.a._2_  (.I(\add_u0.ppa_u0.p_2.a._0_ ),
    .Z(\add_u0.ppa_u0.d3_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \add_u0.ppa_u0.p_2.o._1_  (.A1(\add_u0.b_in[2] ),
    .A2(\add_u0.a_in[2] ),
    .Z(\add_u0.ppa_u0.p_2.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.p_2.o._2_  (.I(\add_u0.ppa_u0.p_2.o._0_ ),
    .Z(\add_u0.ppa_u0.d3_0.a1.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \add_u0.ppa_u0.p_3.a._1_  (.A1(\add_u0.b_in[3] ),
    .A2(\add_u0.a_in[3] ),
    .Z(\add_u0.ppa_u0.p_3.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.p_3.a._2_  (.I(\add_u0.ppa_u0.p_3.a._0_ ),
    .Z(\add_u0.ppa_u0.d4_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \add_u0.ppa_u0.p_3.o._1_  (.A1(\add_u0.b_in[3] ),
    .A2(\add_u0.a_in[3] ),
    .Z(\add_u0.ppa_u0.p_3.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.p_3.o._2_  (.I(\add_u0.ppa_u0.p_3.o._0_ ),
    .Z(\add_u0.ppa_u0.d4_0.a2.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \add_u0.ppa_u0.p_4.a._1_  (.A1(\add_u0.b_in[4] ),
    .A2(\add_u0.a_in[4] ),
    .Z(\add_u0.ppa_u0.p_4.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.p_4.a._2_  (.I(\add_u0.ppa_u0.p_4.a._0_ ),
    .Z(\add_u0.ppa_u0.d5_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \add_u0.ppa_u0.p_4.o._1_  (.A1(\add_u0.b_in[4] ),
    .A2(\add_u0.a_in[4] ),
    .Z(\add_u0.ppa_u0.p_4.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.p_4.o._2_  (.I(\add_u0.ppa_u0.p_4.o._0_ ),
    .Z(\add_u0.ppa_u0.d5_0.a1.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \add_u0.ppa_u0.p_5.a._1_  (.A1(\add_u0.b_in[5] ),
    .A2(\add_u0.a_in[5] ),
    .Z(\add_u0.ppa_u0.p_5.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.p_5.a._2_  (.I(\add_u0.ppa_u0.p_5.a._0_ ),
    .Z(\add_u0.ppa_u0.d6_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \add_u0.ppa_u0.p_5.o._1_  (.A1(\add_u0.b_in[5] ),
    .A2(\add_u0.a_in[5] ),
    .Z(\add_u0.ppa_u0.p_5.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.p_5.o._2_  (.I(\add_u0.ppa_u0.p_5.o._0_ ),
    .Z(\add_u0.ppa_u0.d6_0.a1.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \add_u0.ppa_u0.s0.xor2_0._1_  (.A1(\add_u0.b_in[0] ),
    .A2(\add_u0.a_in[0] ),
    .Z(\add_u0.ppa_u0.s0.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.s0.xor2_0._2_  (.I(\add_u0.ppa_u0.s0.xor2_0._0_ ),
    .Z(\add_u0.ppa_u0.s0.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \add_u0.ppa_u0.s0.xor2_1._1_  (.A1(\add_u0.ppa_u0.s0.temp ),
    .A2(\add_u0.c_in ),
    .Z(\add_u0.ppa_u0.s0.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.s0.xor2_1._2_  (.I(\add_u0.ppa_u0.s0.xor2_1._0_ ),
    .Z(\add_u0.ppa_u0.S[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \add_u0.ppa_u0.s1.xor2_0._1_  (.A1(\add_u0.b_in[1] ),
    .A2(\add_u0.a_in[1] ),
    .Z(\add_u0.ppa_u0.s1.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.s1.xor2_0._2_  (.I(\add_u0.ppa_u0.s1.xor2_0._0_ ),
    .Z(\add_u0.ppa_u0.s1.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \add_u0.ppa_u0.s1.xor2_1._1_  (.A1(\add_u0.ppa_u0.s1.temp ),
    .A2(\add_u0.ppa_u0.cg[0] ),
    .Z(\add_u0.ppa_u0.s1.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.s1.xor2_1._2_  (.I(\add_u0.ppa_u0.s1.xor2_1._0_ ),
    .Z(\add_u0.ppa_u0.S[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \add_u0.ppa_u0.s2.xor2_0._1_  (.A1(\add_u0.b_in[2] ),
    .A2(\add_u0.a_in[2] ),
    .Z(\add_u0.ppa_u0.s2.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.s2.xor2_0._2_  (.I(\add_u0.ppa_u0.s2.xor2_0._0_ ),
    .Z(\add_u0.ppa_u0.s2.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \add_u0.ppa_u0.s2.xor2_1._1_  (.A1(\add_u0.ppa_u0.s2.temp ),
    .A2(\add_u0.ppa_u0.cg[1] ),
    .Z(\add_u0.ppa_u0.s2.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.s2.xor2_1._2_  (.I(\add_u0.ppa_u0.s2.xor2_1._0_ ),
    .Z(\add_u0.ppa_u0.S[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \add_u0.ppa_u0.s3.xor2_0._1_  (.A1(\add_u0.b_in[3] ),
    .A2(\add_u0.a_in[3] ),
    .Z(\add_u0.ppa_u0.s3.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.s3.xor2_0._2_  (.I(\add_u0.ppa_u0.s3.xor2_0._0_ ),
    .Z(\add_u0.ppa_u0.s3.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \add_u0.ppa_u0.s3.xor2_1._1_  (.A1(\add_u0.ppa_u0.s3.temp ),
    .A2(\add_u0.ppa_u0.cg[2] ),
    .Z(\add_u0.ppa_u0.s3.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.s3.xor2_1._2_  (.I(\add_u0.ppa_u0.s3.xor2_1._0_ ),
    .Z(\add_u0.ppa_u0.S[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \add_u0.ppa_u0.s4.xor2_0._1_  (.A1(\add_u0.b_in[4] ),
    .A2(\add_u0.a_in[4] ),
    .Z(\add_u0.ppa_u0.s4.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.s4.xor2_0._2_  (.I(\add_u0.ppa_u0.s4.xor2_0._0_ ),
    .Z(\add_u0.ppa_u0.s4.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \add_u0.ppa_u0.s4.xor2_1._1_  (.A1(\add_u0.ppa_u0.s4.temp ),
    .A2(\add_u0.ppa_u0.cg[3] ),
    .Z(\add_u0.ppa_u0.s4.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.s4.xor2_1._2_  (.I(\add_u0.ppa_u0.s4.xor2_1._0_ ),
    .Z(\add_u0.ppa_u0.S[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \add_u0.ppa_u0.s5.xor2_0._1_  (.A1(\add_u0.b_in[5] ),
    .A2(\add_u0.a_in[5] ),
    .Z(\add_u0.ppa_u0.s5.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.s5.xor2_0._2_  (.I(\add_u0.ppa_u0.s5.xor2_0._0_ ),
    .Z(\add_u0.ppa_u0.s5.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \add_u0.ppa_u0.s5.xor2_1._1_  (.A1(\add_u0.ppa_u0.s5.temp ),
    .A2(\add_u0.ppa_u0.cg[4] ),
    .Z(\add_u0.ppa_u0.s5.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.s5.xor2_1._2_  (.I(\add_u0.ppa_u0.s5.xor2_1._0_ ),
    .Z(\add_u0.ppa_u0.S[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \add_u0.ppa_u0.s6.xor2_0._1_  (.A1(\add_u0.b_in[6] ),
    .A2(\add_u0.a_in[6] ),
    .Z(\add_u0.ppa_u0.s6.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.s6.xor2_0._2_  (.I(\add_u0.ppa_u0.s6.xor2_0._0_ ),
    .Z(\add_u0.ppa_u0.s6.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \add_u0.ppa_u0.s6.xor2_1._1_  (.A1(\add_u0.ppa_u0.s6.temp ),
    .A2(\add_u0.ppa_u0.cg[5] ),
    .Z(\add_u0.ppa_u0.s6.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \add_u0.ppa_u0.s6.xor2_1._2_  (.I(\add_u0.ppa_u0.s6.xor2_1._0_ ),
    .Z(\add_u0.ppa_u0.S[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_clk (.I(net114),
    .Z(clknet_0_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_0__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_2__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_2__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_3__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_3__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_4__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_4__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_5__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_5__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_6__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_6__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_7__f_clk (.I(clknet_0_clk),
    .Z(clknet_3_7__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_0_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_0_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_10_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_10_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_11_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_11_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_12_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_12_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_13_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_13_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_14_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_14_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_15_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_15_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_16_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_16_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_17_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_17_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_18_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_18_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_1_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_1_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_20_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_20_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_21_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_21_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_22_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_22_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_23_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_23_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_24_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_24_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_25_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_25_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_26_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_26_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_27_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_27_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_28_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_28_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_29_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_29_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_2_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_2_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_30_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_30_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_31_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_31_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_32_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_32_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_33_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_33_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_34_clk (.I(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_34_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_35_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_35_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_36_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_36_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_37_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_37_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_38_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_38_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_39_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_39_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_3_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_3_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_40_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_40_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_41_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_41_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_42_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_42_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_44_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_44_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_45_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_45_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_46_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_46_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_48_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_48_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_49_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_49_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_4_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_4_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_50_clk (.I(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_50_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_51_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_51_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_53_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_53_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_54_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_54_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_55_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_55_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_56_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_56_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_57_clk (.I(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_57_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_58_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_58_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_59_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_59_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_5_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_5_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_60_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_60_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_61_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_61_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_62_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_62_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_63_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_63_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_64_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_64_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_65_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_65_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_66_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_66_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_67_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_67_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_68_clk (.I(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_68_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_69_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_69_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_6_clk (.I(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_6_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_70_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_70_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_71_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_71_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_72_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_72_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_73_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_73_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_75_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_75_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_76_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_76_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_77_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_77_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_78_clk (.I(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_78_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_79_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_79_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_7_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_7_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_80_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_80_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_81_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_81_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_82_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_82_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_83_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_83_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_84_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_84_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_86_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_86_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_87_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_87_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_88_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_88_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_89_clk (.I(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_89_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_8_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_8_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_90_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_90_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_91_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_91_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_92_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_92_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_93_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_93_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_94_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_94_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_95_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_95_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_96_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_96_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_9_clk (.I(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_9_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel core_alu_63 (.ZN(net63),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold1 (.I(\mult_add_u0.b_in_d4[7] ),
    .Z(net115),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold10 (.I(\mult_add_u0.b_in_d5[3] ),
    .Z(net124),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold11 (.I(\add_out_d0[5] ),
    .Z(net125),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold12 (.I(\add_out_d1[4] ),
    .Z(net126),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold13 (.I(\add_out_d0[1] ),
    .Z(net127),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold14 (.I(\add_out_d1[0] ),
    .Z(net128),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold15 (.I(\mult_add_u0.b_in_d2[0] ),
    .Z(net129),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold16 (.I(\mult_add_u0.b_in_d1[2] ),
    .Z(net130),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold17 (.I(\mult_add_u0.b_in_d2[1] ),
    .Z(net131),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold18 (.I(\mult_add_u0.mult0.mul_sign_s4 ),
    .Z(net132),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold19 (.I(\mult_add_u0.b_in_d2[4] ),
    .Z(net133),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold2 (.I(\mult_add_u0.m[5] ),
    .Z(net116),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold20 (.I(\add_out_d1[7] ),
    .Z(net134),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold21 (.I(\add_out_d0[6] ),
    .Z(net135),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold22 (.I(\mult_add_u0.m[6] ),
    .Z(net136),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold23 (.I(\mult_add_u0.b_in_d1[7] ),
    .Z(net137),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold24 (.I(\add_out_d3[6] ),
    .Z(net138),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold25 (.I(\mult_add_u0.b_in_d1[3] ),
    .Z(net139),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold26 (.I(\add_out_d3[5] ),
    .Z(net140),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold27 (.I(\mult_add_u0.b_in_d6[4] ),
    .Z(net141),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold28 (.I(\sel_d0[0] ),
    .Z(net142),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold29 (.I(\mult_add_u0.b_in_d1[1] ),
    .Z(net143),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold3 (.I(\mult_add_u0.b_in_d4[1] ),
    .Z(net117),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold30 (.I(\mult_add_u0.b_in_d5[6] ),
    .Z(net144),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold31 (.I(\add_out_d4[1] ),
    .Z(net145),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold32 (.I(\mult_u0.product_r[1] ),
    .Z(net146),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold33 (.I(\mult_u0.mul_sign_s4 ),
    .Z(net147),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold34 (.I(\add_out_d5[5] ),
    .Z(net148),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold35 (.I(\add_out_d0[0] ),
    .Z(net149),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold36 (.I(\mult_add_u0.b_in_d5[7] ),
    .Z(net150),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold4 (.I(\mult_add_u0.b_in_d6[7] ),
    .Z(net118),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold5 (.I(\mult_add_u0.b_in_d5[0] ),
    .Z(net119),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold6 (.I(\mult_add_u0.b_in_d1[6] ),
    .Z(net120),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold7 (.I(\mult_u0.multiplicand[0] ),
    .Z(net121),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold8 (.I(\mult_add_u0.m[4] ),
    .Z(net122),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 hold9 (.I(\add_out_d2[3] ),
    .Z(net123),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1 (.I(i_wb_addr[0]),
    .Z(net1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input10 (.I(i_wb_addr[18]),
    .Z(net10),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input11 (.I(i_wb_addr[19]),
    .Z(net11),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input12 (.I(i_wb_addr[1]),
    .Z(net12),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input13 (.I(i_wb_addr[20]),
    .Z(net13),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input14 (.I(i_wb_addr[21]),
    .Z(net14),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input15 (.I(i_wb_addr[22]),
    .Z(net15),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input16 (.I(i_wb_addr[23]),
    .Z(net16),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input17 (.I(i_wb_addr[24]),
    .Z(net17),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input18 (.I(i_wb_addr[25]),
    .Z(net18),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input19 (.I(i_wb_addr[26]),
    .Z(net19),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input2 (.I(i_wb_addr[10]),
    .Z(net2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input20 (.I(i_wb_addr[27]),
    .Z(net20),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input21 (.I(i_wb_addr[28]),
    .Z(net21),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input22 (.I(i_wb_addr[29]),
    .Z(net22),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input23 (.I(i_wb_addr[2]),
    .Z(net23),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input24 (.I(i_wb_addr[30]),
    .Z(net24),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input25 (.I(i_wb_addr[31]),
    .Z(net25),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input26 (.I(i_wb_addr[3]),
    .Z(net26),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input27 (.I(i_wb_addr[4]),
    .Z(net27),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input28 (.I(i_wb_addr[5]),
    .Z(net28),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input29 (.I(i_wb_addr[6]),
    .Z(net29),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(i_wb_addr[11]),
    .Z(net3),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input30 (.I(i_wb_addr[7]),
    .Z(net30),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input31 (.I(i_wb_addr[8]),
    .Z(net31),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input32 (.I(i_wb_addr[9]),
    .Z(net32),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input33 (.I(i_wb_cyc),
    .Z(net33),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input34 (.I(i_wb_data[0]),
    .Z(net34),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input35 (.I(i_wb_data[10]),
    .Z(net35),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input36 (.I(i_wb_data[11]),
    .Z(net36),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input37 (.I(i_wb_data[12]),
    .Z(net37),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input38 (.I(i_wb_data[13]),
    .Z(net38),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input39 (.I(i_wb_data[14]),
    .Z(net39),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input4 (.I(i_wb_addr[12]),
    .Z(net4),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input40 (.I(i_wb_data[15]),
    .Z(net40),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input41 (.I(i_wb_data[16]),
    .Z(net41),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input42 (.I(i_wb_data[17]),
    .Z(net42),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input43 (.I(i_wb_data[18]),
    .Z(net43),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input44 (.I(i_wb_data[19]),
    .Z(net44),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input45 (.I(i_wb_data[1]),
    .Z(net45),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input46 (.I(i_wb_data[20]),
    .Z(net46),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input47 (.I(i_wb_data[21]),
    .Z(net47),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input48 (.I(i_wb_data[22]),
    .Z(net48),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input49 (.I(i_wb_data[23]),
    .Z(net49),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(i_wb_addr[13]),
    .Z(net5),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input50 (.I(i_wb_data[24]),
    .Z(net50),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input51 (.I(i_wb_data[25]),
    .Z(net51),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input52 (.I(i_wb_data[2]),
    .Z(net52),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input53 (.I(i_wb_data[3]),
    .Z(net53),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input54 (.I(i_wb_data[4]),
    .Z(net54),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input55 (.I(i_wb_data[5]),
    .Z(net55),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input56 (.I(i_wb_data[6]),
    .Z(net56),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input57 (.I(i_wb_data[7]),
    .Z(net57),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input58 (.I(i_wb_data[8]),
    .Z(net58),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input59 (.I(i_wb_data[9]),
    .Z(net59),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input6 (.I(i_wb_addr[14]),
    .Z(net6),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input60 (.I(i_wb_stb),
    .Z(net60),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input61 (.I(i_wb_we),
    .Z(net61),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input62 (.I(reset),
    .Z(net62),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(i_wb_addr[15]),
    .Z(net7),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(i_wb_addr[16]),
    .Z(net8),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input9 (.I(i_wb_addr[17]),
    .Z(net9),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \mult_add_u0._017_  (.I(\mult_add_u0.add0.ppa_u0.S[0] ),
    .ZN(\mult_add_u0._008_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 \mult_add_u0._018_  (.I(net62),
    .Z(\mult_add_u0._009_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \mult_add_u0._019_  (.A1(\mult_add_u0._008_ ),
    .A2(\mult_add_u0._009_ ),
    .ZN(\mult_add_u0._000_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \mult_add_u0._020_  (.I(\mult_add_u0.add0.ppa_u0.S[1] ),
    .ZN(\mult_add_u0._010_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \mult_add_u0._021_  (.A1(\mult_add_u0._009_ ),
    .A2(\mult_add_u0._010_ ),
    .ZN(\mult_add_u0._001_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \mult_add_u0._022_  (.I(\mult_add_u0.add0.ppa_u0.S[2] ),
    .ZN(\mult_add_u0._011_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \mult_add_u0._023_  (.A1(\mult_add_u0._009_ ),
    .A2(\mult_add_u0._011_ ),
    .ZN(\mult_add_u0._002_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \mult_add_u0._024_  (.I(\mult_add_u0.add0.ppa_u0.S[3] ),
    .ZN(\mult_add_u0._012_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \mult_add_u0._025_  (.A1(\mult_add_u0._009_ ),
    .A2(\mult_add_u0._012_ ),
    .ZN(\mult_add_u0._003_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \mult_add_u0._026_  (.I(\mult_add_u0.add0.ppa_u0.S[4] ),
    .ZN(\mult_add_u0._013_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \mult_add_u0._027_  (.A1(\mult_add_u0._009_ ),
    .A2(\mult_add_u0._013_ ),
    .ZN(\mult_add_u0._004_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \mult_add_u0._028_  (.I(\mult_add_u0.add0.ppa_u0.S[5] ),
    .ZN(\mult_add_u0._014_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \mult_add_u0._029_  (.A1(\mult_add_u0._009_ ),
    .A2(\mult_add_u0._014_ ),
    .ZN(\mult_add_u0._005_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \mult_add_u0._030_  (.I(\mult_add_u0.add0.ppa_u0.S[6] ),
    .ZN(\mult_add_u0._015_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \mult_add_u0._031_  (.A1(\mult_add_u0._009_ ),
    .A2(\mult_add_u0._015_ ),
    .ZN(\mult_add_u0._006_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \mult_add_u0._032_  (.I(\mult_add_u0.add0.sum[7] ),
    .ZN(\mult_add_u0._016_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \mult_add_u0._033_  (.A1(\mult_add_u0._009_ ),
    .A2(\mult_add_u0._016_ ),
    .ZN(\mult_add_u0._007_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._034_  (.D(\add_u0.b[0] ),
    .CLK(clknet_leaf_82_clk),
    .Q(\mult_add_u0.b_in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._035_  (.D(\add_u0.b[1] ),
    .CLK(clknet_leaf_82_clk),
    .Q(\mult_add_u0.b_in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._036_  (.D(\add_u0.b[2] ),
    .CLK(clknet_leaf_14_clk),
    .Q(\mult_add_u0.b_in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._037_  (.D(\add_u0.b[3] ),
    .CLK(clknet_leaf_80_clk),
    .Q(\mult_add_u0.b_in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._038_  (.D(\add_u0.b[4] ),
    .CLK(clknet_leaf_33_clk),
    .Q(\mult_add_u0.b_in[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._039_  (.D(\add_u0.b[5] ),
    .CLK(clknet_leaf_33_clk),
    .Q(\mult_add_u0.b_in[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._040_  (.D(\add_u0.b[6] ),
    .CLK(clknet_leaf_79_clk),
    .Q(\mult_add_u0.b_in[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._041_  (.D(\add_u0.b[7] ),
    .CLK(clknet_leaf_88_clk),
    .Q(\mult_add_u0.b_in[7] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._042_  (.D(\mult_add_u0.b_in[0] ),
    .CLK(clknet_leaf_82_clk),
    .Q(\mult_add_u0.b_in_d1[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._043_  (.D(\mult_add_u0.b_in[1] ),
    .CLK(clknet_leaf_82_clk),
    .Q(\mult_add_u0.b_in_d1[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._044_  (.D(\mult_add_u0.b_in[2] ),
    .CLK(clknet_leaf_15_clk),
    .Q(\mult_add_u0.b_in_d1[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._045_  (.D(\mult_add_u0.b_in[3] ),
    .CLK(clknet_leaf_10_clk),
    .Q(\mult_add_u0.b_in_d1[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._046_  (.D(\mult_add_u0.b_in[4] ),
    .CLK(clknet_leaf_35_clk),
    .Q(\mult_add_u0.b_in_d1[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._047_  (.D(\mult_add_u0.b_in[5] ),
    .CLK(clknet_leaf_33_clk),
    .Q(\mult_add_u0.b_in_d1[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._048_  (.D(\mult_add_u0.b_in[6] ),
    .CLK(clknet_leaf_79_clk),
    .Q(\mult_add_u0.b_in_d1[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._049_  (.D(\mult_add_u0.b_in[7] ),
    .CLK(clknet_leaf_88_clk),
    .Q(\mult_add_u0.b_in_d1[7] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._050_  (.D(\mult_add_u0.b_in_d1[0] ),
    .CLK(clknet_leaf_82_clk),
    .Q(\mult_add_u0.b_in_d2[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._051_  (.D(net143),
    .CLK(clknet_leaf_81_clk),
    .Q(\mult_add_u0.b_in_d2[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._052_  (.D(net130),
    .CLK(clknet_leaf_13_clk),
    .Q(\mult_add_u0.b_in_d2[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._053_  (.D(net139),
    .CLK(clknet_leaf_79_clk),
    .Q(\mult_add_u0.b_in_d2[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._054_  (.D(\mult_add_u0.b_in_d1[4] ),
    .CLK(clknet_leaf_35_clk),
    .Q(\mult_add_u0.b_in_d2[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._055_  (.D(\mult_add_u0.b_in_d1[5] ),
    .CLK(clknet_leaf_35_clk),
    .Q(\mult_add_u0.b_in_d2[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._056_  (.D(net120),
    .CLK(clknet_leaf_78_clk),
    .Q(\mult_add_u0.b_in_d2[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._057_  (.D(net137),
    .CLK(clknet_leaf_89_clk),
    .Q(\mult_add_u0.b_in_d2[7] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._058_  (.D(net129),
    .CLK(clknet_leaf_80_clk),
    .Q(\mult_add_u0.b_in_d3[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._059_  (.D(net131),
    .CLK(clknet_leaf_80_clk),
    .Q(\mult_add_u0.b_in_d3[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._060_  (.D(\mult_add_u0.b_in_d2[2] ),
    .CLK(clknet_leaf_34_clk),
    .Q(\mult_add_u0.b_in_d3[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._061_  (.D(\mult_add_u0.b_in_d2[3] ),
    .CLK(clknet_leaf_79_clk),
    .Q(\mult_add_u0.b_in_d3[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._062_  (.D(net133),
    .CLK(clknet_leaf_36_clk),
    .Q(\mult_add_u0.b_in_d3[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._063_  (.D(\mult_add_u0.b_in_d2[5] ),
    .CLK(clknet_leaf_35_clk),
    .Q(\mult_add_u0.b_in_d3[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._064_  (.D(\mult_add_u0.b_in_d2[6] ),
    .CLK(clknet_leaf_78_clk),
    .Q(\mult_add_u0.b_in_d3[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._065_  (.D(\mult_add_u0.b_in_d2[7] ),
    .CLK(clknet_leaf_87_clk),
    .Q(\mult_add_u0.b_in_d3[7] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._066_  (.D(\mult_add_u0.b_in_d3[0] ),
    .CLK(clknet_leaf_80_clk),
    .Q(\mult_add_u0.b_in_d4[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._067_  (.D(\mult_add_u0.b_in_d3[1] ),
    .CLK(clknet_leaf_80_clk),
    .Q(\mult_add_u0.b_in_d4[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._068_  (.D(\mult_add_u0.b_in_d3[2] ),
    .CLK(clknet_leaf_34_clk),
    .Q(\mult_add_u0.b_in_d4[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._069_  (.D(\mult_add_u0.b_in_d3[3] ),
    .CLK(clknet_leaf_79_clk),
    .Q(\mult_add_u0.b_in_d4[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._070_  (.D(\mult_add_u0.b_in_d3[4] ),
    .CLK(clknet_leaf_36_clk),
    .Q(\mult_add_u0.b_in_d4[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._071_  (.D(\mult_add_u0.b_in_d3[5] ),
    .CLK(clknet_leaf_35_clk),
    .Q(\mult_add_u0.b_in_d4[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._072_  (.D(\mult_add_u0.b_in_d3[6] ),
    .CLK(clknet_leaf_78_clk),
    .Q(\mult_add_u0.b_in_d4[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._073_  (.D(\mult_add_u0.b_in_d3[7] ),
    .CLK(clknet_3_1__leaf_clk),
    .Q(\mult_add_u0.b_in_d4[7] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._074_  (.D(\mult_add_u0.b_in_d4[0] ),
    .CLK(clknet_leaf_80_clk),
    .Q(\mult_add_u0.b_in_d5[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._075_  (.D(net117),
    .CLK(clknet_leaf_77_clk),
    .Q(\mult_add_u0.b_in_d5[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._076_  (.D(\mult_add_u0.b_in_d4[2] ),
    .CLK(clknet_leaf_34_clk),
    .Q(\mult_add_u0.b_in_d5[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._077_  (.D(\mult_add_u0.b_in_d4[3] ),
    .CLK(clknet_leaf_79_clk),
    .Q(\mult_add_u0.b_in_d5[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._078_  (.D(\mult_add_u0.b_in_d4[4] ),
    .CLK(clknet_leaf_37_clk),
    .Q(\mult_add_u0.b_in_d5[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._079_  (.D(\mult_add_u0.b_in_d4[5] ),
    .CLK(clknet_leaf_37_clk),
    .Q(\mult_add_u0.b_in_d5[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._080_  (.D(\mult_add_u0.b_in_d4[6] ),
    .CLK(clknet_leaf_53_clk),
    .Q(\mult_add_u0.b_in_d5[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._081_  (.D(net115),
    .CLK(clknet_leaf_81_clk),
    .Q(\mult_add_u0.b_in_d5[7] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._082_  (.D(net119),
    .CLK(clknet_leaf_78_clk),
    .Q(\mult_add_u0.b_in_d6[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._083_  (.D(\mult_add_u0.b_in_d5[1] ),
    .CLK(clknet_leaf_77_clk),
    .Q(\mult_add_u0.b_in_d6[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._084_  (.D(\mult_add_u0.b_in_d5[2] ),
    .CLK(clknet_leaf_33_clk),
    .Q(\mult_add_u0.b_in_d6[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._085_  (.D(net124),
    .CLK(clknet_leaf_78_clk),
    .Q(\mult_add_u0.b_in_d6[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._086_  (.D(\mult_add_u0.b_in_d5[4] ),
    .CLK(clknet_leaf_37_clk),
    .Q(\mult_add_u0.b_in_d6[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._087_  (.D(\mult_add_u0.b_in_d5[5] ),
    .CLK(clknet_leaf_37_clk),
    .Q(\mult_add_u0.b_in_d6[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._088_  (.D(net144),
    .CLK(clknet_leaf_55_clk),
    .Q(\mult_add_u0.b_in_d6[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._089_  (.D(net150),
    .CLK(clknet_leaf_80_clk),
    .Q(\mult_add_u0.b_in_d6[7] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._090_  (.D(\mult_add_u0.b_in_d6[0] ),
    .CLK(clknet_leaf_78_clk),
    .Q(\mult_add_u0.add0.b[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._091_  (.D(\mult_add_u0.b_in_d6[1] ),
    .CLK(clknet_leaf_77_clk),
    .Q(\mult_add_u0.add0.b[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._092_  (.D(\mult_add_u0.b_in_d6[2] ),
    .CLK(clknet_leaf_35_clk),
    .Q(\mult_add_u0.add0.b[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._093_  (.D(\mult_add_u0.b_in_d6[3] ),
    .CLK(clknet_3_6__leaf_clk),
    .Q(\mult_add_u0.add0.b[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._094_  (.D(net141),
    .CLK(clknet_leaf_50_clk),
    .Q(\mult_add_u0.add0.b[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._095_  (.D(\mult_add_u0.b_in_d6[5] ),
    .CLK(clknet_leaf_37_clk),
    .Q(\mult_add_u0.add0.b[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._096_  (.D(\mult_add_u0.b_in_d6[6] ),
    .CLK(clknet_leaf_53_clk),
    .Q(\mult_add_u0.add0.b[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._097_  (.D(net118),
    .CLK(clknet_leaf_77_clk),
    .Q(\mult_add_u0.add0.b[7] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._098_  (.D(\mult_add_u0._000_ ),
    .CLK(clknet_leaf_79_clk),
    .Q(\mult_add_u0.out[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._099_  (.D(\mult_add_u0._001_ ),
    .CLK(clknet_leaf_79_clk),
    .Q(\mult_add_u0.out[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._100_  (.D(\mult_add_u0._002_ ),
    .CLK(clknet_leaf_12_clk),
    .Q(\mult_add_u0.out[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._101_  (.D(\mult_add_u0._003_ ),
    .CLK(clknet_leaf_12_clk),
    .Q(\mult_add_u0.out[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._102_  (.D(\mult_add_u0._004_ ),
    .CLK(clknet_leaf_12_clk),
    .Q(\mult_add_u0.out[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._103_  (.D(\mult_add_u0._005_ ),
    .CLK(clknet_leaf_12_clk),
    .Q(\mult_add_u0.out[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._104_  (.D(\mult_add_u0._006_ ),
    .CLK(clknet_leaf_12_clk),
    .Q(\mult_add_u0.out[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0._105_  (.D(\mult_add_u0._007_ ),
    .CLK(clknet_leaf_79_clk),
    .Q(\mult_add_u0.out[7] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.add0._053_  (.A1(\mult_add_u0.add0.b[7] ),
    .A2(\mult_add_u0.add0.a[7] ),
    .Z(\mult_add_u0.add0._001_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 \mult_add_u0.add0._054_  (.I(\mult_add_u0.add0._001_ ),
    .Z(\mult_add_u0.add0.c_in ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \mult_add_u0.add0._055_  (.I(\mult_add_u0.add0.b[5] ),
    .ZN(\mult_add_u0.add0._002_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 \mult_add_u0.add0._056_  (.I(\mult_add_u0.add0.b[4] ),
    .ZN(\mult_add_u0.add0._003_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 \mult_add_u0.add0._057_  (.A1(\mult_add_u0.add0._002_ ),
    .A2(\mult_add_u0.add0.a[5] ),
    .B1(\mult_add_u0.add0._003_ ),
    .B2(\mult_add_u0.add0.a[4] ),
    .ZN(\mult_add_u0.add0._004_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \mult_add_u0.add0._058_  (.I(\mult_add_u0.add0.a[3] ),
    .ZN(\mult_add_u0.add0._005_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \mult_add_u0.add0._059_  (.I(\mult_add_u0.add0.a[2] ),
    .ZN(\mult_add_u0.add0._006_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 \mult_add_u0.add0._060_  (.A1(\mult_add_u0.add0.b[3] ),
    .A2(\mult_add_u0.add0._005_ ),
    .B1(\mult_add_u0.add0.b[2] ),
    .B2(\mult_add_u0.add0._006_ ),
    .ZN(\mult_add_u0.add0._007_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \mult_add_u0.add0._061_  (.I(\mult_add_u0.add0.b[6] ),
    .ZN(\mult_add_u0.add0._008_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \mult_add_u0.add0._062_  (.A1(\mult_add_u0.add0.a[6] ),
    .A2(\mult_add_u0.add0._008_ ),
    .ZN(\mult_add_u0.add0._009_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \mult_add_u0.add0._063_  (.I(\mult_add_u0.add0.a[1] ),
    .ZN(\mult_add_u0.add0._010_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \mult_add_u0.add0._064_  (.A1(\mult_add_u0.add0.b[1] ),
    .A2(\mult_add_u0.add0._010_ ),
    .ZN(\mult_add_u0.add0._011_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \mult_add_u0.add0._065_  (.I(\mult_add_u0.add0.a[0] ),
    .ZN(\mult_add_u0.add0._012_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 \mult_add_u0.add0._066_  (.A1(\mult_add_u0.add0.b[1] ),
    .A2(\mult_add_u0.add0._010_ ),
    .B1(\mult_add_u0.add0.b[0] ),
    .B2(\mult_add_u0.add0._012_ ),
    .ZN(\mult_add_u0.add0._013_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \mult_add_u0.add0._067_  (.A1(\mult_add_u0.add0.b[2] ),
    .A2(\mult_add_u0.add0._006_ ),
    .ZN(\mult_add_u0.add0._014_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 \mult_add_u0.add0._068_  (.A1(\mult_add_u0.add0._011_ ),
    .A2(\mult_add_u0.add0._013_ ),
    .B(\mult_add_u0.add0._014_ ),
    .ZN(\mult_add_u0.add0._015_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \mult_add_u0.add0._069_  (.I(\mult_add_u0.add0.a[5] ),
    .ZN(\mult_add_u0.add0._016_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.add0._070_  (.A1(\mult_add_u0.add0.a[6] ),
    .A2(\mult_add_u0.add0.b[6] ),
    .Z(\mult_add_u0.add0._017_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0._071_  (.I(\mult_add_u0.add0._017_ ),
    .Z(\mult_add_u0.add0.a_in[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \mult_add_u0.add0._072_  (.A1(\mult_add_u0.add0.a[6] ),
    .A2(\mult_add_u0.add0.b[6] ),
    .ZN(\mult_add_u0.add0._018_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 \mult_add_u0.add0._073_  (.A1(\mult_add_u0.add0.b[5] ),
    .A2(\mult_add_u0.add0._016_ ),
    .B1(\mult_add_u0.add0.a_in[6] ),
    .B2(\mult_add_u0.add0._018_ ),
    .ZN(\mult_add_u0.add0._019_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \mult_add_u0.add0._074_  (.I(\mult_add_u0.add0.b[1] ),
    .ZN(\mult_add_u0.add0._020_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \mult_add_u0.add0._075_  (.A1(\mult_add_u0.add0._020_ ),
    .A2(\mult_add_u0.add0.a[1] ),
    .ZN(\mult_add_u0.add0._021_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \mult_add_u0.add0._076_  (.I(\mult_add_u0.add0.a[4] ),
    .ZN(\mult_add_u0.add0._022_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \mult_add_u0.add0._077_  (.I(\mult_add_u0.add0.b[0] ),
    .ZN(\mult_add_u0.add0._023_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 \mult_add_u0.add0._078_  (.A1(\mult_add_u0.add0.b[4] ),
    .A2(\mult_add_u0.add0._022_ ),
    .B1(\mult_add_u0.add0.b[3] ),
    .B2(\mult_add_u0.add0._005_ ),
    .C1(\mult_add_u0.add0._023_ ),
    .C2(\mult_add_u0.add0.a[0] ),
    .ZN(\mult_add_u0.add0._024_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 \mult_add_u0.add0._079_  (.A1(\mult_add_u0.add0._014_ ),
    .A2(\mult_add_u0.add0._021_ ),
    .A3(\mult_add_u0.add0._013_ ),
    .A4(\mult_add_u0.add0._024_ ),
    .Z(\mult_add_u0.add0._025_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 \mult_add_u0.add0._080_  (.A1(\mult_add_u0.add0._009_ ),
    .A2(\mult_add_u0.add0._015_ ),
    .B1(\mult_add_u0.add0._019_ ),
    .B2(\mult_add_u0.add0._025_ ),
    .ZN(\mult_add_u0.add0._026_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \mult_add_u0.add0._081_  (.I(\mult_add_u0.add0.b[3] ),
    .ZN(\mult_add_u0.add0._027_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 \mult_add_u0.add0._082_  (.A1(\mult_add_u0.add0._003_ ),
    .A2(\mult_add_u0.add0.a[4] ),
    .B1(\mult_add_u0.add0._027_ ),
    .B2(\mult_add_u0.add0.a[3] ),
    .ZN(\mult_add_u0.add0._028_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \mult_add_u0.add0._083_  (.A1(\mult_add_u0.add0._009_ ),
    .A2(\mult_add_u0.add0._028_ ),
    .ZN(\mult_add_u0.add0._029_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 \mult_add_u0.add0._084_  (.A1(\mult_add_u0.add0._007_ ),
    .A2(\mult_add_u0.add0._026_ ),
    .B(\mult_add_u0.add0._029_ ),
    .ZN(\mult_add_u0.add0._030_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \mult_add_u0.add0._085_  (.A1(\mult_add_u0.add0.a[6] ),
    .A2(\mult_add_u0.add0._008_ ),
    .B(\mult_add_u0.add0._019_ ),
    .ZN(\mult_add_u0.add0._031_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \mult_add_u0.add0._086_  (.A1(\mult_add_u0.add0._004_ ),
    .A2(\mult_add_u0.add0._030_ ),
    .B(\mult_add_u0.add0._031_ ),
    .ZN(\mult_add_u0.add0._032_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 \mult_add_u0.add0._087_  (.I(\mult_add_u0.add0._032_ ),
    .Z(\mult_add_u0.add0._033_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.add0._088_  (.I0(\mult_add_u0.add0.a[0] ),
    .I1(\mult_add_u0.add0.b[0] ),
    .S(\mult_add_u0.add0._033_ ),
    .Z(\mult_add_u0.add0._034_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.add0._089_  (.A1(\mult_add_u0.add0.c_in ),
    .A2(\mult_add_u0.add0._034_ ),
    .Z(\mult_add_u0.add0._035_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0._090_  (.I(\mult_add_u0.add0._035_ ),
    .Z(\mult_add_u0.add0.b_in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.add0._091_  (.I0(\mult_add_u0.add0.a[1] ),
    .I1(\mult_add_u0.add0.b[1] ),
    .S(\mult_add_u0.add0._033_ ),
    .Z(\mult_add_u0.add0._036_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.add0._092_  (.A1(\mult_add_u0.add0.c_in ),
    .A2(\mult_add_u0.add0._036_ ),
    .Z(\mult_add_u0.add0._037_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0._093_  (.I(\mult_add_u0.add0._037_ ),
    .Z(\mult_add_u0.add0.b_in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.add0._094_  (.I0(\mult_add_u0.add0.a[2] ),
    .I1(\mult_add_u0.add0.b[2] ),
    .S(\mult_add_u0.add0._033_ ),
    .Z(\mult_add_u0.add0._038_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.add0._095_  (.A1(\mult_add_u0.add0.c_in ),
    .A2(\mult_add_u0.add0._038_ ),
    .Z(\mult_add_u0.add0._039_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0._096_  (.I(\mult_add_u0.add0._039_ ),
    .Z(\mult_add_u0.add0.b_in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.add0._097_  (.I0(\mult_add_u0.add0.a[3] ),
    .I1(\mult_add_u0.add0.b[3] ),
    .S(\mult_add_u0.add0._033_ ),
    .Z(\mult_add_u0.add0._040_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.add0._098_  (.A1(\mult_add_u0.add0.c_in ),
    .A2(\mult_add_u0.add0._040_ ),
    .Z(\mult_add_u0.add0._041_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0._099_  (.I(\mult_add_u0.add0._041_ ),
    .Z(\mult_add_u0.add0.b_in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.add0._100_  (.I0(\mult_add_u0.add0.a[4] ),
    .I1(\mult_add_u0.add0.b[4] ),
    .S(\mult_add_u0.add0._033_ ),
    .Z(\mult_add_u0.add0._042_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.add0._101_  (.A1(\mult_add_u0.add0.c_in ),
    .A2(\mult_add_u0.add0._042_ ),
    .Z(\mult_add_u0.add0._043_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0._102_  (.I(\mult_add_u0.add0._043_ ),
    .Z(\mult_add_u0.add0.b_in[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.add0._103_  (.I0(\mult_add_u0.add0.a[5] ),
    .I1(\mult_add_u0.add0.b[5] ),
    .S(\mult_add_u0.add0._033_ ),
    .Z(\mult_add_u0.add0._044_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.add0._104_  (.A1(\mult_add_u0.add0.c_in ),
    .A2(\mult_add_u0.add0._044_ ),
    .Z(\mult_add_u0.add0._045_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0._105_  (.I(\mult_add_u0.add0._045_ ),
    .Z(\mult_add_u0.add0.b_in[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 \mult_add_u0.add0._106_  (.A1(\mult_add_u0.add0.c_in ),
    .A2(\mult_add_u0.add0._018_ ),
    .ZN(\mult_add_u0.add0._046_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0._107_  (.I(\mult_add_u0.add0._046_ ),
    .Z(\mult_add_u0.add0.b_in[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.add0._108_  (.I0(\mult_add_u0.add0.b[7] ),
    .I1(\mult_add_u0.add0.a[7] ),
    .S(\mult_add_u0.add0._033_ ),
    .Z(\mult_add_u0.add0._047_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0._109_  (.I(\mult_add_u0.add0._047_ ),
    .Z(\mult_add_u0.add0.sign ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \mult_add_u0.add0._110_  (.A1(\mult_add_u0.add0.a[0] ),
    .A2(\mult_add_u0.add0._033_ ),
    .ZN(\mult_add_u0.add0._048_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 \mult_add_u0.add0._111_  (.A1(\mult_add_u0.add0._023_ ),
    .A2(\mult_add_u0.add0._033_ ),
    .B(\mult_add_u0.add0._048_ ),
    .ZN(\mult_add_u0.add0.a_in[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \mult_add_u0.add0._112_  (.A1(\mult_add_u0.add0.a[1] ),
    .A2(\mult_add_u0.add0._033_ ),
    .ZN(\mult_add_u0.add0._049_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 \mult_add_u0.add0._113_  (.A1(\mult_add_u0.add0._020_ ),
    .A2(\mult_add_u0.add0._033_ ),
    .B(\mult_add_u0.add0._049_ ),
    .ZN(\mult_add_u0.add0.a_in[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \mult_add_u0.add0._114_  (.A1(\mult_add_u0.add0.b[2] ),
    .A2(\mult_add_u0.add0._033_ ),
    .ZN(\mult_add_u0.add0._050_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 \mult_add_u0.add0._115_  (.A1(\mult_add_u0.add0._006_ ),
    .A2(\mult_add_u0.add0._033_ ),
    .B(\mult_add_u0.add0._050_ ),
    .ZN(\mult_add_u0.add0.a_in[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \mult_add_u0.add0._116_  (.A1(\mult_add_u0.add0.a[3] ),
    .A2(\mult_add_u0.add0._033_ ),
    .ZN(\mult_add_u0.add0._051_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 \mult_add_u0.add0._117_  (.A1(\mult_add_u0.add0._027_ ),
    .A2(\mult_add_u0.add0._033_ ),
    .B(\mult_add_u0.add0._051_ ),
    .ZN(\mult_add_u0.add0.a_in[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \mult_add_u0.add0._118_  (.A1(\mult_add_u0.add0.a[4] ),
    .A2(\mult_add_u0.add0._033_ ),
    .ZN(\mult_add_u0.add0._052_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 \mult_add_u0.add0._119_  (.A1(\mult_add_u0.add0._003_ ),
    .A2(\mult_add_u0.add0._033_ ),
    .B(\mult_add_u0.add0._052_ ),
    .ZN(\mult_add_u0.add0.a_in[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \mult_add_u0.add0._120_  (.A1(\mult_add_u0.add0.a[5] ),
    .A2(\mult_add_u0.add0._033_ ),
    .ZN(\mult_add_u0.add0._000_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 \mult_add_u0.add0._121_  (.A1(\mult_add_u0.add0._002_ ),
    .A2(\mult_add_u0.add0._033_ ),
    .B(\mult_add_u0.add0._000_ ),
    .ZN(\mult_add_u0.add0.a_in[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0._122_  (.I(\mult_add_u0.add0.sign ),
    .Z(\mult_add_u0.add0.sum[7] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.add0.ppa_u0.d1_0.a2._1_  (.A1(\mult_add_u0.add0.c_in ),
    .A2(\mult_add_u0.add0.ppa_u0.d1_0.a2.in0 ),
    .Z(\mult_add_u0.add0.ppa_u0.d1_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0.ppa_u0.d1_0.a2._2_  (.I(\mult_add_u0.add0.ppa_u0.d1_0.a2._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.d1_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.add0.ppa_u0.d1_0.o2._1_  (.A1(\mult_add_u0.add0.ppa_u0.d1_0.g1 ),
    .A2(\mult_add_u0.add0.ppa_u0.d1_0.a2.out ),
    .Z(\mult_add_u0.add0.ppa_u0.d1_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0.ppa_u0.d1_0.o2._2_  (.I(\mult_add_u0.add0.ppa_u0.d1_0.o2._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.cg[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.add0.ppa_u0.d2_0.a2._1_  (.A1(\mult_add_u0.add0.ppa_u0.cg[0] ),
    .A2(\mult_add_u0.add0.ppa_u0.d2_0.a2.in0 ),
    .Z(\mult_add_u0.add0.ppa_u0.d2_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0.ppa_u0.d2_0.a2._2_  (.I(\mult_add_u0.add0.ppa_u0.d2_0.a2._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.d2_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.add0.ppa_u0.d2_0.o2._1_  (.A1(\mult_add_u0.add0.ppa_u0.d2_0.g1 ),
    .A2(\mult_add_u0.add0.ppa_u0.d2_0.a2.out ),
    .Z(\mult_add_u0.add0.ppa_u0.d2_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0.ppa_u0.d2_0.o2._2_  (.I(\mult_add_u0.add0.ppa_u0.d2_0.o2._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.cg[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.add0.ppa_u0.d3_0.a1._1_  (.A1(\mult_add_u0.add0.ppa_u0.d2_0.a2.in0 ),
    .A2(\mult_add_u0.add0.ppa_u0.d3_0.a1.in0 ),
    .Z(\mult_add_u0.add0.ppa_u0.d3_0.a1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0.ppa_u0.d3_0.a1._2_  (.I(\mult_add_u0.add0.ppa_u0.d3_0.a1._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.cp21 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.add0.ppa_u0.d3_0.a2._1_  (.A1(\mult_add_u0.add0.ppa_u0.d2_0.g1 ),
    .A2(\mult_add_u0.add0.ppa_u0.d3_0.a1.in0 ),
    .Z(\mult_add_u0.add0.ppa_u0.d3_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0.ppa_u0.d3_0.a2._2_  (.I(\mult_add_u0.add0.ppa_u0.d3_0.a2._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.d3_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.add0.ppa_u0.d3_0.o2._1_  (.A1(\mult_add_u0.add0.ppa_u0.d3_0.g1 ),
    .A2(\mult_add_u0.add0.ppa_u0.d3_0.a2.out ),
    .Z(\mult_add_u0.add0.ppa_u0.d3_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0.ppa_u0.d3_0.o2._2_  (.I(\mult_add_u0.add0.ppa_u0.d3_0.o2._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.cg21 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.add0.ppa_u0.d3_1.a2._1_  (.A1(\mult_add_u0.add0.ppa_u0.cg[0] ),
    .A2(\mult_add_u0.add0.ppa_u0.cp21 ),
    .Z(\mult_add_u0.add0.ppa_u0.d3_1.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0.ppa_u0.d3_1.a2._2_  (.I(\mult_add_u0.add0.ppa_u0.d3_1.a2._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.d3_1.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.add0.ppa_u0.d3_1.o2._1_  (.A1(\mult_add_u0.add0.ppa_u0.cg21 ),
    .A2(\mult_add_u0.add0.ppa_u0.d3_1.a2.out ),
    .Z(\mult_add_u0.add0.ppa_u0.d3_1.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 \mult_add_u0.add0.ppa_u0.d3_1.o2._2_  (.I(\mult_add_u0.add0.ppa_u0.d3_1.o2._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.cg[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.add0.ppa_u0.d4_0.a2._1_  (.A1(\mult_add_u0.add0.ppa_u0.cg[2] ),
    .A2(\mult_add_u0.add0.ppa_u0.d4_0.a2.in0 ),
    .Z(\mult_add_u0.add0.ppa_u0.d4_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0.ppa_u0.d4_0.a2._2_  (.I(\mult_add_u0.add0.ppa_u0.d4_0.a2._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.d4_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.add0.ppa_u0.d4_0.o2._1_  (.A1(\mult_add_u0.add0.ppa_u0.d4_0.g1 ),
    .A2(\mult_add_u0.add0.ppa_u0.d4_0.a2.out ),
    .Z(\mult_add_u0.add0.ppa_u0.d4_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0.ppa_u0.d4_0.o2._2_  (.I(\mult_add_u0.add0.ppa_u0.d4_0.o2._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.cg[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.add0.ppa_u0.d5_0.a1._1_  (.A1(\mult_add_u0.add0.ppa_u0.d4_0.a2.in0 ),
    .A2(\mult_add_u0.add0.ppa_u0.d5_0.a1.in0 ),
    .Z(\mult_add_u0.add0.ppa_u0.d5_0.a1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0.ppa_u0.d5_0.a1._2_  (.I(\mult_add_u0.add0.ppa_u0.d5_0.a1._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.cp43 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.add0.ppa_u0.d5_0.a2._1_  (.A1(\mult_add_u0.add0.ppa_u0.d4_0.g1 ),
    .A2(\mult_add_u0.add0.ppa_u0.d5_0.a1.in0 ),
    .Z(\mult_add_u0.add0.ppa_u0.d5_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0.ppa_u0.d5_0.a2._2_  (.I(\mult_add_u0.add0.ppa_u0.d5_0.a2._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.d5_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.add0.ppa_u0.d5_0.o2._1_  (.A1(\mult_add_u0.add0.ppa_u0.d5_0.g1 ),
    .A2(\mult_add_u0.add0.ppa_u0.d5_0.a2.out ),
    .Z(\mult_add_u0.add0.ppa_u0.d5_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0.ppa_u0.d5_0.o2._2_  (.I(\mult_add_u0.add0.ppa_u0.d5_0.o2._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.cg43 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.add0.ppa_u0.d5_1.a2._1_  (.A1(\mult_add_u0.add0.ppa_u0.cg[2] ),
    .A2(\mult_add_u0.add0.ppa_u0.cp43 ),
    .Z(\mult_add_u0.add0.ppa_u0.d5_1.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0.ppa_u0.d5_1.a2._2_  (.I(\mult_add_u0.add0.ppa_u0.d5_1.a2._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.d5_1.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.add0.ppa_u0.d5_1.o2._1_  (.A1(\mult_add_u0.add0.ppa_u0.cg43 ),
    .A2(\mult_add_u0.add0.ppa_u0.d5_1.a2.out ),
    .Z(\mult_add_u0.add0.ppa_u0.d5_1.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0.ppa_u0.d5_1.o2._2_  (.I(\mult_add_u0.add0.ppa_u0.d5_1.o2._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.cg[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.add0.ppa_u0.d6_0.a1._1_  (.A1(\mult_add_u0.add0.ppa_u0.cp43 ),
    .A2(\mult_add_u0.add0.ppa_u0.d6_0.a1.in0 ),
    .Z(\mult_add_u0.add0.ppa_u0.d6_0.a1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0.ppa_u0.d6_0.a1._2_  (.I(\mult_add_u0.add0.ppa_u0.d6_0.a1._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.cp54 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.add0.ppa_u0.d6_0.a2._1_  (.A1(\mult_add_u0.add0.ppa_u0.cg43 ),
    .A2(\mult_add_u0.add0.ppa_u0.d6_0.a1.in0 ),
    .Z(\mult_add_u0.add0.ppa_u0.d6_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0.ppa_u0.d6_0.a2._2_  (.I(\mult_add_u0.add0.ppa_u0.d6_0.a2._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.d6_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.add0.ppa_u0.d6_0.o2._1_  (.A1(\mult_add_u0.add0.ppa_u0.d6_0.g1 ),
    .A2(\mult_add_u0.add0.ppa_u0.d6_0.a2.out ),
    .Z(\mult_add_u0.add0.ppa_u0.d6_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0.ppa_u0.d6_0.o2._2_  (.I(\mult_add_u0.add0.ppa_u0.d6_0.o2._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.cg54 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.add0.ppa_u0.d6_1.a2._1_  (.A1(\mult_add_u0.add0.ppa_u0.cg[2] ),
    .A2(\mult_add_u0.add0.ppa_u0.cp54 ),
    .Z(\mult_add_u0.add0.ppa_u0.d6_1.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0.ppa_u0.d6_1.a2._2_  (.I(\mult_add_u0.add0.ppa_u0.d6_1.a2._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.d6_1.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.add0.ppa_u0.d6_1.o2._1_  (.A1(\mult_add_u0.add0.ppa_u0.cg54 ),
    .A2(\mult_add_u0.add0.ppa_u0.d6_1.a2.out ),
    .Z(\mult_add_u0.add0.ppa_u0.d6_1.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0.ppa_u0.d6_1.o2._2_  (.I(\mult_add_u0.add0.ppa_u0.d6_1.o2._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.cg[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.add0.ppa_u0.p_0.a._1_  (.A1(\mult_add_u0.add0.b_in[0] ),
    .A2(\mult_add_u0.add0.a_in[0] ),
    .Z(\mult_add_u0.add0.ppa_u0.p_0.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0.ppa_u0.p_0.a._2_  (.I(\mult_add_u0.add0.ppa_u0.p_0.a._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.d1_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.add0.ppa_u0.p_0.o._1_  (.A1(\mult_add_u0.add0.b_in[0] ),
    .A2(\mult_add_u0.add0.a_in[0] ),
    .Z(\mult_add_u0.add0.ppa_u0.p_0.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0.ppa_u0.p_0.o._2_  (.I(\mult_add_u0.add0.ppa_u0.p_0.o._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.d1_0.a2.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.add0.ppa_u0.p_1.a._1_  (.A1(\mult_add_u0.add0.b_in[1] ),
    .A2(\mult_add_u0.add0.a_in[1] ),
    .Z(\mult_add_u0.add0.ppa_u0.p_1.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0.ppa_u0.p_1.a._2_  (.I(\mult_add_u0.add0.ppa_u0.p_1.a._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.d2_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.add0.ppa_u0.p_1.o._1_  (.A1(\mult_add_u0.add0.b_in[1] ),
    .A2(\mult_add_u0.add0.a_in[1] ),
    .Z(\mult_add_u0.add0.ppa_u0.p_1.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0.ppa_u0.p_1.o._2_  (.I(\mult_add_u0.add0.ppa_u0.p_1.o._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.d2_0.a2.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.add0.ppa_u0.p_2.a._1_  (.A1(\mult_add_u0.add0.b_in[2] ),
    .A2(\mult_add_u0.add0.a_in[2] ),
    .Z(\mult_add_u0.add0.ppa_u0.p_2.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0.ppa_u0.p_2.a._2_  (.I(\mult_add_u0.add0.ppa_u0.p_2.a._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.d3_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.add0.ppa_u0.p_2.o._1_  (.A1(\mult_add_u0.add0.b_in[2] ),
    .A2(\mult_add_u0.add0.a_in[2] ),
    .Z(\mult_add_u0.add0.ppa_u0.p_2.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0.ppa_u0.p_2.o._2_  (.I(\mult_add_u0.add0.ppa_u0.p_2.o._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.d3_0.a1.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.add0.ppa_u0.p_3.a._1_  (.A1(\mult_add_u0.add0.b_in[3] ),
    .A2(\mult_add_u0.add0.a_in[3] ),
    .Z(\mult_add_u0.add0.ppa_u0.p_3.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0.ppa_u0.p_3.a._2_  (.I(\mult_add_u0.add0.ppa_u0.p_3.a._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.d4_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.add0.ppa_u0.p_3.o._1_  (.A1(\mult_add_u0.add0.b_in[3] ),
    .A2(\mult_add_u0.add0.a_in[3] ),
    .Z(\mult_add_u0.add0.ppa_u0.p_3.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0.ppa_u0.p_3.o._2_  (.I(\mult_add_u0.add0.ppa_u0.p_3.o._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.d4_0.a2.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.add0.ppa_u0.p_4.a._1_  (.A1(\mult_add_u0.add0.b_in[4] ),
    .A2(\mult_add_u0.add0.a_in[4] ),
    .Z(\mult_add_u0.add0.ppa_u0.p_4.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0.ppa_u0.p_4.a._2_  (.I(\mult_add_u0.add0.ppa_u0.p_4.a._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.d5_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.add0.ppa_u0.p_4.o._1_  (.A1(\mult_add_u0.add0.b_in[4] ),
    .A2(\mult_add_u0.add0.a_in[4] ),
    .Z(\mult_add_u0.add0.ppa_u0.p_4.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0.ppa_u0.p_4.o._2_  (.I(\mult_add_u0.add0.ppa_u0.p_4.o._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.d5_0.a1.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.add0.ppa_u0.p_5.a._1_  (.A1(\mult_add_u0.add0.b_in[5] ),
    .A2(\mult_add_u0.add0.a_in[5] ),
    .Z(\mult_add_u0.add0.ppa_u0.p_5.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0.ppa_u0.p_5.a._2_  (.I(\mult_add_u0.add0.ppa_u0.p_5.a._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.d6_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.add0.ppa_u0.p_5.o._1_  (.A1(\mult_add_u0.add0.b_in[5] ),
    .A2(\mult_add_u0.add0.a_in[5] ),
    .Z(\mult_add_u0.add0.ppa_u0.p_5.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0.ppa_u0.p_5.o._2_  (.I(\mult_add_u0.add0.ppa_u0.p_5.o._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.d6_0.a1.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.add0.ppa_u0.s0.xor2_0._1_  (.A1(\mult_add_u0.add0.b_in[0] ),
    .A2(\mult_add_u0.add0.a_in[0] ),
    .Z(\mult_add_u0.add0.ppa_u0.s0.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0.ppa_u0.s0.xor2_0._2_  (.I(\mult_add_u0.add0.ppa_u0.s0.xor2_0._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.s0.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.add0.ppa_u0.s0.xor2_1._1_  (.A1(\mult_add_u0.add0.ppa_u0.s0.temp ),
    .A2(\mult_add_u0.add0.c_in ),
    .Z(\mult_add_u0.add0.ppa_u0.s0.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0.ppa_u0.s0.xor2_1._2_  (.I(\mult_add_u0.add0.ppa_u0.s0.xor2_1._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.S[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.add0.ppa_u0.s1.xor2_0._1_  (.A1(\mult_add_u0.add0.b_in[1] ),
    .A2(\mult_add_u0.add0.a_in[1] ),
    .Z(\mult_add_u0.add0.ppa_u0.s1.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0.ppa_u0.s1.xor2_0._2_  (.I(\mult_add_u0.add0.ppa_u0.s1.xor2_0._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.s1.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.add0.ppa_u0.s1.xor2_1._1_  (.A1(\mult_add_u0.add0.ppa_u0.s1.temp ),
    .A2(\mult_add_u0.add0.ppa_u0.cg[0] ),
    .Z(\mult_add_u0.add0.ppa_u0.s1.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0.ppa_u0.s1.xor2_1._2_  (.I(\mult_add_u0.add0.ppa_u0.s1.xor2_1._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.S[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.add0.ppa_u0.s2.xor2_0._1_  (.A1(\mult_add_u0.add0.b_in[2] ),
    .A2(\mult_add_u0.add0.a_in[2] ),
    .Z(\mult_add_u0.add0.ppa_u0.s2.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0.ppa_u0.s2.xor2_0._2_  (.I(\mult_add_u0.add0.ppa_u0.s2.xor2_0._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.s2.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.add0.ppa_u0.s2.xor2_1._1_  (.A1(\mult_add_u0.add0.ppa_u0.s2.temp ),
    .A2(\mult_add_u0.add0.ppa_u0.cg[1] ),
    .Z(\mult_add_u0.add0.ppa_u0.s2.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0.ppa_u0.s2.xor2_1._2_  (.I(\mult_add_u0.add0.ppa_u0.s2.xor2_1._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.S[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.add0.ppa_u0.s3.xor2_0._1_  (.A1(\mult_add_u0.add0.b_in[3] ),
    .A2(\mult_add_u0.add0.a_in[3] ),
    .Z(\mult_add_u0.add0.ppa_u0.s3.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0.ppa_u0.s3.xor2_0._2_  (.I(\mult_add_u0.add0.ppa_u0.s3.xor2_0._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.s3.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.add0.ppa_u0.s3.xor2_1._1_  (.A1(\mult_add_u0.add0.ppa_u0.s3.temp ),
    .A2(\mult_add_u0.add0.ppa_u0.cg[2] ),
    .Z(\mult_add_u0.add0.ppa_u0.s3.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0.ppa_u0.s3.xor2_1._2_  (.I(\mult_add_u0.add0.ppa_u0.s3.xor2_1._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.S[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.add0.ppa_u0.s4.xor2_0._1_  (.A1(\mult_add_u0.add0.b_in[4] ),
    .A2(\mult_add_u0.add0.a_in[4] ),
    .Z(\mult_add_u0.add0.ppa_u0.s4.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0.ppa_u0.s4.xor2_0._2_  (.I(\mult_add_u0.add0.ppa_u0.s4.xor2_0._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.s4.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.add0.ppa_u0.s4.xor2_1._1_  (.A1(\mult_add_u0.add0.ppa_u0.s4.temp ),
    .A2(\mult_add_u0.add0.ppa_u0.cg[3] ),
    .Z(\mult_add_u0.add0.ppa_u0.s4.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0.ppa_u0.s4.xor2_1._2_  (.I(\mult_add_u0.add0.ppa_u0.s4.xor2_1._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.S[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.add0.ppa_u0.s5.xor2_0._1_  (.A1(\mult_add_u0.add0.b_in[5] ),
    .A2(\mult_add_u0.add0.a_in[5] ),
    .Z(\mult_add_u0.add0.ppa_u0.s5.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0.ppa_u0.s5.xor2_0._2_  (.I(\mult_add_u0.add0.ppa_u0.s5.xor2_0._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.s5.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.add0.ppa_u0.s5.xor2_1._1_  (.A1(\mult_add_u0.add0.ppa_u0.s5.temp ),
    .A2(\mult_add_u0.add0.ppa_u0.cg[4] ),
    .Z(\mult_add_u0.add0.ppa_u0.s5.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0.ppa_u0.s5.xor2_1._2_  (.I(\mult_add_u0.add0.ppa_u0.s5.xor2_1._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.S[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.add0.ppa_u0.s6.xor2_0._1_  (.A1(\mult_add_u0.add0.b_in[6] ),
    .A2(\mult_add_u0.add0.a_in[6] ),
    .Z(\mult_add_u0.add0.ppa_u0.s6.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0.ppa_u0.s6.xor2_0._2_  (.I(\mult_add_u0.add0.ppa_u0.s6.xor2_0._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.s6.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.add0.ppa_u0.s6.xor2_1._1_  (.A1(\mult_add_u0.add0.ppa_u0.s6.temp ),
    .A2(\mult_add_u0.add0.ppa_u0.cg[5] ),
    .Z(\mult_add_u0.add0.ppa_u0.s6.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.add0.ppa_u0.s6.xor2_1._2_  (.I(\mult_add_u0.add0.ppa_u0.s6.xor2_1._0_ ),
    .Z(\mult_add_u0.add0.ppa_u0.S[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \mult_add_u0.mult0._025_  (.I(\mult_add_u0.mult0.product[3] ),
    .ZN(\mult_add_u0.mult0._008_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \mult_add_u0.mult0._026_  (.I(net62),
    .Z(\mult_add_u0.mult0._009_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \mult_add_u0.mult0._027_  (.A1(\mult_add_u0.mult0._008_ ),
    .A2(\mult_add_u0.mult0._009_ ),
    .ZN(\mult_add_u0.mult0._000_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \mult_add_u0.mult0._028_  (.I(\mult_add_u0.mult0.product[4] ),
    .ZN(\mult_add_u0.mult0._010_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \mult_add_u0.mult0._029_  (.A1(\mult_add_u0.mult0._009_ ),
    .A2(\mult_add_u0.mult0._010_ ),
    .ZN(\mult_add_u0.mult0._001_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \mult_add_u0.mult0._030_  (.I(\mult_add_u0.mult0.product[5] ),
    .ZN(\mult_add_u0.mult0._011_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \mult_add_u0.mult0._031_  (.A1(\mult_add_u0.mult0._009_ ),
    .A2(\mult_add_u0.mult0._011_ ),
    .ZN(\mult_add_u0.mult0._002_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \mult_add_u0.mult0._032_  (.I(\mult_add_u0.mult0.product[6] ),
    .ZN(\mult_add_u0.mult0._012_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \mult_add_u0.mult0._033_  (.A1(\mult_add_u0.mult0._009_ ),
    .A2(\mult_add_u0.mult0._012_ ),
    .ZN(\mult_add_u0.mult0._003_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \mult_add_u0.mult0._034_  (.I(\mult_add_u0.mult0.step7.next_acc[0] ),
    .ZN(\mult_add_u0.mult0._013_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \mult_add_u0.mult0._035_  (.A1(\mult_add_u0.mult0._009_ ),
    .A2(\mult_add_u0.mult0._013_ ),
    .ZN(\mult_add_u0.mult0._004_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \mult_add_u0.mult0._036_  (.I(\mult_add_u0.mult0.step7.next_acc[1] ),
    .ZN(\mult_add_u0.mult0._014_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \mult_add_u0.mult0._037_  (.A1(\mult_add_u0.mult0._009_ ),
    .A2(\mult_add_u0.mult0._014_ ),
    .ZN(\mult_add_u0.mult0._005_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \mult_add_u0.mult0._038_  (.I(\mult_add_u0.mult0.step7.next_acc[2] ),
    .ZN(\mult_add_u0.mult0._015_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \mult_add_u0.mult0._039_  (.A1(\mult_add_u0.mult0._009_ ),
    .A2(\mult_add_u0.mult0._015_ ),
    .ZN(\mult_add_u0.mult0._006_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \mult_add_u0.mult0._040_  (.I(\mult_add_u0.mult0.mul_sign_s6 ),
    .ZN(\mult_add_u0.mult0._016_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \mult_add_u0.mult0._041_  (.A1(\mult_add_u0.mult0._009_ ),
    .A2(\mult_add_u0.mult0._016_ ),
    .ZN(\mult_add_u0.mult0._007_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._042_  (.D(\mult_add_u0.mult0._000_ ),
    .CLK(clknet_leaf_54_clk),
    .Q(\mult_add_u0.add0.a[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._043_  (.D(\mult_add_u0.mult0._001_ ),
    .CLK(clknet_leaf_51_clk),
    .Q(\mult_add_u0.add0.a[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._044_  (.D(\mult_add_u0.mult0._002_ ),
    .CLK(clknet_leaf_51_clk),
    .Q(\mult_add_u0.add0.a[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._045_  (.D(\mult_add_u0.mult0._003_ ),
    .CLK(clknet_leaf_51_clk),
    .Q(\mult_add_u0.add0.a[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._046_  (.D(\mult_add_u0.mult0._004_ ),
    .CLK(clknet_leaf_51_clk),
    .Q(\mult_add_u0.add0.a[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._047_  (.D(\mult_add_u0.mult0._005_ ),
    .CLK(clknet_leaf_50_clk),
    .Q(\mult_add_u0.add0.a[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._048_  (.D(\mult_add_u0.mult0._006_ ),
    .CLK(clknet_leaf_50_clk),
    .Q(\mult_add_u0.add0.a[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._049_  (.D(\mult_add_u0.mult0._007_ ),
    .CLK(clknet_leaf_53_clk),
    .Q(\mult_add_u0.add0.a[7] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._050_  (.D(\mult_add_u0.mult0.acc[1][0] ),
    .CLK(clknet_leaf_81_clk),
    .Q(\mult_add_u0.mult0.acc_s1[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._051_  (.D(\mult_add_u0.mult0.acc[1][1] ),
    .CLK(clknet_leaf_73_clk),
    .Q(\mult_add_u0.mult0.acc_s1[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._052_  (.D(\mult_add_u0.mult0.acc[1][2] ),
    .CLK(clknet_leaf_73_clk),
    .Q(\mult_add_u0.mult0.acc_s1[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._053_  (.D(\mult_add_u0.mult0.acc[1][3] ),
    .CLK(clknet_3_4__leaf_clk),
    .Q(\mult_add_u0.mult0.acc_s1[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._054_  (.D(\mult_add_u0.mult0.acc[1][4] ),
    .CLK(clknet_leaf_69_clk),
    .Q(\mult_add_u0.mult0.acc_s1[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._055_  (.D(\mult_add_u0.mult0.acc[1][5] ),
    .CLK(clknet_leaf_67_clk),
    .Q(\mult_add_u0.mult0.acc_s1[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._056_  (.D(\mult_add_u0.mult0.acc[1][6] ),
    .CLK(clknet_leaf_67_clk),
    .Q(\mult_add_u0.mult0.acc_s1[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 \mult_add_u0.mult0._057_  (.D(\mult_add_u0.mult0.Q[0][0] ),
    .CLK(clknet_leaf_71_clk),
    .Q(\mult_add_u0.mult0.Q_s1[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._058_  (.D(\mult_add_u0.mult0.Q[0][1] ),
    .CLK(clknet_leaf_69_clk),
    .Q(\mult_add_u0.mult0.Q_s1[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._059_  (.D(\mult_add_u0.mult0.Q[0][2] ),
    .CLK(clknet_leaf_69_clk),
    .Q(\mult_add_u0.mult0.Q_s1[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._060_  (.D(\mult_add_u0.mult0.Q[0][3] ),
    .CLK(clknet_leaf_65_clk),
    .Q(\mult_add_u0.mult0.Q_s1[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._061_  (.D(\mult_add_u0.mult0.Q[0][4] ),
    .CLK(clknet_leaf_65_clk),
    .Q(\mult_add_u0.mult0.Q_s1[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._062_  (.D(\mult_add_u0.mult0.Q[0][5] ),
    .CLK(clknet_leaf_64_clk),
    .Q(\mult_add_u0.mult0.Q_s1[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._064_  (.D(\mult_add_u0.mult0.acc[2][0] ),
    .CLK(clknet_leaf_76_clk),
    .Q(\mult_add_u0.mult0.acc_s2[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._065_  (.D(\mult_add_u0.mult0.acc[2][1] ),
    .CLK(clknet_leaf_75_clk),
    .Q(\mult_add_u0.mult0.acc_s2[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._066_  (.D(\mult_add_u0.mult0.acc[2][2] ),
    .CLK(clknet_leaf_75_clk),
    .Q(\mult_add_u0.mult0.acc_s2[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._067_  (.D(\mult_add_u0.mult0.acc[2][3] ),
    .CLK(clknet_leaf_61_clk),
    .Q(\mult_add_u0.mult0.acc_s2[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._068_  (.D(\mult_add_u0.mult0.acc[2][4] ),
    .CLK(clknet_leaf_61_clk),
    .Q(\mult_add_u0.mult0.acc_s2[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._069_  (.D(\mult_add_u0.mult0.acc[2][5] ),
    .CLK(clknet_leaf_62_clk),
    .Q(\mult_add_u0.mult0.acc_s2[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._070_  (.D(\mult_add_u0.mult0.acc[2][6] ),
    .CLK(clknet_leaf_62_clk),
    .Q(\mult_add_u0.mult0.acc_s2[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 \mult_add_u0.mult0._071_  (.D(\mult_add_u0.mult0.Q[1][0] ),
    .CLK(clknet_leaf_69_clk),
    .Q(\mult_add_u0.mult0.Q_s2[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._072_  (.D(\mult_add_u0.mult0.Q[1][1] ),
    .CLK(clknet_leaf_69_clk),
    .Q(\mult_add_u0.mult0.Q_s2[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._073_  (.D(\mult_add_u0.mult0.Q[1][2] ),
    .CLK(clknet_leaf_63_clk),
    .Q(\mult_add_u0.mult0.Q_s2[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._074_  (.D(\mult_add_u0.mult0.Q[1][3] ),
    .CLK(clknet_leaf_65_clk),
    .Q(\mult_add_u0.mult0.Q_s2[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._075_  (.D(\mult_add_u0.mult0.Q[1][4] ),
    .CLK(clknet_leaf_63_clk),
    .Q(\mult_add_u0.mult0.Q_s2[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._078_  (.D(\mult_add_u0.mult0.acc[3][0] ),
    .CLK(clknet_leaf_55_clk),
    .Q(\mult_add_u0.mult0.acc_s3[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._079_  (.D(\mult_add_u0.mult0.acc[3][1] ),
    .CLK(clknet_leaf_56_clk),
    .Q(\mult_add_u0.mult0.acc_s3[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._080_  (.D(\mult_add_u0.mult0.acc[3][2] ),
    .CLK(clknet_leaf_56_clk),
    .Q(\mult_add_u0.mult0.acc_s3[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._081_  (.D(\mult_add_u0.mult0.acc[3][3] ),
    .CLK(clknet_leaf_60_clk),
    .Q(\mult_add_u0.mult0.acc_s3[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._082_  (.D(\mult_add_u0.mult0.acc[3][4] ),
    .CLK(clknet_leaf_59_clk),
    .Q(\mult_add_u0.mult0.acc_s3[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._083_  (.D(\mult_add_u0.mult0.acc[3][5] ),
    .CLK(clknet_leaf_59_clk),
    .Q(\mult_add_u0.mult0.acc_s3[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._084_  (.D(\mult_add_u0.mult0.acc[3][6] ),
    .CLK(clknet_leaf_59_clk),
    .Q(\mult_add_u0.mult0.acc_s3[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 \mult_add_u0.mult0._085_  (.D(\mult_add_u0.mult0.Q[2][0] ),
    .CLK(clknet_leaf_66_clk),
    .Q(\mult_add_u0.mult0.Q_s3[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._086_  (.D(\mult_add_u0.mult0.Q[2][1] ),
    .CLK(clknet_leaf_62_clk),
    .Q(\mult_add_u0.mult0.Q_s3[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._087_  (.D(\mult_add_u0.mult0.Q[2][2] ),
    .CLK(clknet_leaf_63_clk),
    .Q(\mult_add_u0.mult0.Q_s3[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._088_  (.D(\mult_add_u0.mult0.Q[2][3] ),
    .CLK(clknet_leaf_63_clk),
    .Q(\mult_add_u0.mult0.Q_s3[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._092_  (.D(\mult_add_u0.mult0.acc[4][0] ),
    .CLK(clknet_leaf_54_clk),
    .Q(\mult_add_u0.mult0.acc_s4[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._093_  (.D(\mult_add_u0.mult0.acc[4][1] ),
    .CLK(clknet_leaf_57_clk),
    .Q(\mult_add_u0.mult0.acc_s4[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._094_  (.D(\mult_add_u0.mult0.acc[4][2] ),
    .CLK(clknet_leaf_57_clk),
    .Q(\mult_add_u0.mult0.acc_s4[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._095_  (.D(\mult_add_u0.mult0.acc[4][3] ),
    .CLK(clknet_leaf_57_clk),
    .Q(\mult_add_u0.mult0.acc_s4[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._096_  (.D(\mult_add_u0.mult0.acc[4][4] ),
    .CLK(clknet_leaf_57_clk),
    .Q(\mult_add_u0.mult0.acc_s4[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._097_  (.D(\mult_add_u0.mult0.acc[4][5] ),
    .CLK(clknet_leaf_57_clk),
    .Q(\mult_add_u0.mult0.acc_s4[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 \mult_add_u0.mult0._099_  (.D(\mult_add_u0.mult0.Q[3][0] ),
    .CLK(clknet_leaf_62_clk),
    .Q(\mult_add_u0.mult0.Q_s4[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._100_  (.D(\mult_add_u0.mult0.Q[3][1] ),
    .CLK(clknet_leaf_46_clk),
    .Q(\mult_add_u0.mult0.Q_s4[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._101_  (.D(\mult_add_u0.mult0.Q[3][2] ),
    .CLK(clknet_leaf_63_clk),
    .Q(\mult_add_u0.mult0.Q_s4[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._105_  (.D(\mult_add_u0.mult0.Q[3][6] ),
    .CLK(clknet_leaf_54_clk),
    .Q(\mult_add_u0.mult0.Q_s4[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._106_  (.D(\mult_add_u0.mult0.acc[5][0] ),
    .CLK(clknet_leaf_48_clk),
    .Q(\mult_add_u0.mult0.acc_s5[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._107_  (.D(\mult_add_u0.mult0.acc[5][1] ),
    .CLK(clknet_leaf_49_clk),
    .Q(\mult_add_u0.mult0.acc_s5[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._108_  (.D(\mult_add_u0.mult0.acc[5][2] ),
    .CLK(clknet_3_7__leaf_clk),
    .Q(\mult_add_u0.mult0.acc_s5[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._109_  (.D(\mult_add_u0.mult0.acc[5][3] ),
    .CLK(clknet_leaf_45_clk),
    .Q(\mult_add_u0.mult0.acc_s5[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._110_  (.D(\mult_add_u0.mult0.acc[5][4] ),
    .CLK(clknet_leaf_45_clk),
    .Q(\mult_add_u0.mult0.acc_s5[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 \mult_add_u0.mult0._113_  (.D(\mult_add_u0.mult0.Q[4][0] ),
    .CLK(clknet_leaf_46_clk),
    .Q(\mult_add_u0.mult0.Q_s5[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._114_  (.D(\mult_add_u0.mult0.Q[4][1] ),
    .CLK(clknet_leaf_58_clk),
    .Q(\mult_add_u0.mult0.Q_s5[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._118_  (.D(\mult_add_u0.mult0.Q[4][5] ),
    .CLK(clknet_leaf_53_clk),
    .Q(\mult_add_u0.mult0.Q_s5[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._119_  (.D(\mult_add_u0.mult0.Q[4][6] ),
    .CLK(clknet_leaf_48_clk),
    .Q(\mult_add_u0.mult0.Q_s5[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._120_  (.D(\mult_add_u0.mult0.acc[6][0] ),
    .CLK(clknet_leaf_50_clk),
    .Q(\mult_add_u0.mult0.acc_s6[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._121_  (.D(\mult_add_u0.mult0.acc[6][1] ),
    .CLK(clknet_leaf_44_clk),
    .Q(\mult_add_u0.mult0.acc_s6[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._122_  (.D(\mult_add_u0.mult0.acc[6][2] ),
    .CLK(clknet_3_7__leaf_clk),
    .Q(\mult_add_u0.mult0.acc_s6[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._123_  (.D(\mult_add_u0.mult0.acc[6][3] ),
    .CLK(clknet_leaf_44_clk),
    .Q(\mult_add_u0.mult0.acc_s6[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 \mult_add_u0.mult0._127_  (.D(\mult_add_u0.mult0.Q[5][0] ),
    .CLK(clknet_leaf_45_clk),
    .Q(\mult_add_u0.mult0.Q_s6[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._131_  (.D(\mult_add_u0.mult0.Q[5][4] ),
    .CLK(clknet_leaf_53_clk),
    .Q(\mult_add_u0.mult0.Q_s6[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._132_  (.D(\mult_add_u0.mult0.Q[5][5] ),
    .CLK(clknet_leaf_51_clk),
    .Q(\mult_add_u0.mult0.Q_s6[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._133_  (.D(\mult_add_u0.mult0.Q[5][6] ),
    .CLK(clknet_leaf_48_clk),
    .Q(\mult_add_u0.mult0.Q_s6[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._134_  (.D(\mult_add_u0.mult0.q0[1] ),
    .CLK(clknet_leaf_73_clk),
    .Q(\mult_add_u0.mult0.q0_s1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._135_  (.D(\mult_add_u0.mult0.q0[2] ),
    .CLK(clknet_leaf_60_clk),
    .Q(\mult_add_u0.mult0.q0_s2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._136_  (.D(\mult_add_u0.mult0.q0[3] ),
    .CLK(clknet_leaf_59_clk),
    .Q(\mult_add_u0.mult0.q0_s3 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._137_  (.D(\mult_add_u0.mult0.q0[4] ),
    .CLK(clknet_leaf_57_clk),
    .Q(\mult_add_u0.mult0.q0_s4 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._138_  (.D(\mult_add_u0.mult0.q0[5] ),
    .CLK(clknet_leaf_46_clk),
    .Q(\mult_add_u0.mult0.q0_s5 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._139_  (.D(\mult_add_u0.mult0.q0[6] ),
    .CLK(clknet_leaf_44_clk),
    .Q(\mult_add_u0.mult0.q0_s6 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._140_  (.D(\mult_add_u0.mult0.multiplicand[0] ),
    .CLK(clknet_leaf_81_clk),
    .Q(\mult_add_u0.mult0.multiplicand_s1[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._141_  (.D(\mult_add_u0.mult0.multiplicand[1] ),
    .CLK(clknet_leaf_77_clk),
    .Q(\mult_add_u0.mult0.multiplicand_s1[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._142_  (.D(\mult_add_u0.mult0.multiplicand[2] ),
    .CLK(clknet_leaf_81_clk),
    .Q(\mult_add_u0.mult0.multiplicand_s1[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._143_  (.D(\mult_add_u0.mult0.multiplicand[3] ),
    .CLK(clknet_leaf_73_clk),
    .Q(\mult_add_u0.mult0.multiplicand_s1[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._144_  (.D(\mult_add_u0.mult0.multiplicand[4] ),
    .CLK(clknet_leaf_69_clk),
    .Q(\mult_add_u0.mult0.multiplicand_s1[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._145_  (.D(\mult_add_u0.mult0.multiplicand[5] ),
    .CLK(clknet_leaf_66_clk),
    .Q(\mult_add_u0.mult0.multiplicand_s1[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._146_  (.D(\mult_add_u0.mult0.multiplicand[6] ),
    .CLK(clknet_leaf_66_clk),
    .Q(\mult_add_u0.mult0.multiplicand_s1[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._147_  (.D(\mult_add_u0.mult0.multiplicand_s1[0] ),
    .CLK(clknet_leaf_76_clk),
    .Q(\mult_add_u0.mult0.multiplicand_s2[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._148_  (.D(\mult_add_u0.mult0.multiplicand_s1[1] ),
    .CLK(clknet_leaf_76_clk),
    .Q(\mult_add_u0.mult0.multiplicand_s2[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._149_  (.D(\mult_add_u0.mult0.multiplicand_s1[2] ),
    .CLK(clknet_leaf_76_clk),
    .Q(\mult_add_u0.mult0.multiplicand_s2[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._150_  (.D(\mult_add_u0.mult0.multiplicand_s1[3] ),
    .CLK(clknet_leaf_68_clk),
    .Q(\mult_add_u0.mult0.multiplicand_s2[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._151_  (.D(\mult_add_u0.mult0.multiplicand_s1[4] ),
    .CLK(clknet_leaf_68_clk),
    .Q(\mult_add_u0.mult0.multiplicand_s2[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._152_  (.D(\mult_add_u0.mult0.multiplicand_s1[5] ),
    .CLK(clknet_leaf_65_clk),
    .Q(\mult_add_u0.mult0.multiplicand_s2[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._153_  (.D(\mult_add_u0.mult0.multiplicand_s1[6] ),
    .CLK(clknet_leaf_65_clk),
    .Q(\mult_add_u0.mult0.multiplicand_s2[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._154_  (.D(\mult_add_u0.mult0.multiplicand_s2[0] ),
    .CLK(clknet_leaf_55_clk),
    .Q(\mult_add_u0.mult0.multiplicand_s3[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._155_  (.D(\mult_add_u0.mult0.multiplicand_s2[1] ),
    .CLK(clknet_leaf_55_clk),
    .Q(\mult_add_u0.mult0.multiplicand_s3[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._156_  (.D(\mult_add_u0.mult0.multiplicand_s2[2] ),
    .CLK(clknet_leaf_55_clk),
    .Q(\mult_add_u0.mult0.multiplicand_s3[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._157_  (.D(\mult_add_u0.mult0.multiplicand_s2[3] ),
    .CLK(clknet_leaf_56_clk),
    .Q(\mult_add_u0.mult0.multiplicand_s3[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._158_  (.D(\mult_add_u0.mult0.multiplicand_s2[4] ),
    .CLK(clknet_leaf_60_clk),
    .Q(\mult_add_u0.mult0.multiplicand_s3[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._159_  (.D(\mult_add_u0.mult0.multiplicand_s2[5] ),
    .CLK(clknet_leaf_59_clk),
    .Q(\mult_add_u0.mult0.multiplicand_s3[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._160_  (.D(\mult_add_u0.mult0.multiplicand_s2[6] ),
    .CLK(clknet_leaf_62_clk),
    .Q(\mult_add_u0.mult0.multiplicand_s3[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._161_  (.D(\mult_add_u0.mult0.multiplicand_s3[0] ),
    .CLK(clknet_leaf_54_clk),
    .Q(\mult_add_u0.mult0.multiplicand_s4[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._162_  (.D(\mult_add_u0.mult0.multiplicand_s3[1] ),
    .CLK(clknet_leaf_51_clk),
    .Q(\mult_add_u0.mult0.multiplicand_s4[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._163_  (.D(\mult_add_u0.mult0.multiplicand_s3[2] ),
    .CLK(clknet_leaf_48_clk),
    .Q(\mult_add_u0.mult0.multiplicand_s4[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._164_  (.D(\mult_add_u0.mult0.multiplicand_s3[3] ),
    .CLK(clknet_leaf_57_clk),
    .Q(\mult_add_u0.mult0.multiplicand_s4[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._165_  (.D(\mult_add_u0.mult0.multiplicand_s3[4] ),
    .CLK(clknet_leaf_57_clk),
    .Q(\mult_add_u0.mult0.multiplicand_s4[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._166_  (.D(\mult_add_u0.mult0.multiplicand_s3[5] ),
    .CLK(clknet_leaf_58_clk),
    .Q(\mult_add_u0.mult0.multiplicand_s4[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._168_  (.D(\mult_add_u0.mult0.multiplicand_s4[0] ),
    .CLK(clknet_leaf_50_clk),
    .Q(\mult_add_u0.mult0.multiplicand_s5[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._169_  (.D(\mult_add_u0.mult0.multiplicand_s4[1] ),
    .CLK(clknet_leaf_48_clk),
    .Q(\mult_add_u0.mult0.multiplicand_s5[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._170_  (.D(\mult_add_u0.mult0.multiplicand_s4[2] ),
    .CLK(clknet_leaf_49_clk),
    .Q(\mult_add_u0.mult0.multiplicand_s5[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._171_  (.D(\mult_add_u0.mult0.multiplicand_s4[3] ),
    .CLK(clknet_leaf_46_clk),
    .Q(\mult_add_u0.mult0.multiplicand_s5[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._172_  (.D(\mult_add_u0.mult0.multiplicand_s4[4] ),
    .CLK(clknet_leaf_46_clk),
    .Q(\mult_add_u0.mult0.multiplicand_s5[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._175_  (.D(\mult_add_u0.mult0.multiplicand_s5[0] ),
    .CLK(clknet_leaf_50_clk),
    .Q(\mult_add_u0.mult0.multiplicand_s6[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._176_  (.D(\mult_add_u0.mult0.multiplicand_s5[1] ),
    .CLK(clknet_leaf_50_clk),
    .Q(\mult_add_u0.mult0.multiplicand_s6[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._177_  (.D(\mult_add_u0.mult0.multiplicand_s5[2] ),
    .CLK(clknet_leaf_44_clk),
    .Q(\mult_add_u0.mult0.multiplicand_s6[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._178_  (.D(\mult_add_u0.mult0.multiplicand_s5[3] ),
    .CLK(clknet_leaf_44_clk),
    .Q(\mult_add_u0.mult0.multiplicand_s6[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._182_  (.D(\add_u0.a[0] ),
    .CLK(clknet_leaf_96_clk),
    .Q(\mult_add_u0.mult0.multiplicand[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._183_  (.D(\add_u0.a[1] ),
    .CLK(clknet_leaf_0_clk),
    .Q(\mult_add_u0.mult0.multiplicand[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._184_  (.D(\add_u0.a[2] ),
    .CLK(clknet_leaf_9_clk),
    .Q(\mult_add_u0.mult0.multiplicand[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._185_  (.D(\add_u0.a[3] ),
    .CLK(clknet_leaf_91_clk),
    .Q(\mult_add_u0.mult0.multiplicand[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._186_  (.D(\add_u0.a[4] ),
    .CLK(clknet_leaf_88_clk),
    .Q(\mult_add_u0.mult0.multiplicand[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._187_  (.D(\add_u0.a[5] ),
    .CLK(clknet_leaf_87_clk),
    .Q(\mult_add_u0.mult0.multiplicand[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._188_  (.D(\add_u0.a[6] ),
    .CLK(clknet_leaf_89_clk),
    .Q(\mult_add_u0.mult0.multiplicand[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 \mult_add_u0.mult0._189_  (.D(\mult_add_u0.m[0] ),
    .CLK(clknet_leaf_71_clk),
    .Q(\mult_add_u0.mult0.multiplier[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._190_  (.D(\mult_add_u0.m[1] ),
    .CLK(clknet_leaf_71_clk),
    .Q(\mult_add_u0.mult0.multiplier[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._191_  (.D(\mult_add_u0.m[2] ),
    .CLK(clknet_leaf_71_clk),
    .Q(\mult_add_u0.mult0.multiplier[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._192_  (.D(\mult_add_u0.m[3] ),
    .CLK(clknet_leaf_70_clk),
    .Q(\mult_add_u0.mult0.multiplier[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._193_  (.D(net122),
    .CLK(clknet_leaf_65_clk),
    .Q(\mult_add_u0.mult0.multiplier[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._194_  (.D(net116),
    .CLK(clknet_leaf_66_clk),
    .Q(\mult_add_u0.mult0.multiplier[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._195_  (.D(net136),
    .CLK(clknet_leaf_64_clk),
    .Q(\mult_add_u0.mult0.multiplier[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._196_  (.D(\mult_add_u0.mult0.mul_sign ),
    .CLK(clknet_leaf_87_clk),
    .Q(\mult_add_u0.mult0.mul_sign_s1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._197_  (.D(\mult_add_u0.mult0.mul_sign_s1 ),
    .CLK(clknet_leaf_87_clk),
    .Q(\mult_add_u0.mult0.mul_sign_s2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._198_  (.D(\mult_add_u0.mult0.mul_sign_s2 ),
    .CLK(clknet_leaf_84_clk),
    .Q(\mult_add_u0.mult0.mul_sign_s3 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._199_  (.D(\mult_add_u0.mult0.mul_sign_s3 ),
    .CLK(clknet_leaf_80_clk),
    .Q(\mult_add_u0.mult0.mul_sign_s4 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._200_  (.D(net132),
    .CLK(clknet_leaf_77_clk),
    .Q(\mult_add_u0.mult0.mul_sign_s5 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_add_u0.mult0._201_  (.D(\mult_add_u0.mult0.mul_sign_s5 ),
    .CLK(clknet_leaf_77_clk),
    .Q(\mult_add_u0.mult0.mul_sign_s6 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step1._09_  (.A1(net88),
    .A2(\mult_add_u0.mult0.multiplier[0] ),
    .Z(\mult_add_u0.mult0.step1._00_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_add_u0.mult0.step1._09__88  (.ZN(net88),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 \mult_add_u0.mult0.step1._10_  (.I(\mult_add_u0.mult0.step1._00_ ),
    .Z(\mult_add_u0.mult0.step1._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.mult0.step1._11_  (.I0(net86),
    .I1(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.S[6] ),
    .S(\mult_add_u0.mult0.step1._01_ ),
    .Z(\mult_add_u0.mult0.step1._02_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_add_u0.mult0.step1._11__86  (.ZN(net86),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1._12_  (.I(\mult_add_u0.mult0.step1._02_ ),
    .Z(\mult_add_u0.mult0.acc[1][6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.mult0.step1._13_  (.I0(net66),
    .I1(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.S[1] ),
    .S(\mult_add_u0.mult0.step1._01_ ),
    .Z(\mult_add_u0.mult0.step1._03_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_add_u0.mult0.step1._13__66  (.ZN(net66),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1._14_  (.I(\mult_add_u0.mult0.step1._03_ ),
    .Z(\mult_add_u0.mult0.acc[1][0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.mult0.step1._15_  (.I0(net70),
    .I1(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.S[2] ),
    .S(\mult_add_u0.mult0.step1._01_ ),
    .Z(\mult_add_u0.mult0.step1._04_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_add_u0.mult0.step1._15__70  (.ZN(net70),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1._16_  (.I(\mult_add_u0.mult0.step1._04_ ),
    .Z(\mult_add_u0.mult0.acc[1][1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.mult0.step1._17_  (.I0(net74),
    .I1(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.S[3] ),
    .S(\mult_add_u0.mult0.step1._01_ ),
    .Z(\mult_add_u0.mult0.step1._05_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_add_u0.mult0.step1._17__74  (.ZN(net74),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1._18_  (.I(\mult_add_u0.mult0.step1._05_ ),
    .Z(\mult_add_u0.mult0.acc[1][2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.mult0.step1._19_  (.I0(net78),
    .I1(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.S[4] ),
    .S(\mult_add_u0.mult0.step1._01_ ),
    .Z(\mult_add_u0.mult0.step1._06_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_add_u0.mult0.step1._19__78  (.ZN(net78),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1._20_  (.I(\mult_add_u0.mult0.step1._06_ ),
    .Z(\mult_add_u0.mult0.acc[1][3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.mult0.step1._21_  (.I0(net82),
    .I1(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.S[5] ),
    .S(\mult_add_u0.mult0.step1._01_ ),
    .Z(\mult_add_u0.mult0.step1._07_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_add_u0.mult0.step1._21__82  (.ZN(net82),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1._22_  (.I(\mult_add_u0.mult0.step1._07_ ),
    .Z(\mult_add_u0.mult0.acc[1][4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1._25_  (.I(\mult_add_u0.mult0.multiplier[1] ),
    .Z(\mult_add_u0.mult0.Q[0][0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1._26_  (.I(\mult_add_u0.mult0.multiplier[2] ),
    .Z(\mult_add_u0.mult0.Q[0][1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1._27_  (.I(\mult_add_u0.mult0.multiplier[3] ),
    .Z(\mult_add_u0.mult0.Q[0][2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1._28_  (.I(\mult_add_u0.mult0.multiplier[4] ),
    .Z(\mult_add_u0.mult0.Q[0][3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1._29_  (.I(\mult_add_u0.mult0.multiplier[5] ),
    .Z(\mult_add_u0.mult0.Q[0][4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1._30_  (.I(\mult_add_u0.mult0.multiplier[6] ),
    .Z(\mult_add_u0.mult0.Q[0][5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1._31_  (.I(\mult_add_u0.mult0.acc[1][6] ),
    .Z(\mult_add_u0.mult0.acc[1][5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1._32_  (.I(\mult_add_u0.mult0.multiplier[0] ),
    .Z(\mult_add_u0.mult0.q0[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d1_0.a2._1_  (.A1(\mult_add_u0.mult0.multiplier[0] ),
    .A2(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d1_0.a2.in0 ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d1_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d1_0.a2._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d1_0.a2._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d1_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d1_0.o2._1_  (.A1(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d1_0.g1 ),
    .A2(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d1_0.a2.out ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d1_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d1_0.o2._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d1_0.o2._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.cg[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d2_0.a2._1_  (.A1(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.cg[0] ),
    .A2(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d2_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d2_0.a2._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d2_0.a2._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d2_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d2_0.o2._1_  (.A1(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d2_0.g1 ),
    .A2(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d2_0.a2.out ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d2_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d2_0.o2._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d2_0.o2._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.cg[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d3_0.a1._1_  (.A1(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ),
    .A2(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d3_0.a1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d3_0.a1._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d3_0.a1._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.cp21 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d3_0.a2._1_  (.A1(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d2_0.g1 ),
    .A2(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d3_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d3_0.a2._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d3_0.a2._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d3_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d3_0.o2._1_  (.A1(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d3_0.g1 ),
    .A2(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d3_0.a2.out ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d3_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d3_0.o2._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d3_0.o2._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.cg21 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d3_1.a2._1_  (.A1(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.cg[0] ),
    .A2(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.cp21 ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d3_1.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d3_1.a2._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d3_1.a2._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d3_1.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d3_1.o2._1_  (.A1(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.cg21 ),
    .A2(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d3_1.a2.out ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d3_1.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d3_1.o2._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d3_1.o2._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.cg[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d4_0.a2._1_  (.A1(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.cg[2] ),
    .A2(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d4_0.a2.in0 ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d4_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d4_0.a2._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d4_0.a2._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d4_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d4_0.o2._1_  (.A1(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d4_0.g1 ),
    .A2(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d4_0.a2.out ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d4_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d4_0.o2._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d4_0.o2._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.cg[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d5_0.a1._1_  (.A1(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d4_0.a2.in0 ),
    .A2(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d5_0.a1.in0 ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d5_0.a1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d5_0.a1._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d5_0.a1._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.cp43 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d5_0.a2._1_  (.A1(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d4_0.g1 ),
    .A2(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d5_0.a1.in0 ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d5_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d5_0.a2._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d5_0.a2._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d5_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d5_0.o2._1_  (.A1(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d5_0.g1 ),
    .A2(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d5_0.a2.out ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d5_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d5_0.o2._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d5_0.o2._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.cg43 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d5_1.a2._1_  (.A1(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.cg[2] ),
    .A2(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.cp43 ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d5_1.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d5_1.a2._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d5_1.a2._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d5_1.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d5_1.o2._1_  (.A1(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.cg43 ),
    .A2(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d5_1.a2.out ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d5_1.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d5_1.o2._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d5_1.o2._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.cg[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d6_0.a1._1_  (.A1(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.cp43 ),
    .A2(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d6_0.a1.in0 ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d6_0.a1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d6_0.a1._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d6_0.a1._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.cp54 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d6_0.a2._1_  (.A1(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.cg43 ),
    .A2(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d6_0.a1.in0 ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d6_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d6_0.a2._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d6_0.a2._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d6_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d6_0.o2._1_  (.A1(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d6_0.g1 ),
    .A2(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d6_0.a2.out ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d6_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d6_0.o2._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d6_0.o2._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.cg54 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d6_1.a2._1_  (.A1(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.cg[2] ),
    .A2(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.cp54 ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d6_1.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d6_1.a2._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d6_1.a2._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d6_1.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d6_1.o2._1_  (.A1(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.cg54 ),
    .A2(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d6_1.a2.out ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d6_1.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d6_1.o2._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d6_1.o2._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.cg[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_0.a._1_  (.A1(\mult_add_u0.mult0.step1.add_sub4_u0.int_ip[0] ),
    .A2(net64),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_0.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_0.a._1__64  (.ZN(net64),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_0.a._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_0.a._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d1_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_0.o._1_  (.A1(\mult_add_u0.mult0.step1.add_sub4_u0.int_ip[0] ),
    .A2(net65),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_0.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_0.o._1__65  (.ZN(net65),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_0.o._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_0.o._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d1_0.a2.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_1.a._1_  (.A1(\mult_add_u0.mult0.step1.add_sub4_u0.int_ip[1] ),
    .A2(net67),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_1.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_1.a._1__67  (.ZN(net67),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_1.a._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_1.a._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d2_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_1.o._1_  (.A1(\mult_add_u0.mult0.step1.add_sub4_u0.int_ip[1] ),
    .A2(net68),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_1.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_1.o._1__68  (.ZN(net68),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_1.o._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_1.o._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_2.a._1_  (.A1(\mult_add_u0.mult0.step1.add_sub4_u0.int_ip[2] ),
    .A2(net71),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_2.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_2.a._1__71  (.ZN(net71),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_2.a._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_2.a._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d3_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_2.o._1_  (.A1(\mult_add_u0.mult0.step1.add_sub4_u0.int_ip[2] ),
    .A2(net72),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_2.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_2.o._1__72  (.ZN(net72),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_2.o._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_2.o._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_3.a._1_  (.A1(\mult_add_u0.mult0.step1.add_sub4_u0.int_ip[3] ),
    .A2(net75),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_3.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_3.a._1__75  (.ZN(net75),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_3.a._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_3.a._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d4_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_3.o._1_  (.A1(\mult_add_u0.mult0.step1.add_sub4_u0.int_ip[3] ),
    .A2(net76),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_3.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_3.o._1__76  (.ZN(net76),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_3.o._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_3.o._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d4_0.a2.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_4.a._1_  (.A1(\mult_add_u0.mult0.step1.add_sub4_u0.int_ip[4] ),
    .A2(net79),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_4.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_4.a._1__79  (.ZN(net79),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_4.a._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_4.a._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d5_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_4.o._1_  (.A1(\mult_add_u0.mult0.step1.add_sub4_u0.int_ip[4] ),
    .A2(net80),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_4.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_4.o._1__80  (.ZN(net80),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_4.o._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_4.o._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d5_0.a1.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_5.a._1_  (.A1(\mult_add_u0.mult0.step1.add_sub4_u0.int_ip[5] ),
    .A2(net83),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_5.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_5.a._1__83  (.ZN(net83),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_5.a._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_5.a._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d6_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_5.o._1_  (.A1(\mult_add_u0.mult0.step1.add_sub4_u0.int_ip[5] ),
    .A2(net84),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_5.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_5.o._1__84  (.ZN(net84),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_5.o._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.p_5.o._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.d6_0.a1.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s1.xor2_0._1_  (.A1(\mult_add_u0.mult0.step1.add_sub4_u0.int_ip[1] ),
    .A2(net69),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s1.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s1.xor2_0._1__69  (.ZN(net69),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s1.xor2_0._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s1.xor2_0._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s1.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s1.xor2_1._1_  (.A1(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s1.temp ),
    .A2(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.cg[0] ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s1.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s1.xor2_1._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s1.xor2_1._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.S[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s2.xor2_0._1_  (.A1(\mult_add_u0.mult0.step1.add_sub4_u0.int_ip[2] ),
    .A2(net73),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s2.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s2.xor2_0._1__73  (.ZN(net73),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s2.xor2_0._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s2.xor2_0._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s2.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s2.xor2_1._1_  (.A1(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s2.temp ),
    .A2(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.cg[1] ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s2.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s2.xor2_1._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s2.xor2_1._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.S[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s3.xor2_0._1_  (.A1(\mult_add_u0.mult0.step1.add_sub4_u0.int_ip[3] ),
    .A2(net77),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s3.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s3.xor2_0._1__77  (.ZN(net77),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s3.xor2_0._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s3.xor2_0._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s3.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s3.xor2_1._1_  (.A1(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s3.temp ),
    .A2(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.cg[2] ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s3.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s3.xor2_1._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s3.xor2_1._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.S[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s4.xor2_0._1_  (.A1(\mult_add_u0.mult0.step1.add_sub4_u0.int_ip[4] ),
    .A2(net81),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s4.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s4.xor2_0._1__81  (.ZN(net81),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s4.xor2_0._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s4.xor2_0._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s4.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s4.xor2_1._1_  (.A1(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s4.temp ),
    .A2(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.cg[3] ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s4.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s4.xor2_1._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s4.xor2_1._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.S[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s5.xor2_0._1_  (.A1(\mult_add_u0.mult0.step1.add_sub4_u0.int_ip[5] ),
    .A2(net85),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s5.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s5.xor2_0._1__85  (.ZN(net85),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s5.xor2_0._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s5.xor2_0._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s5.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s5.xor2_1._1_  (.A1(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s5.temp ),
    .A2(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.cg[4] ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s5.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s5.xor2_1._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s5.xor2_1._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.S[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s6.xor2_0._1_  (.A1(\mult_add_u0.mult0.step1.add_sub4_u0.int_ip[6] ),
    .A2(net87),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s6.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s6.xor2_0._1__87  (.ZN(net87),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s6.xor2_0._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s6.xor2_0._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s6.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s6.xor2_1._1_  (.A1(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s6.temp ),
    .A2(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.cg[5] ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s6.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s6.xor2_1._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.s6.xor2_1._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.ppa8_u0.S[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step1.add_sub4_u0.x0._1_  (.A1(\mult_add_u0.mult0.multiplier[0] ),
    .A2(\mult_add_u0.mult0.multiplicand[0] ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.x0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1.add_sub4_u0.x0._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.x0._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.int_ip[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step1.add_sub4_u0.x1._1_  (.A1(\mult_add_u0.mult0.multiplier[0] ),
    .A2(\mult_add_u0.mult0.multiplicand[1] ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.x1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1.add_sub4_u0.x1._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.x1._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.int_ip[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step1.add_sub4_u0.x2._1_  (.A1(\mult_add_u0.mult0.multiplier[0] ),
    .A2(\mult_add_u0.mult0.multiplicand[2] ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.x2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1.add_sub4_u0.x2._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.x2._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.int_ip[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step1.add_sub4_u0.x3._1_  (.A1(\mult_add_u0.mult0.multiplier[0] ),
    .A2(\mult_add_u0.mult0.multiplicand[3] ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.x3._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1.add_sub4_u0.x3._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.x3._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.int_ip[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step1.add_sub4_u0.x4._1_  (.A1(\mult_add_u0.mult0.multiplier[0] ),
    .A2(\mult_add_u0.mult0.multiplicand[4] ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.x4._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1.add_sub4_u0.x4._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.x4._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.int_ip[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step1.add_sub4_u0.x5._1_  (.A1(\mult_add_u0.mult0.multiplier[0] ),
    .A2(\mult_add_u0.mult0.multiplicand[5] ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.x5._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1.add_sub4_u0.x5._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.x5._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.int_ip[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step1.add_sub4_u0.x6._1_  (.A1(\mult_add_u0.mult0.multiplier[0] ),
    .A2(\mult_add_u0.mult0.multiplicand[6] ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.x6._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step1.add_sub4_u0.x6._2_  (.I(\mult_add_u0.mult0.step1.add_sub4_u0.x6._0_ ),
    .Z(\mult_add_u0.mult0.step1.add_sub4_u0.int_ip[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step2._09_  (.A1(\mult_add_u0.mult0.q0_s1 ),
    .A2(\mult_add_u0.mult0.Q_s1[0] ),
    .Z(\mult_add_u0.mult0.step2._00_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 \mult_add_u0.mult0.step2._10_  (.I(\mult_add_u0.mult0.step2._00_ ),
    .Z(\mult_add_u0.mult0.step2._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.mult0.step2._11_  (.I0(\mult_add_u0.mult0.acc_s1[6] ),
    .I1(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.S[6] ),
    .S(\mult_add_u0.mult0.step2._01_ ),
    .Z(\mult_add_u0.mult0.step2._02_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2._12_  (.I(\mult_add_u0.mult0.step2._02_ ),
    .Z(\mult_add_u0.mult0.acc[2][6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.mult0.step2._13_  (.I0(\mult_add_u0.mult0.acc_s1[1] ),
    .I1(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.S[1] ),
    .S(\mult_add_u0.mult0.step2._01_ ),
    .Z(\mult_add_u0.mult0.step2._03_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2._14_  (.I(\mult_add_u0.mult0.step2._03_ ),
    .Z(\mult_add_u0.mult0.acc[2][0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.mult0.step2._15_  (.I0(\mult_add_u0.mult0.acc_s1[2] ),
    .I1(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.S[2] ),
    .S(\mult_add_u0.mult0.step2._01_ ),
    .Z(\mult_add_u0.mult0.step2._04_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2._16_  (.I(\mult_add_u0.mult0.step2._04_ ),
    .Z(\mult_add_u0.mult0.acc[2][1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.mult0.step2._17_  (.I0(\mult_add_u0.mult0.acc_s1[3] ),
    .I1(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.S[3] ),
    .S(\mult_add_u0.mult0.step2._01_ ),
    .Z(\mult_add_u0.mult0.step2._05_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2._18_  (.I(\mult_add_u0.mult0.step2._05_ ),
    .Z(\mult_add_u0.mult0.acc[2][2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.mult0.step2._19_  (.I0(\mult_add_u0.mult0.acc_s1[4] ),
    .I1(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.S[4] ),
    .S(\mult_add_u0.mult0.step2._01_ ),
    .Z(\mult_add_u0.mult0.step2._06_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2._20_  (.I(\mult_add_u0.mult0.step2._06_ ),
    .Z(\mult_add_u0.mult0.acc[2][3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.mult0.step2._21_  (.I0(\mult_add_u0.mult0.acc_s1[5] ),
    .I1(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.S[5] ),
    .S(\mult_add_u0.mult0.step2._01_ ),
    .Z(\mult_add_u0.mult0.step2._07_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2._22_  (.I(\mult_add_u0.mult0.step2._07_ ),
    .Z(\mult_add_u0.mult0.acc[2][4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2._25_  (.I(\mult_add_u0.mult0.Q_s1[1] ),
    .Z(\mult_add_u0.mult0.Q[1][0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2._26_  (.I(\mult_add_u0.mult0.Q_s1[2] ),
    .Z(\mult_add_u0.mult0.Q[1][1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2._27_  (.I(\mult_add_u0.mult0.Q_s1[3] ),
    .Z(\mult_add_u0.mult0.Q[1][2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2._28_  (.I(\mult_add_u0.mult0.Q_s1[4] ),
    .Z(\mult_add_u0.mult0.Q[1][3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2._29_  (.I(\mult_add_u0.mult0.Q_s1[5] ),
    .Z(\mult_add_u0.mult0.Q[1][4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2._31_  (.I(\mult_add_u0.mult0.acc[2][6] ),
    .Z(\mult_add_u0.mult0.acc[2][5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2._32_  (.I(\mult_add_u0.mult0.Q_s1[0] ),
    .Z(\mult_add_u0.mult0.q0[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d1_0.a2._1_  (.A1(\mult_add_u0.mult0.Q_s1[0] ),
    .A2(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d1_0.a2.in0 ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d1_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d1_0.a2._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d1_0.a2._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d1_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d1_0.o2._1_  (.A1(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d1_0.g1 ),
    .A2(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d1_0.a2.out ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d1_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d1_0.o2._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d1_0.o2._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.cg[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d2_0.a2._1_  (.A1(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.cg[0] ),
    .A2(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d2_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d2_0.a2._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d2_0.a2._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d2_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d2_0.o2._1_  (.A1(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d2_0.g1 ),
    .A2(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d2_0.a2.out ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d2_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d2_0.o2._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d2_0.o2._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.cg[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d3_0.a1._1_  (.A1(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ),
    .A2(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d3_0.a1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d3_0.a1._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d3_0.a1._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.cp21 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d3_0.a2._1_  (.A1(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d2_0.g1 ),
    .A2(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d3_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d3_0.a2._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d3_0.a2._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d3_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d3_0.o2._1_  (.A1(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d3_0.g1 ),
    .A2(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d3_0.a2.out ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d3_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d3_0.o2._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d3_0.o2._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.cg21 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d3_1.a2._1_  (.A1(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.cg[0] ),
    .A2(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.cp21 ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d3_1.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d3_1.a2._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d3_1.a2._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d3_1.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d3_1.o2._1_  (.A1(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.cg21 ),
    .A2(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d3_1.a2.out ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d3_1.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d3_1.o2._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d3_1.o2._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.cg[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d4_0.a2._1_  (.A1(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.cg[2] ),
    .A2(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d4_0.a2.in0 ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d4_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d4_0.a2._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d4_0.a2._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d4_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d4_0.o2._1_  (.A1(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d4_0.g1 ),
    .A2(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d4_0.a2.out ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d4_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d4_0.o2._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d4_0.o2._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.cg[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d5_0.a1._1_  (.A1(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d4_0.a2.in0 ),
    .A2(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d5_0.a1.in0 ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d5_0.a1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d5_0.a1._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d5_0.a1._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.cp43 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d5_0.a2._1_  (.A1(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d4_0.g1 ),
    .A2(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d5_0.a1.in0 ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d5_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d5_0.a2._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d5_0.a2._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d5_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d5_0.o2._1_  (.A1(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d5_0.g1 ),
    .A2(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d5_0.a2.out ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d5_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d5_0.o2._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d5_0.o2._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.cg43 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d5_1.a2._1_  (.A1(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.cg[2] ),
    .A2(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.cp43 ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d5_1.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d5_1.a2._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d5_1.a2._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d5_1.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d5_1.o2._1_  (.A1(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.cg43 ),
    .A2(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d5_1.a2.out ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d5_1.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d5_1.o2._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d5_1.o2._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.cg[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d6_0.a1._1_  (.A1(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.cp43 ),
    .A2(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d6_0.a1.in0 ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d6_0.a1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d6_0.a1._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d6_0.a1._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.cp54 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d6_0.a2._1_  (.A1(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.cg43 ),
    .A2(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d6_0.a1.in0 ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d6_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d6_0.a2._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d6_0.a2._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d6_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d6_0.o2._1_  (.A1(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d6_0.g1 ),
    .A2(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d6_0.a2.out ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d6_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d6_0.o2._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d6_0.o2._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.cg54 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d6_1.a2._1_  (.A1(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.cg[2] ),
    .A2(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.cp54 ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d6_1.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d6_1.a2._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d6_1.a2._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d6_1.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d6_1.o2._1_  (.A1(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.cg54 ),
    .A2(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d6_1.a2.out ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d6_1.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d6_1.o2._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d6_1.o2._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.cg[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_0.a._1_  (.A1(\mult_add_u0.mult0.step2.add_sub4_u0.int_ip[0] ),
    .A2(\mult_add_u0.mult0.acc_s1[0] ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_0.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_0.a._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_0.a._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d1_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_0.o._1_  (.A1(\mult_add_u0.mult0.step2.add_sub4_u0.int_ip[0] ),
    .A2(\mult_add_u0.mult0.acc_s1[0] ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_0.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_0.o._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_0.o._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d1_0.a2.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_1.a._1_  (.A1(\mult_add_u0.mult0.step2.add_sub4_u0.int_ip[1] ),
    .A2(\mult_add_u0.mult0.acc_s1[1] ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_1.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_1.a._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_1.a._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d2_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_1.o._1_  (.A1(\mult_add_u0.mult0.step2.add_sub4_u0.int_ip[1] ),
    .A2(\mult_add_u0.mult0.acc_s1[1] ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_1.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_1.o._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_1.o._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_2.a._1_  (.A1(\mult_add_u0.mult0.step2.add_sub4_u0.int_ip[2] ),
    .A2(\mult_add_u0.mult0.acc_s1[2] ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_2.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_2.a._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_2.a._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d3_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_2.o._1_  (.A1(\mult_add_u0.mult0.step2.add_sub4_u0.int_ip[2] ),
    .A2(\mult_add_u0.mult0.acc_s1[2] ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_2.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_2.o._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_2.o._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_3.a._1_  (.A1(\mult_add_u0.mult0.step2.add_sub4_u0.int_ip[3] ),
    .A2(\mult_add_u0.mult0.acc_s1[3] ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_3.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_3.a._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_3.a._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d4_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_3.o._1_  (.A1(\mult_add_u0.mult0.step2.add_sub4_u0.int_ip[3] ),
    .A2(\mult_add_u0.mult0.acc_s1[3] ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_3.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_3.o._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_3.o._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d4_0.a2.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_4.a._1_  (.A1(\mult_add_u0.mult0.step2.add_sub4_u0.int_ip[4] ),
    .A2(\mult_add_u0.mult0.acc_s1[4] ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_4.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_4.a._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_4.a._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d5_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_4.o._1_  (.A1(\mult_add_u0.mult0.step2.add_sub4_u0.int_ip[4] ),
    .A2(\mult_add_u0.mult0.acc_s1[4] ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_4.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_4.o._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_4.o._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d5_0.a1.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_5.a._1_  (.A1(\mult_add_u0.mult0.step2.add_sub4_u0.int_ip[5] ),
    .A2(\mult_add_u0.mult0.acc_s1[5] ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_5.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_5.a._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_5.a._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d6_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_5.o._1_  (.A1(\mult_add_u0.mult0.step2.add_sub4_u0.int_ip[5] ),
    .A2(\mult_add_u0.mult0.acc_s1[5] ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_5.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_5.o._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.p_5.o._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.d6_0.a1.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s1.xor2_0._1_  (.A1(\mult_add_u0.mult0.step2.add_sub4_u0.int_ip[1] ),
    .A2(\mult_add_u0.mult0.acc_s1[1] ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s1.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s1.xor2_0._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s1.xor2_0._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s1.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s1.xor2_1._1_  (.A1(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s1.temp ),
    .A2(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.cg[0] ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s1.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s1.xor2_1._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s1.xor2_1._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.S[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s2.xor2_0._1_  (.A1(\mult_add_u0.mult0.step2.add_sub4_u0.int_ip[2] ),
    .A2(\mult_add_u0.mult0.acc_s1[2] ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s2.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s2.xor2_0._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s2.xor2_0._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s2.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s2.xor2_1._1_  (.A1(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s2.temp ),
    .A2(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.cg[1] ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s2.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s2.xor2_1._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s2.xor2_1._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.S[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s3.xor2_0._1_  (.A1(\mult_add_u0.mult0.step2.add_sub4_u0.int_ip[3] ),
    .A2(\mult_add_u0.mult0.acc_s1[3] ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s3.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s3.xor2_0._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s3.xor2_0._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s3.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s3.xor2_1._1_  (.A1(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s3.temp ),
    .A2(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.cg[2] ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s3.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s3.xor2_1._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s3.xor2_1._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.S[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s4.xor2_0._1_  (.A1(\mult_add_u0.mult0.step2.add_sub4_u0.int_ip[4] ),
    .A2(\mult_add_u0.mult0.acc_s1[4] ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s4.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s4.xor2_0._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s4.xor2_0._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s4.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s4.xor2_1._1_  (.A1(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s4.temp ),
    .A2(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.cg[3] ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s4.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s4.xor2_1._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s4.xor2_1._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.S[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s5.xor2_0._1_  (.A1(\mult_add_u0.mult0.step2.add_sub4_u0.int_ip[5] ),
    .A2(\mult_add_u0.mult0.acc_s1[5] ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s5.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s5.xor2_0._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s5.xor2_0._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s5.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s5.xor2_1._1_  (.A1(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s5.temp ),
    .A2(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.cg[4] ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s5.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s5.xor2_1._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s5.xor2_1._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.S[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s6.xor2_0._1_  (.A1(\mult_add_u0.mult0.step2.add_sub4_u0.int_ip[6] ),
    .A2(\mult_add_u0.mult0.acc_s1[6] ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s6.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s6.xor2_0._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s6.xor2_0._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s6.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s6.xor2_1._1_  (.A1(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s6.temp ),
    .A2(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.cg[5] ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s6.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s6.xor2_1._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.s6.xor2_1._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.ppa8_u0.S[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step2.add_sub4_u0.x0._1_  (.A1(\mult_add_u0.mult0.Q_s1[0] ),
    .A2(\mult_add_u0.mult0.multiplicand_s1[0] ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.x0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.x0._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.x0._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.int_ip[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step2.add_sub4_u0.x1._1_  (.A1(\mult_add_u0.mult0.Q_s1[0] ),
    .A2(\mult_add_u0.mult0.multiplicand_s1[1] ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.x1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.x1._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.x1._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.int_ip[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step2.add_sub4_u0.x2._1_  (.A1(\mult_add_u0.mult0.Q_s1[0] ),
    .A2(\mult_add_u0.mult0.multiplicand_s1[2] ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.x2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.x2._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.x2._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.int_ip[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step2.add_sub4_u0.x3._1_  (.A1(\mult_add_u0.mult0.Q_s1[0] ),
    .A2(\mult_add_u0.mult0.multiplicand_s1[3] ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.x3._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.x3._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.x3._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.int_ip[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step2.add_sub4_u0.x4._1_  (.A1(\mult_add_u0.mult0.Q_s1[0] ),
    .A2(\mult_add_u0.mult0.multiplicand_s1[4] ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.x4._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.x4._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.x4._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.int_ip[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step2.add_sub4_u0.x5._1_  (.A1(\mult_add_u0.mult0.Q_s1[0] ),
    .A2(\mult_add_u0.mult0.multiplicand_s1[5] ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.x5._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.x5._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.x5._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.int_ip[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step2.add_sub4_u0.x6._1_  (.A1(\mult_add_u0.mult0.Q_s1[0] ),
    .A2(\mult_add_u0.mult0.multiplicand_s1[6] ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.x6._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step2.add_sub4_u0.x6._2_  (.I(\mult_add_u0.mult0.step2.add_sub4_u0.x6._0_ ),
    .Z(\mult_add_u0.mult0.step2.add_sub4_u0.int_ip[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step3._09_  (.A1(\mult_add_u0.mult0.q0_s2 ),
    .A2(\mult_add_u0.mult0.Q_s2[0] ),
    .Z(\mult_add_u0.mult0.step3._00_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 \mult_add_u0.mult0.step3._10_  (.I(\mult_add_u0.mult0.step3._00_ ),
    .Z(\mult_add_u0.mult0.step3._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.mult0.step3._11_  (.I0(\mult_add_u0.mult0.acc_s2[6] ),
    .I1(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.S[6] ),
    .S(\mult_add_u0.mult0.step3._01_ ),
    .Z(\mult_add_u0.mult0.step3._02_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3._12_  (.I(\mult_add_u0.mult0.step3._02_ ),
    .Z(\mult_add_u0.mult0.acc[3][6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.mult0.step3._13_  (.I0(\mult_add_u0.mult0.acc_s2[1] ),
    .I1(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.S[1] ),
    .S(\mult_add_u0.mult0.step3._01_ ),
    .Z(\mult_add_u0.mult0.step3._03_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3._14_  (.I(\mult_add_u0.mult0.step3._03_ ),
    .Z(\mult_add_u0.mult0.acc[3][0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.mult0.step3._15_  (.I0(\mult_add_u0.mult0.acc_s2[2] ),
    .I1(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.S[2] ),
    .S(\mult_add_u0.mult0.step3._01_ ),
    .Z(\mult_add_u0.mult0.step3._04_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3._16_  (.I(\mult_add_u0.mult0.step3._04_ ),
    .Z(\mult_add_u0.mult0.acc[3][1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.mult0.step3._17_  (.I0(\mult_add_u0.mult0.acc_s2[3] ),
    .I1(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.S[3] ),
    .S(\mult_add_u0.mult0.step3._01_ ),
    .Z(\mult_add_u0.mult0.step3._05_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3._18_  (.I(\mult_add_u0.mult0.step3._05_ ),
    .Z(\mult_add_u0.mult0.acc[3][2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.mult0.step3._19_  (.I0(\mult_add_u0.mult0.acc_s2[4] ),
    .I1(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.S[4] ),
    .S(\mult_add_u0.mult0.step3._01_ ),
    .Z(\mult_add_u0.mult0.step3._06_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3._20_  (.I(\mult_add_u0.mult0.step3._06_ ),
    .Z(\mult_add_u0.mult0.acc[3][3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.mult0.step3._21_  (.I0(\mult_add_u0.mult0.acc_s2[5] ),
    .I1(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.S[5] ),
    .S(\mult_add_u0.mult0.step3._01_ ),
    .Z(\mult_add_u0.mult0.step3._07_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3._22_  (.I(\mult_add_u0.mult0.step3._07_ ),
    .Z(\mult_add_u0.mult0.acc[3][4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3._25_  (.I(\mult_add_u0.mult0.Q_s2[1] ),
    .Z(\mult_add_u0.mult0.Q[2][0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3._26_  (.I(\mult_add_u0.mult0.Q_s2[2] ),
    .Z(\mult_add_u0.mult0.Q[2][1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3._27_  (.I(\mult_add_u0.mult0.Q_s2[3] ),
    .Z(\mult_add_u0.mult0.Q[2][2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3._28_  (.I(\mult_add_u0.mult0.Q_s2[4] ),
    .Z(\mult_add_u0.mult0.Q[2][3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3._31_  (.I(\mult_add_u0.mult0.acc[3][6] ),
    .Z(\mult_add_u0.mult0.acc[3][5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3._32_  (.I(\mult_add_u0.mult0.Q_s2[0] ),
    .Z(\mult_add_u0.mult0.q0[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d1_0.a2._1_  (.A1(\mult_add_u0.mult0.Q_s2[0] ),
    .A2(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d1_0.a2.in0 ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d1_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d1_0.a2._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d1_0.a2._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d1_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d1_0.o2._1_  (.A1(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d1_0.g1 ),
    .A2(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d1_0.a2.out ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d1_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d1_0.o2._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d1_0.o2._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.cg[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d2_0.a2._1_  (.A1(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.cg[0] ),
    .A2(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d2_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d2_0.a2._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d2_0.a2._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d2_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d2_0.o2._1_  (.A1(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d2_0.g1 ),
    .A2(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d2_0.a2.out ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d2_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d2_0.o2._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d2_0.o2._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.cg[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d3_0.a1._1_  (.A1(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ),
    .A2(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d3_0.a1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d3_0.a1._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d3_0.a1._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.cp21 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d3_0.a2._1_  (.A1(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d2_0.g1 ),
    .A2(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d3_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d3_0.a2._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d3_0.a2._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d3_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d3_0.o2._1_  (.A1(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d3_0.g1 ),
    .A2(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d3_0.a2.out ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d3_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d3_0.o2._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d3_0.o2._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.cg21 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d3_1.a2._1_  (.A1(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.cg[0] ),
    .A2(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.cp21 ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d3_1.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d3_1.a2._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d3_1.a2._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d3_1.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d3_1.o2._1_  (.A1(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.cg21 ),
    .A2(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d3_1.a2.out ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d3_1.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d3_1.o2._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d3_1.o2._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.cg[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d4_0.a2._1_  (.A1(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.cg[2] ),
    .A2(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d4_0.a2.in0 ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d4_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d4_0.a2._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d4_0.a2._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d4_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d4_0.o2._1_  (.A1(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d4_0.g1 ),
    .A2(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d4_0.a2.out ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d4_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d4_0.o2._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d4_0.o2._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.cg[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d5_0.a1._1_  (.A1(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d4_0.a2.in0 ),
    .A2(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d5_0.a1.in0 ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d5_0.a1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d5_0.a1._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d5_0.a1._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.cp43 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d5_0.a2._1_  (.A1(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d4_0.g1 ),
    .A2(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d5_0.a1.in0 ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d5_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d5_0.a2._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d5_0.a2._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d5_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d5_0.o2._1_  (.A1(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d5_0.g1 ),
    .A2(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d5_0.a2.out ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d5_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d5_0.o2._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d5_0.o2._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.cg43 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d5_1.a2._1_  (.A1(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.cg[2] ),
    .A2(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.cp43 ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d5_1.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d5_1.a2._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d5_1.a2._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d5_1.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d5_1.o2._1_  (.A1(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.cg43 ),
    .A2(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d5_1.a2.out ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d5_1.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d5_1.o2._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d5_1.o2._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.cg[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d6_0.a1._1_  (.A1(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.cp43 ),
    .A2(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d6_0.a1.in0 ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d6_0.a1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d6_0.a1._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d6_0.a1._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.cp54 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d6_0.a2._1_  (.A1(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.cg43 ),
    .A2(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d6_0.a1.in0 ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d6_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d6_0.a2._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d6_0.a2._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d6_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d6_0.o2._1_  (.A1(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d6_0.g1 ),
    .A2(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d6_0.a2.out ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d6_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d6_0.o2._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d6_0.o2._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.cg54 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d6_1.a2._1_  (.A1(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.cg[2] ),
    .A2(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.cp54 ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d6_1.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d6_1.a2._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d6_1.a2._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d6_1.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d6_1.o2._1_  (.A1(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.cg54 ),
    .A2(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d6_1.a2.out ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d6_1.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d6_1.o2._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d6_1.o2._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.cg[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_0.a._1_  (.A1(\mult_add_u0.mult0.step3.add_sub4_u0.int_ip[0] ),
    .A2(\mult_add_u0.mult0.acc_s2[0] ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_0.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_0.a._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_0.a._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d1_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_0.o._1_  (.A1(\mult_add_u0.mult0.step3.add_sub4_u0.int_ip[0] ),
    .A2(\mult_add_u0.mult0.acc_s2[0] ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_0.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_0.o._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_0.o._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d1_0.a2.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_1.a._1_  (.A1(\mult_add_u0.mult0.step3.add_sub4_u0.int_ip[1] ),
    .A2(\mult_add_u0.mult0.acc_s2[1] ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_1.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_1.a._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_1.a._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d2_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_1.o._1_  (.A1(\mult_add_u0.mult0.step3.add_sub4_u0.int_ip[1] ),
    .A2(\mult_add_u0.mult0.acc_s2[1] ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_1.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_1.o._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_1.o._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_2.a._1_  (.A1(\mult_add_u0.mult0.step3.add_sub4_u0.int_ip[2] ),
    .A2(\mult_add_u0.mult0.acc_s2[2] ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_2.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_2.a._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_2.a._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d3_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_2.o._1_  (.A1(\mult_add_u0.mult0.step3.add_sub4_u0.int_ip[2] ),
    .A2(\mult_add_u0.mult0.acc_s2[2] ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_2.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_2.o._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_2.o._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_3.a._1_  (.A1(\mult_add_u0.mult0.step3.add_sub4_u0.int_ip[3] ),
    .A2(\mult_add_u0.mult0.acc_s2[3] ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_3.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_3.a._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_3.a._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d4_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_3.o._1_  (.A1(\mult_add_u0.mult0.step3.add_sub4_u0.int_ip[3] ),
    .A2(\mult_add_u0.mult0.acc_s2[3] ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_3.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_3.o._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_3.o._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d4_0.a2.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_4.a._1_  (.A1(\mult_add_u0.mult0.step3.add_sub4_u0.int_ip[4] ),
    .A2(\mult_add_u0.mult0.acc_s2[4] ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_4.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_4.a._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_4.a._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d5_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_4.o._1_  (.A1(\mult_add_u0.mult0.step3.add_sub4_u0.int_ip[4] ),
    .A2(\mult_add_u0.mult0.acc_s2[4] ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_4.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_4.o._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_4.o._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d5_0.a1.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_5.a._1_  (.A1(\mult_add_u0.mult0.step3.add_sub4_u0.int_ip[5] ),
    .A2(\mult_add_u0.mult0.acc_s2[5] ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_5.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_5.a._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_5.a._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d6_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_5.o._1_  (.A1(\mult_add_u0.mult0.step3.add_sub4_u0.int_ip[5] ),
    .A2(\mult_add_u0.mult0.acc_s2[5] ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_5.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_5.o._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.p_5.o._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.d6_0.a1.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s1.xor2_0._1_  (.A1(\mult_add_u0.mult0.step3.add_sub4_u0.int_ip[1] ),
    .A2(\mult_add_u0.mult0.acc_s2[1] ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s1.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s1.xor2_0._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s1.xor2_0._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s1.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s1.xor2_1._1_  (.A1(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s1.temp ),
    .A2(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.cg[0] ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s1.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s1.xor2_1._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s1.xor2_1._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.S[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s2.xor2_0._1_  (.A1(\mult_add_u0.mult0.step3.add_sub4_u0.int_ip[2] ),
    .A2(\mult_add_u0.mult0.acc_s2[2] ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s2.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s2.xor2_0._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s2.xor2_0._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s2.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s2.xor2_1._1_  (.A1(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s2.temp ),
    .A2(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.cg[1] ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s2.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s2.xor2_1._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s2.xor2_1._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.S[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s3.xor2_0._1_  (.A1(\mult_add_u0.mult0.step3.add_sub4_u0.int_ip[3] ),
    .A2(\mult_add_u0.mult0.acc_s2[3] ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s3.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s3.xor2_0._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s3.xor2_0._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s3.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s3.xor2_1._1_  (.A1(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s3.temp ),
    .A2(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.cg[2] ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s3.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s3.xor2_1._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s3.xor2_1._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.S[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s4.xor2_0._1_  (.A1(\mult_add_u0.mult0.step3.add_sub4_u0.int_ip[4] ),
    .A2(\mult_add_u0.mult0.acc_s2[4] ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s4.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s4.xor2_0._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s4.xor2_0._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s4.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s4.xor2_1._1_  (.A1(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s4.temp ),
    .A2(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.cg[3] ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s4.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s4.xor2_1._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s4.xor2_1._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.S[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s5.xor2_0._1_  (.A1(\mult_add_u0.mult0.step3.add_sub4_u0.int_ip[5] ),
    .A2(\mult_add_u0.mult0.acc_s2[5] ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s5.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s5.xor2_0._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s5.xor2_0._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s5.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s5.xor2_1._1_  (.A1(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s5.temp ),
    .A2(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.cg[4] ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s5.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s5.xor2_1._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s5.xor2_1._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.S[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s6.xor2_0._1_  (.A1(\mult_add_u0.mult0.step3.add_sub4_u0.int_ip[6] ),
    .A2(\mult_add_u0.mult0.acc_s2[6] ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s6.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s6.xor2_0._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s6.xor2_0._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s6.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s6.xor2_1._1_  (.A1(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s6.temp ),
    .A2(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.cg[5] ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s6.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s6.xor2_1._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.s6.xor2_1._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.ppa8_u0.S[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step3.add_sub4_u0.x0._1_  (.A1(\mult_add_u0.mult0.Q_s2[0] ),
    .A2(\mult_add_u0.mult0.multiplicand_s2[0] ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.x0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.x0._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.x0._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.int_ip[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step3.add_sub4_u0.x1._1_  (.A1(\mult_add_u0.mult0.Q_s2[0] ),
    .A2(\mult_add_u0.mult0.multiplicand_s2[1] ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.x1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.x1._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.x1._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.int_ip[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step3.add_sub4_u0.x2._1_  (.A1(\mult_add_u0.mult0.Q_s2[0] ),
    .A2(\mult_add_u0.mult0.multiplicand_s2[2] ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.x2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.x2._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.x2._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.int_ip[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step3.add_sub4_u0.x3._1_  (.A1(\mult_add_u0.mult0.Q_s2[0] ),
    .A2(\mult_add_u0.mult0.multiplicand_s2[3] ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.x3._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.x3._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.x3._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.int_ip[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step3.add_sub4_u0.x4._1_  (.A1(\mult_add_u0.mult0.Q_s2[0] ),
    .A2(\mult_add_u0.mult0.multiplicand_s2[4] ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.x4._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.x4._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.x4._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.int_ip[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step3.add_sub4_u0.x5._1_  (.A1(\mult_add_u0.mult0.Q_s2[0] ),
    .A2(\mult_add_u0.mult0.multiplicand_s2[5] ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.x5._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.x5._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.x5._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.int_ip[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step3.add_sub4_u0.x6._1_  (.A1(\mult_add_u0.mult0.Q_s2[0] ),
    .A2(\mult_add_u0.mult0.multiplicand_s2[6] ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.x6._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step3.add_sub4_u0.x6._2_  (.I(\mult_add_u0.mult0.step3.add_sub4_u0.x6._0_ ),
    .Z(\mult_add_u0.mult0.step3.add_sub4_u0.int_ip[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step4._09_  (.A1(\mult_add_u0.mult0.q0_s3 ),
    .A2(\mult_add_u0.mult0.Q_s3[0] ),
    .Z(\mult_add_u0.mult0.step4._00_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 \mult_add_u0.mult0.step4._10_  (.I(\mult_add_u0.mult0.step4._00_ ),
    .Z(\mult_add_u0.mult0.step4._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.mult0.step4._11_  (.I0(\mult_add_u0.mult0.acc_s3[6] ),
    .I1(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.S[6] ),
    .S(\mult_add_u0.mult0.step4._01_ ),
    .Z(\mult_add_u0.mult0.step4._02_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4._12_  (.I(\mult_add_u0.mult0.step4._02_ ),
    .Z(\mult_add_u0.mult0.acc[4][6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.mult0.step4._13_  (.I0(\mult_add_u0.mult0.acc_s3[1] ),
    .I1(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.S[1] ),
    .S(\mult_add_u0.mult0.step4._01_ ),
    .Z(\mult_add_u0.mult0.step4._03_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4._14_  (.I(\mult_add_u0.mult0.step4._03_ ),
    .Z(\mult_add_u0.mult0.acc[4][0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.mult0.step4._15_  (.I0(\mult_add_u0.mult0.acc_s3[2] ),
    .I1(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.S[2] ),
    .S(\mult_add_u0.mult0.step4._01_ ),
    .Z(\mult_add_u0.mult0.step4._04_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4._16_  (.I(\mult_add_u0.mult0.step4._04_ ),
    .Z(\mult_add_u0.mult0.acc[4][1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.mult0.step4._17_  (.I0(\mult_add_u0.mult0.acc_s3[3] ),
    .I1(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.S[3] ),
    .S(\mult_add_u0.mult0.step4._01_ ),
    .Z(\mult_add_u0.mult0.step4._05_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4._18_  (.I(\mult_add_u0.mult0.step4._05_ ),
    .Z(\mult_add_u0.mult0.acc[4][2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.mult0.step4._19_  (.I0(\mult_add_u0.mult0.acc_s3[4] ),
    .I1(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.S[4] ),
    .S(\mult_add_u0.mult0.step4._01_ ),
    .Z(\mult_add_u0.mult0.step4._06_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4._20_  (.I(\mult_add_u0.mult0.step4._06_ ),
    .Z(\mult_add_u0.mult0.acc[4][3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.mult0.step4._21_  (.I0(\mult_add_u0.mult0.acc_s3[5] ),
    .I1(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.S[5] ),
    .S(\mult_add_u0.mult0.step4._01_ ),
    .Z(\mult_add_u0.mult0.step4._07_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4._22_  (.I(\mult_add_u0.mult0.step4._07_ ),
    .Z(\mult_add_u0.mult0.acc[4][4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.mult0.step4._23_  (.I0(\mult_add_u0.mult0.acc_s3[0] ),
    .I1(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.S[0] ),
    .S(\mult_add_u0.mult0.step4._01_ ),
    .Z(\mult_add_u0.mult0.step4._08_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4._24_  (.I(\mult_add_u0.mult0.step4._08_ ),
    .Z(\mult_add_u0.mult0.Q[3][6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4._25_  (.I(\mult_add_u0.mult0.Q_s3[1] ),
    .Z(\mult_add_u0.mult0.Q[3][0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4._26_  (.I(\mult_add_u0.mult0.Q_s3[2] ),
    .Z(\mult_add_u0.mult0.Q[3][1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4._27_  (.I(\mult_add_u0.mult0.Q_s3[3] ),
    .Z(\mult_add_u0.mult0.Q[3][2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4._31_  (.I(\mult_add_u0.mult0.acc[4][6] ),
    .Z(\mult_add_u0.mult0.acc[4][5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4._32_  (.I(\mult_add_u0.mult0.Q_s3[0] ),
    .Z(\mult_add_u0.mult0.q0[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d1_0.a2._1_  (.A1(\mult_add_u0.mult0.Q_s3[0] ),
    .A2(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d1_0.a2.in0 ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d1_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d1_0.a2._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d1_0.a2._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d1_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d1_0.o2._1_  (.A1(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d1_0.g1 ),
    .A2(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d1_0.a2.out ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d1_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d1_0.o2._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d1_0.o2._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.cg[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d2_0.a2._1_  (.A1(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.cg[0] ),
    .A2(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d2_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d2_0.a2._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d2_0.a2._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d2_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d2_0.o2._1_  (.A1(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d2_0.g1 ),
    .A2(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d2_0.a2.out ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d2_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d2_0.o2._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d2_0.o2._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.cg[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d3_0.a1._1_  (.A1(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ),
    .A2(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d3_0.a1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d3_0.a1._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d3_0.a1._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.cp21 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d3_0.a2._1_  (.A1(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d2_0.g1 ),
    .A2(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d3_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d3_0.a2._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d3_0.a2._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d3_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d3_0.o2._1_  (.A1(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d3_0.g1 ),
    .A2(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d3_0.a2.out ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d3_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d3_0.o2._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d3_0.o2._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.cg21 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d3_1.a2._1_  (.A1(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.cg[0] ),
    .A2(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.cp21 ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d3_1.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d3_1.a2._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d3_1.a2._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d3_1.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d3_1.o2._1_  (.A1(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.cg21 ),
    .A2(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d3_1.a2.out ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d3_1.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d3_1.o2._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d3_1.o2._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.cg[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d4_0.a2._1_  (.A1(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.cg[2] ),
    .A2(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d4_0.a2.in0 ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d4_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d4_0.a2._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d4_0.a2._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d4_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d4_0.o2._1_  (.A1(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d4_0.g1 ),
    .A2(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d4_0.a2.out ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d4_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d4_0.o2._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d4_0.o2._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.cg[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d5_0.a1._1_  (.A1(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d4_0.a2.in0 ),
    .A2(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d5_0.a1.in0 ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d5_0.a1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d5_0.a1._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d5_0.a1._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.cp43 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d5_0.a2._1_  (.A1(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d4_0.g1 ),
    .A2(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d5_0.a1.in0 ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d5_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d5_0.a2._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d5_0.a2._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d5_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d5_0.o2._1_  (.A1(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d5_0.g1 ),
    .A2(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d5_0.a2.out ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d5_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d5_0.o2._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d5_0.o2._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.cg43 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d5_1.a2._1_  (.A1(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.cg[2] ),
    .A2(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.cp43 ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d5_1.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d5_1.a2._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d5_1.a2._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d5_1.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d5_1.o2._1_  (.A1(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.cg43 ),
    .A2(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d5_1.a2.out ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d5_1.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d5_1.o2._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d5_1.o2._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.cg[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d6_0.a1._1_  (.A1(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.cp43 ),
    .A2(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d6_0.a1.in0 ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d6_0.a1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d6_0.a1._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d6_0.a1._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.cp54 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d6_0.a2._1_  (.A1(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.cg43 ),
    .A2(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d6_0.a1.in0 ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d6_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d6_0.a2._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d6_0.a2._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d6_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d6_0.o2._1_  (.A1(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d6_0.g1 ),
    .A2(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d6_0.a2.out ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d6_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d6_0.o2._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d6_0.o2._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.cg54 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d6_1.a2._1_  (.A1(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.cg[2] ),
    .A2(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.cp54 ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d6_1.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d6_1.a2._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d6_1.a2._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d6_1.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d6_1.o2._1_  (.A1(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.cg54 ),
    .A2(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d6_1.a2.out ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d6_1.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d6_1.o2._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d6_1.o2._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.cg[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_0.a._1_  (.A1(\mult_add_u0.mult0.step4.add_sub4_u0.int_ip[0] ),
    .A2(\mult_add_u0.mult0.acc_s3[0] ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_0.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_0.a._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_0.a._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d1_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_0.o._1_  (.A1(\mult_add_u0.mult0.step4.add_sub4_u0.int_ip[0] ),
    .A2(\mult_add_u0.mult0.acc_s3[0] ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_0.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_0.o._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_0.o._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d1_0.a2.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_1.a._1_  (.A1(\mult_add_u0.mult0.step4.add_sub4_u0.int_ip[1] ),
    .A2(\mult_add_u0.mult0.acc_s3[1] ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_1.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_1.a._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_1.a._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d2_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_1.o._1_  (.A1(\mult_add_u0.mult0.step4.add_sub4_u0.int_ip[1] ),
    .A2(\mult_add_u0.mult0.acc_s3[1] ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_1.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_1.o._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_1.o._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_2.a._1_  (.A1(\mult_add_u0.mult0.step4.add_sub4_u0.int_ip[2] ),
    .A2(\mult_add_u0.mult0.acc_s3[2] ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_2.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_2.a._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_2.a._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d3_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_2.o._1_  (.A1(\mult_add_u0.mult0.step4.add_sub4_u0.int_ip[2] ),
    .A2(\mult_add_u0.mult0.acc_s3[2] ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_2.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_2.o._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_2.o._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_3.a._1_  (.A1(\mult_add_u0.mult0.step4.add_sub4_u0.int_ip[3] ),
    .A2(\mult_add_u0.mult0.acc_s3[3] ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_3.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_3.a._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_3.a._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d4_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_3.o._1_  (.A1(\mult_add_u0.mult0.step4.add_sub4_u0.int_ip[3] ),
    .A2(\mult_add_u0.mult0.acc_s3[3] ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_3.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_3.o._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_3.o._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d4_0.a2.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_4.a._1_  (.A1(\mult_add_u0.mult0.step4.add_sub4_u0.int_ip[4] ),
    .A2(\mult_add_u0.mult0.acc_s3[4] ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_4.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_4.a._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_4.a._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d5_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_4.o._1_  (.A1(\mult_add_u0.mult0.step4.add_sub4_u0.int_ip[4] ),
    .A2(\mult_add_u0.mult0.acc_s3[4] ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_4.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_4.o._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_4.o._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d5_0.a1.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_5.a._1_  (.A1(\mult_add_u0.mult0.step4.add_sub4_u0.int_ip[5] ),
    .A2(\mult_add_u0.mult0.acc_s3[5] ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_5.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_5.a._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_5.a._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d6_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_5.o._1_  (.A1(\mult_add_u0.mult0.step4.add_sub4_u0.int_ip[5] ),
    .A2(\mult_add_u0.mult0.acc_s3[5] ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_5.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_5.o._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.p_5.o._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.d6_0.a1.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s0.xor2_0._1_  (.A1(\mult_add_u0.mult0.step4.add_sub4_u0.int_ip[0] ),
    .A2(\mult_add_u0.mult0.acc_s3[0] ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s0.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s0.xor2_0._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s0.xor2_0._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s0.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s0.xor2_1._1_  (.A1(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s0.temp ),
    .A2(\mult_add_u0.mult0.Q_s3[0] ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s0.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s0.xor2_1._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s0.xor2_1._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.S[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s1.xor2_0._1_  (.A1(\mult_add_u0.mult0.step4.add_sub4_u0.int_ip[1] ),
    .A2(\mult_add_u0.mult0.acc_s3[1] ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s1.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s1.xor2_0._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s1.xor2_0._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s1.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s1.xor2_1._1_  (.A1(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s1.temp ),
    .A2(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.cg[0] ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s1.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s1.xor2_1._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s1.xor2_1._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.S[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s2.xor2_0._1_  (.A1(\mult_add_u0.mult0.step4.add_sub4_u0.int_ip[2] ),
    .A2(\mult_add_u0.mult0.acc_s3[2] ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s2.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s2.xor2_0._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s2.xor2_0._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s2.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s2.xor2_1._1_  (.A1(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s2.temp ),
    .A2(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.cg[1] ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s2.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s2.xor2_1._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s2.xor2_1._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.S[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s3.xor2_0._1_  (.A1(\mult_add_u0.mult0.step4.add_sub4_u0.int_ip[3] ),
    .A2(\mult_add_u0.mult0.acc_s3[3] ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s3.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s3.xor2_0._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s3.xor2_0._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s3.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s3.xor2_1._1_  (.A1(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s3.temp ),
    .A2(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.cg[2] ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s3.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s3.xor2_1._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s3.xor2_1._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.S[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s4.xor2_0._1_  (.A1(\mult_add_u0.mult0.step4.add_sub4_u0.int_ip[4] ),
    .A2(\mult_add_u0.mult0.acc_s3[4] ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s4.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s4.xor2_0._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s4.xor2_0._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s4.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s4.xor2_1._1_  (.A1(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s4.temp ),
    .A2(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.cg[3] ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s4.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s4.xor2_1._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s4.xor2_1._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.S[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s5.xor2_0._1_  (.A1(\mult_add_u0.mult0.step4.add_sub4_u0.int_ip[5] ),
    .A2(\mult_add_u0.mult0.acc_s3[5] ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s5.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s5.xor2_0._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s5.xor2_0._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s5.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s5.xor2_1._1_  (.A1(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s5.temp ),
    .A2(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.cg[4] ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s5.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s5.xor2_1._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s5.xor2_1._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.S[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s6.xor2_0._1_  (.A1(\mult_add_u0.mult0.step4.add_sub4_u0.int_ip[6] ),
    .A2(\mult_add_u0.mult0.acc_s3[6] ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s6.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s6.xor2_0._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s6.xor2_0._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s6.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s6.xor2_1._1_  (.A1(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s6.temp ),
    .A2(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.cg[5] ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s6.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s6.xor2_1._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.s6.xor2_1._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.ppa8_u0.S[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step4.add_sub4_u0.x0._1_  (.A1(\mult_add_u0.mult0.Q_s3[0] ),
    .A2(\mult_add_u0.mult0.multiplicand_s3[0] ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.x0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.x0._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.x0._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.int_ip[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step4.add_sub4_u0.x1._1_  (.A1(\mult_add_u0.mult0.Q_s3[0] ),
    .A2(\mult_add_u0.mult0.multiplicand_s3[1] ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.x1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.x1._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.x1._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.int_ip[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step4.add_sub4_u0.x2._1_  (.A1(\mult_add_u0.mult0.Q_s3[0] ),
    .A2(\mult_add_u0.mult0.multiplicand_s3[2] ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.x2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.x2._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.x2._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.int_ip[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step4.add_sub4_u0.x3._1_  (.A1(\mult_add_u0.mult0.Q_s3[0] ),
    .A2(\mult_add_u0.mult0.multiplicand_s3[3] ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.x3._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.x3._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.x3._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.int_ip[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step4.add_sub4_u0.x4._1_  (.A1(\mult_add_u0.mult0.Q_s3[0] ),
    .A2(\mult_add_u0.mult0.multiplicand_s3[4] ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.x4._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.x4._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.x4._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.int_ip[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step4.add_sub4_u0.x5._1_  (.A1(\mult_add_u0.mult0.Q_s3[0] ),
    .A2(\mult_add_u0.mult0.multiplicand_s3[5] ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.x5._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.x5._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.x5._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.int_ip[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step4.add_sub4_u0.x6._1_  (.A1(\mult_add_u0.mult0.Q_s3[0] ),
    .A2(\mult_add_u0.mult0.multiplicand_s3[6] ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.x6._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step4.add_sub4_u0.x6._2_  (.I(\mult_add_u0.mult0.step4.add_sub4_u0.x6._0_ ),
    .Z(\mult_add_u0.mult0.step4.add_sub4_u0.int_ip[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step5._09_  (.A1(\mult_add_u0.mult0.q0_s4 ),
    .A2(\mult_add_u0.mult0.Q_s4[0] ),
    .Z(\mult_add_u0.mult0.step5._00_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 \mult_add_u0.mult0.step5._10_  (.I(\mult_add_u0.mult0.step5._00_ ),
    .Z(\mult_add_u0.mult0.step5._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.mult0.step5._13_  (.I0(\mult_add_u0.mult0.acc_s4[1] ),
    .I1(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.S[1] ),
    .S(\mult_add_u0.mult0.step5._01_ ),
    .Z(\mult_add_u0.mult0.step5._03_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5._14_  (.I(\mult_add_u0.mult0.step5._03_ ),
    .Z(\mult_add_u0.mult0.acc[5][0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.mult0.step5._15_  (.I0(\mult_add_u0.mult0.acc_s4[2] ),
    .I1(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.S[2] ),
    .S(\mult_add_u0.mult0.step5._01_ ),
    .Z(\mult_add_u0.mult0.step5._04_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5._16_  (.I(\mult_add_u0.mult0.step5._04_ ),
    .Z(\mult_add_u0.mult0.acc[5][1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.mult0.step5._17_  (.I0(\mult_add_u0.mult0.acc_s4[3] ),
    .I1(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.S[3] ),
    .S(\mult_add_u0.mult0.step5._01_ ),
    .Z(\mult_add_u0.mult0.step5._05_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5._18_  (.I(\mult_add_u0.mult0.step5._05_ ),
    .Z(\mult_add_u0.mult0.acc[5][2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.mult0.step5._19_  (.I0(\mult_add_u0.mult0.acc_s4[4] ),
    .I1(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.S[4] ),
    .S(\mult_add_u0.mult0.step5._01_ ),
    .Z(\mult_add_u0.mult0.step5._06_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5._20_  (.I(\mult_add_u0.mult0.step5._06_ ),
    .Z(\mult_add_u0.mult0.acc[5][3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.mult0.step5._21_  (.I0(\mult_add_u0.mult0.acc_s4[5] ),
    .I1(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.S[5] ),
    .S(\mult_add_u0.mult0.step5._01_ ),
    .Z(\mult_add_u0.mult0.step5._07_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5._22_  (.I(\mult_add_u0.mult0.step5._07_ ),
    .Z(\mult_add_u0.mult0.acc[5][4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.mult0.step5._23_  (.I0(\mult_add_u0.mult0.acc_s4[0] ),
    .I1(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.S[0] ),
    .S(\mult_add_u0.mult0.step5._01_ ),
    .Z(\mult_add_u0.mult0.step5._08_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5._24_  (.I(\mult_add_u0.mult0.step5._08_ ),
    .Z(\mult_add_u0.mult0.Q[4][6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5._25_  (.I(\mult_add_u0.mult0.Q_s4[1] ),
    .Z(\mult_add_u0.mult0.Q[4][0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5._26_  (.I(\mult_add_u0.mult0.Q_s4[2] ),
    .Z(\mult_add_u0.mult0.Q[4][1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5._30_  (.I(\mult_add_u0.mult0.Q_s4[6] ),
    .Z(\mult_add_u0.mult0.Q[4][5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5._32_  (.I(\mult_add_u0.mult0.Q_s4[0] ),
    .Z(\mult_add_u0.mult0.q0[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d1_0.a2._1_  (.A1(\mult_add_u0.mult0.Q_s4[0] ),
    .A2(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d1_0.a2.in0 ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d1_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d1_0.a2._2_  (.I(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d1_0.a2._0_ ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d1_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d1_0.o2._1_  (.A1(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d1_0.g1 ),
    .A2(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d1_0.a2.out ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d1_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d1_0.o2._2_  (.I(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d1_0.o2._0_ ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.cg[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d2_0.a2._1_  (.A1(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.cg[0] ),
    .A2(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d2_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d2_0.a2._2_  (.I(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d2_0.a2._0_ ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d2_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d2_0.o2._1_  (.A1(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d2_0.g1 ),
    .A2(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d2_0.a2.out ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d2_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d2_0.o2._2_  (.I(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d2_0.o2._0_ ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.cg[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d3_0.a1._1_  (.A1(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ),
    .A2(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d3_0.a1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d3_0.a1._2_  (.I(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d3_0.a1._0_ ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.cp21 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d3_0.a2._1_  (.A1(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d2_0.g1 ),
    .A2(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d3_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d3_0.a2._2_  (.I(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d3_0.a2._0_ ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d3_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d3_0.o2._1_  (.A1(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d3_0.g1 ),
    .A2(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d3_0.a2.out ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d3_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d3_0.o2._2_  (.I(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d3_0.o2._0_ ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.cg21 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d3_1.a2._1_  (.A1(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.cg[0] ),
    .A2(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.cp21 ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d3_1.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d3_1.a2._2_  (.I(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d3_1.a2._0_ ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d3_1.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d3_1.o2._1_  (.A1(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.cg21 ),
    .A2(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d3_1.a2.out ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d3_1.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d3_1.o2._2_  (.I(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d3_1.o2._0_ ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.cg[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d4_0.a2._1_  (.A1(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.cg[2] ),
    .A2(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d4_0.a2.in0 ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d4_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d4_0.a2._2_  (.I(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d4_0.a2._0_ ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d4_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d4_0.o2._1_  (.A1(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d4_0.g1 ),
    .A2(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d4_0.a2.out ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d4_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d4_0.o2._2_  (.I(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d4_0.o2._0_ ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.cg[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d5_0.a1._1_  (.A1(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d4_0.a2.in0 ),
    .A2(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d5_0.a1.in0 ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d5_0.a1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d5_0.a1._2_  (.I(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d5_0.a1._0_ ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.cp43 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d5_0.a2._1_  (.A1(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d4_0.g1 ),
    .A2(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d5_0.a1.in0 ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d5_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d5_0.a2._2_  (.I(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d5_0.a2._0_ ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d5_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d5_0.o2._1_  (.A1(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d5_0.g1 ),
    .A2(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d5_0.a2.out ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d5_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d5_0.o2._2_  (.I(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d5_0.o2._0_ ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.cg43 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d5_1.a2._1_  (.A1(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.cg[2] ),
    .A2(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.cp43 ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d5_1.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d5_1.a2._2_  (.I(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d5_1.a2._0_ ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d5_1.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d5_1.o2._1_  (.A1(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.cg43 ),
    .A2(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d5_1.a2.out ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d5_1.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d5_1.o2._2_  (.I(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d5_1.o2._0_ ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.cg[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_0.a._1_  (.A1(\mult_add_u0.mult0.step5.add_sub4_u0.int_ip[0] ),
    .A2(\mult_add_u0.mult0.acc_s4[0] ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_0.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_0.a._2_  (.I(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_0.a._0_ ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d1_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_0.o._1_  (.A1(\mult_add_u0.mult0.step5.add_sub4_u0.int_ip[0] ),
    .A2(\mult_add_u0.mult0.acc_s4[0] ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_0.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_0.o._2_  (.I(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_0.o._0_ ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d1_0.a2.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_1.a._1_  (.A1(\mult_add_u0.mult0.step5.add_sub4_u0.int_ip[1] ),
    .A2(\mult_add_u0.mult0.acc_s4[1] ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_1.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_1.a._2_  (.I(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_1.a._0_ ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d2_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_1.o._1_  (.A1(\mult_add_u0.mult0.step5.add_sub4_u0.int_ip[1] ),
    .A2(\mult_add_u0.mult0.acc_s4[1] ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_1.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_1.o._2_  (.I(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_1.o._0_ ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_2.a._1_  (.A1(\mult_add_u0.mult0.step5.add_sub4_u0.int_ip[2] ),
    .A2(\mult_add_u0.mult0.acc_s4[2] ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_2.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_2.a._2_  (.I(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_2.a._0_ ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d3_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_2.o._1_  (.A1(\mult_add_u0.mult0.step5.add_sub4_u0.int_ip[2] ),
    .A2(\mult_add_u0.mult0.acc_s4[2] ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_2.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_2.o._2_  (.I(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_2.o._0_ ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_3.a._1_  (.A1(\mult_add_u0.mult0.step5.add_sub4_u0.int_ip[3] ),
    .A2(\mult_add_u0.mult0.acc_s4[3] ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_3.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_3.a._2_  (.I(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_3.a._0_ ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d4_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_3.o._1_  (.A1(\mult_add_u0.mult0.step5.add_sub4_u0.int_ip[3] ),
    .A2(\mult_add_u0.mult0.acc_s4[3] ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_3.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_3.o._2_  (.I(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_3.o._0_ ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d4_0.a2.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_4.a._1_  (.A1(\mult_add_u0.mult0.step5.add_sub4_u0.int_ip[4] ),
    .A2(\mult_add_u0.mult0.acc_s4[4] ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_4.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_4.a._2_  (.I(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_4.a._0_ ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d5_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_4.o._1_  (.A1(\mult_add_u0.mult0.step5.add_sub4_u0.int_ip[4] ),
    .A2(\mult_add_u0.mult0.acc_s4[4] ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_4.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_4.o._2_  (.I(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.p_4.o._0_ ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.d5_0.a1.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s0.xor2_0._1_  (.A1(\mult_add_u0.mult0.step5.add_sub4_u0.int_ip[0] ),
    .A2(\mult_add_u0.mult0.acc_s4[0] ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s0.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s0.xor2_0._2_  (.I(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s0.xor2_0._0_ ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s0.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s0.xor2_1._1_  (.A1(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s0.temp ),
    .A2(\mult_add_u0.mult0.Q_s4[0] ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s0.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s0.xor2_1._2_  (.I(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s0.xor2_1._0_ ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.S[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s1.xor2_0._1_  (.A1(\mult_add_u0.mult0.step5.add_sub4_u0.int_ip[1] ),
    .A2(\mult_add_u0.mult0.acc_s4[1] ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s1.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s1.xor2_0._2_  (.I(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s1.xor2_0._0_ ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s1.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s1.xor2_1._1_  (.A1(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s1.temp ),
    .A2(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.cg[0] ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s1.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s1.xor2_1._2_  (.I(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s1.xor2_1._0_ ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.S[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s2.xor2_0._1_  (.A1(\mult_add_u0.mult0.step5.add_sub4_u0.int_ip[2] ),
    .A2(\mult_add_u0.mult0.acc_s4[2] ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s2.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s2.xor2_0._2_  (.I(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s2.xor2_0._0_ ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s2.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s2.xor2_1._1_  (.A1(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s2.temp ),
    .A2(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.cg[1] ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s2.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s2.xor2_1._2_  (.I(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s2.xor2_1._0_ ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.S[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s3.xor2_0._1_  (.A1(\mult_add_u0.mult0.step5.add_sub4_u0.int_ip[3] ),
    .A2(\mult_add_u0.mult0.acc_s4[3] ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s3.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s3.xor2_0._2_  (.I(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s3.xor2_0._0_ ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s3.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s3.xor2_1._1_  (.A1(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s3.temp ),
    .A2(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.cg[2] ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s3.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s3.xor2_1._2_  (.I(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s3.xor2_1._0_ ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.S[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s4.xor2_0._1_  (.A1(\mult_add_u0.mult0.step5.add_sub4_u0.int_ip[4] ),
    .A2(\mult_add_u0.mult0.acc_s4[4] ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s4.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s4.xor2_0._2_  (.I(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s4.xor2_0._0_ ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s4.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s4.xor2_1._1_  (.A1(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s4.temp ),
    .A2(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.cg[3] ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s4.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s4.xor2_1._2_  (.I(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s4.xor2_1._0_ ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.S[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s5.xor2_0._1_  (.A1(\mult_add_u0.mult0.step5.add_sub4_u0.int_ip[5] ),
    .A2(\mult_add_u0.mult0.acc_s4[5] ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s5.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s5.xor2_0._2_  (.I(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s5.xor2_0._0_ ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s5.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s5.xor2_1._1_  (.A1(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s5.temp ),
    .A2(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.cg[4] ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s5.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s5.xor2_1._2_  (.I(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.s5.xor2_1._0_ ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.ppa8_u0.S[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step5.add_sub4_u0.x0._1_  (.A1(\mult_add_u0.mult0.Q_s4[0] ),
    .A2(\mult_add_u0.mult0.multiplicand_s4[0] ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.x0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5.add_sub4_u0.x0._2_  (.I(\mult_add_u0.mult0.step5.add_sub4_u0.x0._0_ ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.int_ip[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step5.add_sub4_u0.x1._1_  (.A1(\mult_add_u0.mult0.Q_s4[0] ),
    .A2(\mult_add_u0.mult0.multiplicand_s4[1] ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.x1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5.add_sub4_u0.x1._2_  (.I(\mult_add_u0.mult0.step5.add_sub4_u0.x1._0_ ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.int_ip[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step5.add_sub4_u0.x2._1_  (.A1(\mult_add_u0.mult0.Q_s4[0] ),
    .A2(\mult_add_u0.mult0.multiplicand_s4[2] ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.x2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5.add_sub4_u0.x2._2_  (.I(\mult_add_u0.mult0.step5.add_sub4_u0.x2._0_ ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.int_ip[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step5.add_sub4_u0.x3._1_  (.A1(\mult_add_u0.mult0.Q_s4[0] ),
    .A2(\mult_add_u0.mult0.multiplicand_s4[3] ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.x3._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5.add_sub4_u0.x3._2_  (.I(\mult_add_u0.mult0.step5.add_sub4_u0.x3._0_ ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.int_ip[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step5.add_sub4_u0.x4._1_  (.A1(\mult_add_u0.mult0.Q_s4[0] ),
    .A2(\mult_add_u0.mult0.multiplicand_s4[4] ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.x4._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5.add_sub4_u0.x4._2_  (.I(\mult_add_u0.mult0.step5.add_sub4_u0.x4._0_ ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.int_ip[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step5.add_sub4_u0.x5._1_  (.A1(\mult_add_u0.mult0.Q_s4[0] ),
    .A2(\mult_add_u0.mult0.multiplicand_s4[5] ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.x5._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step5.add_sub4_u0.x5._2_  (.I(\mult_add_u0.mult0.step5.add_sub4_u0.x5._0_ ),
    .Z(\mult_add_u0.mult0.step5.add_sub4_u0.int_ip[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step6._09_  (.A1(\mult_add_u0.mult0.q0_s5 ),
    .A2(\mult_add_u0.mult0.Q_s5[0] ),
    .Z(\mult_add_u0.mult0.step6._00_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 \mult_add_u0.mult0.step6._10_  (.I(\mult_add_u0.mult0.step6._00_ ),
    .Z(\mult_add_u0.mult0.step6._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.mult0.step6._13_  (.I0(\mult_add_u0.mult0.acc_s5[1] ),
    .I1(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.S[1] ),
    .S(\mult_add_u0.mult0.step6._01_ ),
    .Z(\mult_add_u0.mult0.step6._03_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step6._14_  (.I(\mult_add_u0.mult0.step6._03_ ),
    .Z(\mult_add_u0.mult0.acc[6][0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.mult0.step6._15_  (.I0(\mult_add_u0.mult0.acc_s5[2] ),
    .I1(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.S[2] ),
    .S(\mult_add_u0.mult0.step6._01_ ),
    .Z(\mult_add_u0.mult0.step6._04_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step6._16_  (.I(\mult_add_u0.mult0.step6._04_ ),
    .Z(\mult_add_u0.mult0.acc[6][1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.mult0.step6._17_  (.I0(\mult_add_u0.mult0.acc_s5[3] ),
    .I1(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.S[3] ),
    .S(\mult_add_u0.mult0.step6._01_ ),
    .Z(\mult_add_u0.mult0.step6._05_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step6._18_  (.I(\mult_add_u0.mult0.step6._05_ ),
    .Z(\mult_add_u0.mult0.acc[6][2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.mult0.step6._19_  (.I0(\mult_add_u0.mult0.acc_s5[4] ),
    .I1(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.S[4] ),
    .S(\mult_add_u0.mult0.step6._01_ ),
    .Z(\mult_add_u0.mult0.step6._06_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step6._20_  (.I(\mult_add_u0.mult0.step6._06_ ),
    .Z(\mult_add_u0.mult0.acc[6][3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.mult0.step6._23_  (.I0(\mult_add_u0.mult0.acc_s5[0] ),
    .I1(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.S[0] ),
    .S(\mult_add_u0.mult0.step6._01_ ),
    .Z(\mult_add_u0.mult0.step6._08_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step6._24_  (.I(\mult_add_u0.mult0.step6._08_ ),
    .Z(\mult_add_u0.mult0.Q[5][6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step6._25_  (.I(\mult_add_u0.mult0.Q_s5[1] ),
    .Z(\mult_add_u0.mult0.Q[5][0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step6._29_  (.I(\mult_add_u0.mult0.Q_s5[5] ),
    .Z(\mult_add_u0.mult0.Q[5][4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step6._30_  (.I(\mult_add_u0.mult0.Q_s5[6] ),
    .Z(\mult_add_u0.mult0.Q[5][5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step6._32_  (.I(\mult_add_u0.mult0.Q_s5[0] ),
    .Z(\mult_add_u0.mult0.q0[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d1_0.a2._1_  (.A1(\mult_add_u0.mult0.Q_s5[0] ),
    .A2(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d1_0.a2.in0 ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d1_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d1_0.a2._2_  (.I(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d1_0.a2._0_ ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d1_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d1_0.o2._1_  (.A1(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d1_0.g1 ),
    .A2(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d1_0.a2.out ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d1_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d1_0.o2._2_  (.I(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d1_0.o2._0_ ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.cg[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d2_0.a2._1_  (.A1(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.cg[0] ),
    .A2(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d2_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d2_0.a2._2_  (.I(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d2_0.a2._0_ ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d2_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d2_0.o2._1_  (.A1(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d2_0.g1 ),
    .A2(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d2_0.a2.out ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d2_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d2_0.o2._2_  (.I(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d2_0.o2._0_ ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.cg[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d3_0.a1._1_  (.A1(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ),
    .A2(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d3_0.a1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d3_0.a1._2_  (.I(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d3_0.a1._0_ ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.cp21 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d3_0.a2._1_  (.A1(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d2_0.g1 ),
    .A2(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d3_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d3_0.a2._2_  (.I(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d3_0.a2._0_ ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d3_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d3_0.o2._1_  (.A1(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d3_0.g1 ),
    .A2(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d3_0.a2.out ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d3_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d3_0.o2._2_  (.I(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d3_0.o2._0_ ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.cg21 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d3_1.a2._1_  (.A1(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.cg[0] ),
    .A2(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.cp21 ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d3_1.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d3_1.a2._2_  (.I(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d3_1.a2._0_ ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d3_1.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d3_1.o2._1_  (.A1(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.cg21 ),
    .A2(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d3_1.a2.out ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d3_1.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d3_1.o2._2_  (.I(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d3_1.o2._0_ ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.cg[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d4_0.a2._1_  (.A1(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.cg[2] ),
    .A2(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d4_0.a2.in0 ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d4_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d4_0.a2._2_  (.I(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d4_0.a2._0_ ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d4_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d4_0.o2._1_  (.A1(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d4_0.g1 ),
    .A2(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d4_0.a2.out ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d4_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d4_0.o2._2_  (.I(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d4_0.o2._0_ ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.cg[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.p_0.a._1_  (.A1(\mult_add_u0.mult0.step6.add_sub4_u0.int_ip[0] ),
    .A2(\mult_add_u0.mult0.acc_s5[0] ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.p_0.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.p_0.a._2_  (.I(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.p_0.a._0_ ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d1_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.p_0.o._1_  (.A1(\mult_add_u0.mult0.step6.add_sub4_u0.int_ip[0] ),
    .A2(\mult_add_u0.mult0.acc_s5[0] ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.p_0.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.p_0.o._2_  (.I(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.p_0.o._0_ ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d1_0.a2.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.p_1.a._1_  (.A1(\mult_add_u0.mult0.step6.add_sub4_u0.int_ip[1] ),
    .A2(\mult_add_u0.mult0.acc_s5[1] ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.p_1.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.p_1.a._2_  (.I(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.p_1.a._0_ ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d2_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.p_1.o._1_  (.A1(\mult_add_u0.mult0.step6.add_sub4_u0.int_ip[1] ),
    .A2(\mult_add_u0.mult0.acc_s5[1] ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.p_1.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.p_1.o._2_  (.I(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.p_1.o._0_ ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.p_2.a._1_  (.A1(\mult_add_u0.mult0.step6.add_sub4_u0.int_ip[2] ),
    .A2(\mult_add_u0.mult0.acc_s5[2] ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.p_2.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.p_2.a._2_  (.I(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.p_2.a._0_ ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d3_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.p_2.o._1_  (.A1(\mult_add_u0.mult0.step6.add_sub4_u0.int_ip[2] ),
    .A2(\mult_add_u0.mult0.acc_s5[2] ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.p_2.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.p_2.o._2_  (.I(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.p_2.o._0_ ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.p_3.a._1_  (.A1(\mult_add_u0.mult0.step6.add_sub4_u0.int_ip[3] ),
    .A2(\mult_add_u0.mult0.acc_s5[3] ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.p_3.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.p_3.a._2_  (.I(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.p_3.a._0_ ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d4_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.p_3.o._1_  (.A1(\mult_add_u0.mult0.step6.add_sub4_u0.int_ip[3] ),
    .A2(\mult_add_u0.mult0.acc_s5[3] ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.p_3.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.p_3.o._2_  (.I(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.p_3.o._0_ ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.d4_0.a2.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s0.xor2_0._1_  (.A1(\mult_add_u0.mult0.step6.add_sub4_u0.int_ip[0] ),
    .A2(\mult_add_u0.mult0.acc_s5[0] ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s0.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s0.xor2_0._2_  (.I(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s0.xor2_0._0_ ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s0.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s0.xor2_1._1_  (.A1(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s0.temp ),
    .A2(\mult_add_u0.mult0.Q_s5[0] ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s0.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s0.xor2_1._2_  (.I(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s0.xor2_1._0_ ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.S[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s1.xor2_0._1_  (.A1(\mult_add_u0.mult0.step6.add_sub4_u0.int_ip[1] ),
    .A2(\mult_add_u0.mult0.acc_s5[1] ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s1.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s1.xor2_0._2_  (.I(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s1.xor2_0._0_ ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s1.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s1.xor2_1._1_  (.A1(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s1.temp ),
    .A2(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.cg[0] ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s1.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s1.xor2_1._2_  (.I(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s1.xor2_1._0_ ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.S[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s2.xor2_0._1_  (.A1(\mult_add_u0.mult0.step6.add_sub4_u0.int_ip[2] ),
    .A2(\mult_add_u0.mult0.acc_s5[2] ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s2.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s2.xor2_0._2_  (.I(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s2.xor2_0._0_ ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s2.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s2.xor2_1._1_  (.A1(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s2.temp ),
    .A2(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.cg[1] ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s2.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s2.xor2_1._2_  (.I(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s2.xor2_1._0_ ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.S[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s3.xor2_0._1_  (.A1(\mult_add_u0.mult0.step6.add_sub4_u0.int_ip[3] ),
    .A2(\mult_add_u0.mult0.acc_s5[3] ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s3.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s3.xor2_0._2_  (.I(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s3.xor2_0._0_ ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s3.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s3.xor2_1._1_  (.A1(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s3.temp ),
    .A2(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.cg[2] ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s3.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s3.xor2_1._2_  (.I(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s3.xor2_1._0_ ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.S[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s4.xor2_0._1_  (.A1(\mult_add_u0.mult0.step6.add_sub4_u0.int_ip[4] ),
    .A2(\mult_add_u0.mult0.acc_s5[4] ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s4.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s4.xor2_0._2_  (.I(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s4.xor2_0._0_ ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s4.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s4.xor2_1._1_  (.A1(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s4.temp ),
    .A2(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.cg[3] ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s4.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s4.xor2_1._2_  (.I(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.s4.xor2_1._0_ ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.ppa8_u0.S[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step6.add_sub4_u0.x0._1_  (.A1(\mult_add_u0.mult0.Q_s5[0] ),
    .A2(\mult_add_u0.mult0.multiplicand_s5[0] ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.x0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step6.add_sub4_u0.x0._2_  (.I(\mult_add_u0.mult0.step6.add_sub4_u0.x0._0_ ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.int_ip[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step6.add_sub4_u0.x1._1_  (.A1(\mult_add_u0.mult0.Q_s5[0] ),
    .A2(\mult_add_u0.mult0.multiplicand_s5[1] ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.x1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step6.add_sub4_u0.x1._2_  (.I(\mult_add_u0.mult0.step6.add_sub4_u0.x1._0_ ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.int_ip[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step6.add_sub4_u0.x2._1_  (.A1(\mult_add_u0.mult0.Q_s5[0] ),
    .A2(\mult_add_u0.mult0.multiplicand_s5[2] ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.x2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step6.add_sub4_u0.x2._2_  (.I(\mult_add_u0.mult0.step6.add_sub4_u0.x2._0_ ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.int_ip[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step6.add_sub4_u0.x3._1_  (.A1(\mult_add_u0.mult0.Q_s5[0] ),
    .A2(\mult_add_u0.mult0.multiplicand_s5[3] ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.x3._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step6.add_sub4_u0.x3._2_  (.I(\mult_add_u0.mult0.step6.add_sub4_u0.x3._0_ ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.int_ip[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step6.add_sub4_u0.x4._1_  (.A1(\mult_add_u0.mult0.Q_s5[0] ),
    .A2(\mult_add_u0.mult0.multiplicand_s5[4] ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.x4._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step6.add_sub4_u0.x4._2_  (.I(\mult_add_u0.mult0.step6.add_sub4_u0.x4._0_ ),
    .Z(\mult_add_u0.mult0.step6.add_sub4_u0.int_ip[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step7._09_  (.A1(\mult_add_u0.mult0.q0_s6 ),
    .A2(\mult_add_u0.mult0.Q_s6[0] ),
    .Z(\mult_add_u0.mult0.step7._00_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \mult_add_u0.mult0.step7._10_  (.I(\mult_add_u0.mult0.step7._00_ ),
    .Z(\mult_add_u0.mult0.step7._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.mult0.step7._13_  (.I0(\mult_add_u0.mult0.acc_s6[1] ),
    .I1(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.S[1] ),
    .S(\mult_add_u0.mult0.step7._01_ ),
    .Z(\mult_add_u0.mult0.step7._03_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step7._14_  (.I(\mult_add_u0.mult0.step7._03_ ),
    .Z(\mult_add_u0.mult0.step7.next_acc[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.mult0.step7._15_  (.I0(\mult_add_u0.mult0.acc_s6[2] ),
    .I1(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.S[2] ),
    .S(\mult_add_u0.mult0.step7._01_ ),
    .Z(\mult_add_u0.mult0.step7._04_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step7._16_  (.I(\mult_add_u0.mult0.step7._04_ ),
    .Z(\mult_add_u0.mult0.step7.next_acc[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.mult0.step7._17_  (.I0(\mult_add_u0.mult0.acc_s6[3] ),
    .I1(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.S[3] ),
    .S(\mult_add_u0.mult0.step7._01_ ),
    .Z(\mult_add_u0.mult0.step7._05_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step7._18_  (.I(\mult_add_u0.mult0.step7._05_ ),
    .Z(\mult_add_u0.mult0.step7.next_acc[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_add_u0.mult0.step7._23_  (.I0(\mult_add_u0.mult0.acc_s6[0] ),
    .I1(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.S[0] ),
    .S(\mult_add_u0.mult0.step7._01_ ),
    .Z(\mult_add_u0.mult0.step7._08_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step7._24_  (.I(\mult_add_u0.mult0.step7._08_ ),
    .Z(\mult_add_u0.mult0.product[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step7._28_  (.I(\mult_add_u0.mult0.Q_s6[4] ),
    .Z(\mult_add_u0.mult0.product[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step7._29_  (.I(\mult_add_u0.mult0.Q_s6[5] ),
    .Z(\mult_add_u0.mult0.product[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step7._30_  (.I(\mult_add_u0.mult0.Q_s6[6] ),
    .Z(\mult_add_u0.mult0.product[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d1_0.a2._1_  (.A1(\mult_add_u0.mult0.Q_s6[0] ),
    .A2(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d1_0.a2.in0 ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d1_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d1_0.a2._2_  (.I(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d1_0.a2._0_ ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d1_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d1_0.o2._1_  (.A1(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d1_0.g1 ),
    .A2(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d1_0.a2.out ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d1_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d1_0.o2._2_  (.I(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d1_0.o2._0_ ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.cg[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d2_0.a2._1_  (.A1(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.cg[0] ),
    .A2(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d2_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d2_0.a2._2_  (.I(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d2_0.a2._0_ ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d2_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d2_0.o2._1_  (.A1(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d2_0.g1 ),
    .A2(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d2_0.a2.out ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d2_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d2_0.o2._2_  (.I(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d2_0.o2._0_ ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.cg[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d3_0.a1._1_  (.A1(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ),
    .A2(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d3_0.a1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d3_0.a1._2_  (.I(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d3_0.a1._0_ ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.cp21 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d3_0.a2._1_  (.A1(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d2_0.g1 ),
    .A2(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d3_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d3_0.a2._2_  (.I(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d3_0.a2._0_ ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d3_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d3_0.o2._1_  (.A1(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d3_0.g1 ),
    .A2(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d3_0.a2.out ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d3_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d3_0.o2._2_  (.I(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d3_0.o2._0_ ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.cg21 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d3_1.a2._1_  (.A1(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.cg[0] ),
    .A2(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.cp21 ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d3_1.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d3_1.a2._2_  (.I(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d3_1.a2._0_ ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d3_1.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d3_1.o2._1_  (.A1(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.cg21 ),
    .A2(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d3_1.a2.out ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d3_1.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d3_1.o2._2_  (.I(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d3_1.o2._0_ ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.cg[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.p_0.a._1_  (.A1(\mult_add_u0.mult0.step7.add_sub4_u0.int_ip[0] ),
    .A2(\mult_add_u0.mult0.acc_s6[0] ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.p_0.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.p_0.a._2_  (.I(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.p_0.a._0_ ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d1_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.p_0.o._1_  (.A1(\mult_add_u0.mult0.step7.add_sub4_u0.int_ip[0] ),
    .A2(\mult_add_u0.mult0.acc_s6[0] ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.p_0.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.p_0.o._2_  (.I(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.p_0.o._0_ ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d1_0.a2.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.p_1.a._1_  (.A1(\mult_add_u0.mult0.step7.add_sub4_u0.int_ip[1] ),
    .A2(\mult_add_u0.mult0.acc_s6[1] ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.p_1.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.p_1.a._2_  (.I(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.p_1.a._0_ ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d2_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.p_1.o._1_  (.A1(\mult_add_u0.mult0.step7.add_sub4_u0.int_ip[1] ),
    .A2(\mult_add_u0.mult0.acc_s6[1] ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.p_1.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.p_1.o._2_  (.I(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.p_1.o._0_ ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.p_2.a._1_  (.A1(\mult_add_u0.mult0.step7.add_sub4_u0.int_ip[2] ),
    .A2(\mult_add_u0.mult0.acc_s6[2] ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.p_2.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.p_2.a._2_  (.I(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.p_2.a._0_ ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d3_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.p_2.o._1_  (.A1(\mult_add_u0.mult0.step7.add_sub4_u0.int_ip[2] ),
    .A2(\mult_add_u0.mult0.acc_s6[2] ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.p_2.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.p_2.o._2_  (.I(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.p_2.o._0_ ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s0.xor2_0._1_  (.A1(\mult_add_u0.mult0.step7.add_sub4_u0.int_ip[0] ),
    .A2(\mult_add_u0.mult0.acc_s6[0] ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s0.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s0.xor2_0._2_  (.I(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s0.xor2_0._0_ ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s0.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s0.xor2_1._1_  (.A1(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s0.temp ),
    .A2(\mult_add_u0.mult0.Q_s6[0] ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s0.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s0.xor2_1._2_  (.I(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s0.xor2_1._0_ ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.S[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s1.xor2_0._1_  (.A1(\mult_add_u0.mult0.step7.add_sub4_u0.int_ip[1] ),
    .A2(\mult_add_u0.mult0.acc_s6[1] ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s1.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s1.xor2_0._2_  (.I(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s1.xor2_0._0_ ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s1.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s1.xor2_1._1_  (.A1(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s1.temp ),
    .A2(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.cg[0] ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s1.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s1.xor2_1._2_  (.I(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s1.xor2_1._0_ ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.S[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s2.xor2_0._1_  (.A1(\mult_add_u0.mult0.step7.add_sub4_u0.int_ip[2] ),
    .A2(\mult_add_u0.mult0.acc_s6[2] ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s2.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s2.xor2_0._2_  (.I(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s2.xor2_0._0_ ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s2.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s2.xor2_1._1_  (.A1(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s2.temp ),
    .A2(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.cg[1] ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s2.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s2.xor2_1._2_  (.I(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s2.xor2_1._0_ ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.S[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s3.xor2_0._1_  (.A1(\mult_add_u0.mult0.step7.add_sub4_u0.int_ip[3] ),
    .A2(\mult_add_u0.mult0.acc_s6[3] ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s3.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s3.xor2_0._2_  (.I(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s3.xor2_0._0_ ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s3.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s3.xor2_1._1_  (.A1(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s3.temp ),
    .A2(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.cg[2] ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s3.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s3.xor2_1._2_  (.I(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.s3.xor2_1._0_ ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.ppa8_u0.S[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step7.add_sub4_u0.x0._1_  (.A1(\mult_add_u0.mult0.Q_s6[0] ),
    .A2(\mult_add_u0.mult0.multiplicand_s6[0] ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.x0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step7.add_sub4_u0.x0._2_  (.I(\mult_add_u0.mult0.step7.add_sub4_u0.x0._0_ ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.int_ip[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step7.add_sub4_u0.x1._1_  (.A1(\mult_add_u0.mult0.Q_s6[0] ),
    .A2(\mult_add_u0.mult0.multiplicand_s6[1] ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.x1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step7.add_sub4_u0.x1._2_  (.I(\mult_add_u0.mult0.step7.add_sub4_u0.x1._0_ ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.int_ip[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step7.add_sub4_u0.x2._1_  (.A1(\mult_add_u0.mult0.Q_s6[0] ),
    .A2(\mult_add_u0.mult0.multiplicand_s6[2] ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.x2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step7.add_sub4_u0.x2._2_  (.I(\mult_add_u0.mult0.step7.add_sub4_u0.x2._0_ ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.int_ip[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.step7.add_sub4_u0.x3._1_  (.A1(\mult_add_u0.mult0.Q_s6[0] ),
    .A2(\mult_add_u0.mult0.multiplicand_s6[3] ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.x3._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.step7.add_sub4_u0.x3._2_  (.I(\mult_add_u0.mult0.step7.add_sub4_u0.x3._0_ ),
    .Z(\mult_add_u0.mult0.step7.add_sub4_u0.int_ip[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_add_u0.mult0.x_sign._1_  (.A1(\add_u0.a[7] ),
    .A2(\mult_add_u0.m[7] ),
    .Z(\mult_add_u0.mult0.x_sign._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_add_u0.mult0.x_sign._2_  (.I(\mult_add_u0.mult0.x_sign._0_ ),
    .Z(\mult_add_u0.mult0.mul_sign ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \mult_u0._025_  (.I(\mult_u0.product[3] ),
    .ZN(\mult_u0._008_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \mult_u0._026_  (.I(net62),
    .Z(\mult_u0._009_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \mult_u0._027_  (.A1(\mult_u0._008_ ),
    .A2(\mult_u0._009_ ),
    .ZN(\mult_u0._000_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \mult_u0._028_  (.I(\mult_u0.product[4] ),
    .ZN(\mult_u0._010_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \mult_u0._029_  (.A1(\mult_u0._009_ ),
    .A2(\mult_u0._010_ ),
    .ZN(\mult_u0._001_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \mult_u0._030_  (.I(\mult_u0.product[5] ),
    .ZN(\mult_u0._011_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \mult_u0._031_  (.A1(\mult_u0._009_ ),
    .A2(\mult_u0._011_ ),
    .ZN(\mult_u0._002_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \mult_u0._032_  (.I(\mult_u0.product[6] ),
    .ZN(\mult_u0._012_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \mult_u0._033_  (.A1(\mult_u0._009_ ),
    .A2(\mult_u0._012_ ),
    .ZN(\mult_u0._003_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \mult_u0._034_  (.I(\mult_u0.step7.next_acc[0] ),
    .ZN(\mult_u0._013_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \mult_u0._035_  (.A1(\mult_u0._009_ ),
    .A2(\mult_u0._013_ ),
    .ZN(\mult_u0._004_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \mult_u0._036_  (.I(\mult_u0.step7.next_acc[1] ),
    .ZN(\mult_u0._014_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \mult_u0._037_  (.A1(\mult_u0._009_ ),
    .A2(\mult_u0._014_ ),
    .ZN(\mult_u0._005_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \mult_u0._038_  (.I(\mult_u0.step7.next_acc[2] ),
    .ZN(\mult_u0._015_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \mult_u0._039_  (.A1(\mult_u0._009_ ),
    .A2(\mult_u0._015_ ),
    .ZN(\mult_u0._006_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \mult_u0._040_  (.I(\mult_u0.mul_sign_s6 ),
    .ZN(\mult_u0._016_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \mult_u0._041_  (.A1(\mult_u0._009_ ),
    .A2(\mult_u0._016_ ),
    .ZN(\mult_u0._007_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._042_  (.D(\mult_u0._000_ ),
    .CLK(clknet_leaf_10_clk),
    .Q(\mult_u0.product_r[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._043_  (.D(\mult_u0._001_ ),
    .CLK(clknet_leaf_14_clk),
    .Q(\mult_u0.product_r[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._044_  (.D(\mult_u0._002_ ),
    .CLK(clknet_leaf_14_clk),
    .Q(\mult_u0.product_r[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._045_  (.D(\mult_u0._003_ ),
    .CLK(clknet_leaf_13_clk),
    .Q(\mult_u0.product_r[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._046_  (.D(\mult_u0._004_ ),
    .CLK(clknet_leaf_14_clk),
    .Q(\mult_u0.product_r[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._047_  (.D(\mult_u0._005_ ),
    .CLK(clknet_leaf_13_clk),
    .Q(\mult_u0.product_r[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._048_  (.D(\mult_u0._006_ ),
    .CLK(clknet_leaf_13_clk),
    .Q(\mult_u0.product_r[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._049_  (.D(\mult_u0._007_ ),
    .CLK(clknet_leaf_10_clk),
    .Q(\mult_u0.product_r[7] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._050_  (.D(\mult_u0.acc[1][0] ),
    .CLK(clknet_leaf_18_clk),
    .Q(\mult_u0.acc_s1[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._051_  (.D(\mult_u0.acc[1][1] ),
    .CLK(clknet_leaf_18_clk),
    .Q(\mult_u0.acc_s1[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._052_  (.D(\mult_u0.acc[1][2] ),
    .CLK(clknet_leaf_20_clk),
    .Q(\mult_u0.acc_s1[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._053_  (.D(\mult_u0.acc[1][3] ),
    .CLK(clknet_leaf_21_clk),
    .Q(\mult_u0.acc_s1[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._054_  (.D(\mult_u0.acc[1][4] ),
    .CLK(clknet_leaf_23_clk),
    .Q(\mult_u0.acc_s1[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._055_  (.D(\mult_u0.acc[1][5] ),
    .CLK(clknet_leaf_23_clk),
    .Q(\mult_u0.acc_s1[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._056_  (.D(\mult_u0.acc[1][6] ),
    .CLK(clknet_leaf_24_clk),
    .Q(\mult_u0.acc_s1[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 \mult_u0._057_  (.D(\mult_u0.Q[0][0] ),
    .CLK(clknet_leaf_6_clk),
    .Q(\mult_u0.Q_s1[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._058_  (.D(\mult_u0.Q[0][1] ),
    .CLK(clknet_leaf_6_clk),
    .Q(\mult_u0.Q_s1[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._059_  (.D(\mult_u0.Q[0][2] ),
    .CLK(clknet_leaf_90_clk),
    .Q(\mult_u0.Q_s1[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._060_  (.D(\mult_u0.Q[0][3] ),
    .CLK(clknet_leaf_83_clk),
    .Q(\mult_u0.Q_s1[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._061_  (.D(\mult_u0.Q[0][4] ),
    .CLK(clknet_leaf_84_clk),
    .Q(\mult_u0.Q_s1[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._062_  (.D(\mult_u0.Q[0][5] ),
    .CLK(clknet_leaf_89_clk),
    .Q(\mult_u0.Q_s1[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._064_  (.D(\mult_u0.acc[2][0] ),
    .CLK(clknet_leaf_16_clk),
    .Q(\mult_u0.acc_s2[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._065_  (.D(\mult_u0.acc[2][1] ),
    .CLK(clknet_leaf_16_clk),
    .Q(\mult_u0.acc_s2[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._066_  (.D(\mult_u0.acc[2][2] ),
    .CLK(clknet_leaf_21_clk),
    .Q(\mult_u0.acc_s2[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._067_  (.D(\mult_u0.acc[2][3] ),
    .CLK(clknet_leaf_26_clk),
    .Q(\mult_u0.acc_s2[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._068_  (.D(\mult_u0.acc[2][4] ),
    .CLK(clknet_leaf_26_clk),
    .Q(\mult_u0.acc_s2[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._069_  (.D(\mult_u0.acc[2][5] ),
    .CLK(clknet_leaf_25_clk),
    .Q(\mult_u0.acc_s2[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._070_  (.D(\mult_u0.acc[2][6] ),
    .CLK(clknet_leaf_25_clk),
    .Q(\mult_u0.acc_s2[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 \mult_u0._071_  (.D(\mult_u0.Q[1][0] ),
    .CLK(clknet_leaf_17_clk),
    .Q(\mult_u0.Q_s2[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._072_  (.D(\mult_u0.Q[1][1] ),
    .CLK(clknet_leaf_6_clk),
    .Q(\mult_u0.Q_s2[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._073_  (.D(\mult_u0.Q[1][2] ),
    .CLK(clknet_leaf_15_clk),
    .Q(\mult_u0.Q_s2[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._074_  (.D(\mult_u0.Q[1][3] ),
    .CLK(clknet_leaf_84_clk),
    .Q(\mult_u0.Q_s2[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._075_  (.D(\mult_u0.Q[1][4] ),
    .CLK(clknet_leaf_84_clk),
    .Q(\mult_u0.Q_s2[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._078_  (.D(\mult_u0.acc[3][0] ),
    .CLK(clknet_leaf_15_clk),
    .Q(\mult_u0.acc_s3[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._079_  (.D(\mult_u0.acc[3][1] ),
    .CLK(clknet_leaf_31_clk),
    .Q(\mult_u0.acc_s3[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._080_  (.D(\mult_u0.acc[3][2] ),
    .CLK(clknet_leaf_31_clk),
    .Q(\mult_u0.acc_s3[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._081_  (.D(\mult_u0.acc[3][3] ),
    .CLK(clknet_leaf_27_clk),
    .Q(\mult_u0.acc_s3[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._082_  (.D(\mult_u0.acc[3][4] ),
    .CLK(clknet_leaf_27_clk),
    .Q(\mult_u0.acc_s3[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._083_  (.D(\mult_u0.acc[3][5] ),
    .CLK(clknet_leaf_28_clk),
    .Q(\mult_u0.acc_s3[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._084_  (.D(\mult_u0.acc[3][6] ),
    .CLK(clknet_leaf_28_clk),
    .Q(\mult_u0.acc_s3[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 \mult_u0._085_  (.D(\mult_u0.Q[2][0] ),
    .CLK(clknet_leaf_11_clk),
    .Q(\mult_u0.Q_s3[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._086_  (.D(\mult_u0.Q[2][1] ),
    .CLK(clknet_leaf_32_clk),
    .Q(\mult_u0.Q_s3[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._087_  (.D(\mult_u0.Q[2][2] ),
    .CLK(clknet_leaf_34_clk),
    .Q(\mult_u0.Q_s3[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._088_  (.D(\mult_u0.Q[2][3] ),
    .CLK(clknet_leaf_84_clk),
    .Q(\mult_u0.Q_s3[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._092_  (.D(\mult_u0.acc[4][0] ),
    .CLK(clknet_leaf_32_clk),
    .Q(\mult_u0.acc_s4[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._093_  (.D(\mult_u0.acc[4][1] ),
    .CLK(clknet_leaf_30_clk),
    .Q(\mult_u0.acc_s4[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._094_  (.D(\mult_u0.acc[4][2] ),
    .CLK(clknet_leaf_30_clk),
    .Q(\mult_u0.acc_s4[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._095_  (.D(\mult_u0.acc[4][3] ),
    .CLK(clknet_leaf_29_clk),
    .Q(\mult_u0.acc_s4[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._096_  (.D(\mult_u0.acc[4][4] ),
    .CLK(clknet_leaf_29_clk),
    .Q(\mult_u0.acc_s4[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._097_  (.D(\mult_u0.acc[4][5] ),
    .CLK(clknet_leaf_29_clk),
    .Q(\mult_u0.acc_s4[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 \mult_u0._099_  (.D(\mult_u0.Q[3][0] ),
    .CLK(clknet_leaf_32_clk),
    .Q(\mult_u0.Q_s4[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._100_  (.D(\mult_u0.Q[3][1] ),
    .CLK(clknet_leaf_33_clk),
    .Q(\mult_u0.Q_s4[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._101_  (.D(\mult_u0.Q[3][2] ),
    .CLK(clknet_leaf_33_clk),
    .Q(\mult_u0.Q_s4[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._105_  (.D(\mult_u0.Q[3][6] ),
    .CLK(clknet_leaf_17_clk),
    .Q(\mult_u0.Q_s4[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._106_  (.D(\mult_u0.acc[5][0] ),
    .CLK(clknet_leaf_39_clk),
    .Q(\mult_u0.acc_s5[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._107_  (.D(\mult_u0.acc[5][1] ),
    .CLK(clknet_leaf_39_clk),
    .Q(\mult_u0.acc_s5[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._108_  (.D(\mult_u0.acc[5][2] ),
    .CLK(clknet_leaf_40_clk),
    .Q(\mult_u0.acc_s5[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._109_  (.D(\mult_u0.acc[5][3] ),
    .CLK(clknet_leaf_40_clk),
    .Q(\mult_u0.acc_s5[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._110_  (.D(\mult_u0.acc[5][4] ),
    .CLK(clknet_leaf_41_clk),
    .Q(\mult_u0.acc_s5[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 \mult_u0._113_  (.D(\mult_u0.Q[4][0] ),
    .CLK(clknet_leaf_36_clk),
    .Q(\mult_u0.Q_s5[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._114_  (.D(\mult_u0.Q[4][1] ),
    .CLK(clknet_leaf_36_clk),
    .Q(\mult_u0.Q_s5[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._118_  (.D(\mult_u0.Q[4][5] ),
    .CLK(clknet_leaf_17_clk),
    .Q(\mult_u0.Q_s5[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._119_  (.D(\mult_u0.Q[4][6] ),
    .CLK(clknet_leaf_32_clk),
    .Q(\mult_u0.Q_s5[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._120_  (.D(\mult_u0.acc[6][0] ),
    .CLK(clknet_leaf_38_clk),
    .Q(\mult_u0.acc_s6[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._121_  (.D(\mult_u0.acc[6][1] ),
    .CLK(clknet_leaf_38_clk),
    .Q(\mult_u0.acc_s6[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._122_  (.D(\mult_u0.acc[6][2] ),
    .CLK(clknet_leaf_42_clk),
    .Q(\mult_u0.acc_s6[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._123_  (.D(\mult_u0.acc[6][3] ),
    .CLK(clknet_leaf_41_clk),
    .Q(\mult_u0.acc_s6[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 \mult_u0._127_  (.D(\mult_u0.Q[5][0] ),
    .CLK(clknet_leaf_36_clk),
    .Q(\mult_u0.Q_s6[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._131_  (.D(\mult_u0.Q[5][4] ),
    .CLK(clknet_leaf_11_clk),
    .Q(\mult_u0.Q_s6[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._132_  (.D(\mult_u0.Q[5][5] ),
    .CLK(clknet_leaf_34_clk),
    .Q(\mult_u0.Q_s6[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._133_  (.D(\mult_u0.Q[5][6] ),
    .CLK(clknet_leaf_36_clk),
    .Q(\mult_u0.Q_s6[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._134_  (.D(\mult_u0.q0[1] ),
    .CLK(clknet_leaf_21_clk),
    .Q(\mult_u0.q0_s1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._135_  (.D(\mult_u0.q0[2] ),
    .CLK(clknet_leaf_22_clk),
    .Q(\mult_u0.q0_s2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._136_  (.D(\mult_u0.q0[3] ),
    .CLK(clknet_leaf_15_clk),
    .Q(\mult_u0.q0_s3 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._137_  (.D(\mult_u0.q0[4] ),
    .CLK(clknet_leaf_30_clk),
    .Q(\mult_u0.q0_s4 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._138_  (.D(\mult_u0.q0[5] ),
    .CLK(clknet_leaf_40_clk),
    .Q(\mult_u0.q0_s5 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._139_  (.D(\mult_u0.q0[6] ),
    .CLK(clknet_leaf_36_clk),
    .Q(\mult_u0.q0_s6 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._140_  (.D(net121),
    .CLK(clknet_leaf_5_clk),
    .Q(\mult_u0.multiplicand_s1[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._141_  (.D(\mult_u0.multiplicand[1] ),
    .CLK(clknet_leaf_18_clk),
    .Q(\mult_u0.multiplicand_s1[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._142_  (.D(\mult_u0.multiplicand[2] ),
    .CLK(clknet_leaf_20_clk),
    .Q(\mult_u0.multiplicand_s1[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._143_  (.D(\mult_u0.multiplicand[3] ),
    .CLK(clknet_leaf_21_clk),
    .Q(\mult_u0.multiplicand_s1[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._144_  (.D(\mult_u0.multiplicand[4] ),
    .CLK(clknet_leaf_21_clk),
    .Q(\mult_u0.multiplicand_s1[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._145_  (.D(\mult_u0.multiplicand[5] ),
    .CLK(clknet_leaf_22_clk),
    .Q(\mult_u0.multiplicand_s1[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._146_  (.D(\mult_u0.multiplicand[6] ),
    .CLK(clknet_leaf_24_clk),
    .Q(\mult_u0.multiplicand_s1[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._147_  (.D(\mult_u0.multiplicand_s1[0] ),
    .CLK(clknet_leaf_17_clk),
    .Q(\mult_u0.multiplicand_s2[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._148_  (.D(\mult_u0.multiplicand_s1[1] ),
    .CLK(clknet_leaf_16_clk),
    .Q(\mult_u0.multiplicand_s2[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._149_  (.D(\mult_u0.multiplicand_s1[2] ),
    .CLK(clknet_leaf_21_clk),
    .Q(\mult_u0.multiplicand_s2[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._150_  (.D(\mult_u0.multiplicand_s1[3] ),
    .CLK(clknet_leaf_22_clk),
    .Q(\mult_u0.multiplicand_s2[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._151_  (.D(\mult_u0.multiplicand_s1[4] ),
    .CLK(clknet_leaf_26_clk),
    .Q(\mult_u0.multiplicand_s2[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._152_  (.D(\mult_u0.multiplicand_s1[5] ),
    .CLK(clknet_leaf_24_clk),
    .Q(\mult_u0.multiplicand_s2[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._153_  (.D(\mult_u0.multiplicand_s1[6] ),
    .CLK(clknet_leaf_25_clk),
    .Q(\mult_u0.multiplicand_s2[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._154_  (.D(\mult_u0.multiplicand_s2[0] ),
    .CLK(clknet_leaf_16_clk),
    .Q(\mult_u0.multiplicand_s3[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._155_  (.D(\mult_u0.multiplicand_s2[1] ),
    .CLK(clknet_leaf_31_clk),
    .Q(\mult_u0.multiplicand_s3[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._156_  (.D(\mult_u0.multiplicand_s2[2] ),
    .CLK(clknet_leaf_31_clk),
    .Q(\mult_u0.multiplicand_s3[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._157_  (.D(\mult_u0.multiplicand_s2[3] ),
    .CLK(clknet_leaf_27_clk),
    .Q(\mult_u0.multiplicand_s3[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._158_  (.D(\mult_u0.multiplicand_s2[4] ),
    .CLK(clknet_leaf_27_clk),
    .Q(\mult_u0.multiplicand_s3[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._159_  (.D(\mult_u0.multiplicand_s2[5] ),
    .CLK(clknet_leaf_28_clk),
    .Q(\mult_u0.multiplicand_s3[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._160_  (.D(\mult_u0.multiplicand_s2[6] ),
    .CLK(clknet_leaf_25_clk),
    .Q(\mult_u0.multiplicand_s3[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._161_  (.D(\mult_u0.multiplicand_s3[0] ),
    .CLK(clknet_leaf_32_clk),
    .Q(\mult_u0.multiplicand_s4[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._162_  (.D(\mult_u0.multiplicand_s3[1] ),
    .CLK(clknet_leaf_30_clk),
    .Q(\mult_u0.multiplicand_s4[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._163_  (.D(\mult_u0.multiplicand_s3[2] ),
    .CLK(clknet_leaf_30_clk),
    .Q(\mult_u0.multiplicand_s4[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._164_  (.D(\mult_u0.multiplicand_s3[3] ),
    .CLK(clknet_leaf_29_clk),
    .Q(\mult_u0.multiplicand_s4[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._165_  (.D(\mult_u0.multiplicand_s3[4] ),
    .CLK(clknet_leaf_29_clk),
    .Q(\mult_u0.multiplicand_s4[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._166_  (.D(\mult_u0.multiplicand_s3[5] ),
    .CLK(clknet_leaf_29_clk),
    .Q(\mult_u0.multiplicand_s4[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._168_  (.D(\mult_u0.multiplicand_s4[0] ),
    .CLK(clknet_leaf_33_clk),
    .Q(\mult_u0.multiplicand_s5[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._169_  (.D(\mult_u0.multiplicand_s4[1] ),
    .CLK(clknet_leaf_39_clk),
    .Q(\mult_u0.multiplicand_s5[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._170_  (.D(\mult_u0.multiplicand_s4[2] ),
    .CLK(clknet_leaf_39_clk),
    .Q(\mult_u0.multiplicand_s5[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._171_  (.D(\mult_u0.multiplicand_s4[3] ),
    .CLK(clknet_leaf_40_clk),
    .Q(\mult_u0.multiplicand_s5[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._172_  (.D(\mult_u0.multiplicand_s4[4] ),
    .CLK(clknet_leaf_29_clk),
    .Q(\mult_u0.multiplicand_s5[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._175_  (.D(\mult_u0.multiplicand_s5[0] ),
    .CLK(clknet_leaf_36_clk),
    .Q(\mult_u0.multiplicand_s6[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._176_  (.D(\mult_u0.multiplicand_s5[1] ),
    .CLK(clknet_leaf_38_clk),
    .Q(\mult_u0.multiplicand_s6[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._177_  (.D(\mult_u0.multiplicand_s5[2] ),
    .CLK(clknet_leaf_42_clk),
    .Q(\mult_u0.multiplicand_s6[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._178_  (.D(\mult_u0.multiplicand_s5[3] ),
    .CLK(clknet_leaf_41_clk),
    .Q(\mult_u0.multiplicand_s6[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._182_  (.D(\add_u0.b[0] ),
    .CLK(clknet_leaf_6_clk),
    .Q(\mult_u0.multiplicand[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._183_  (.D(\add_u0.b[1] ),
    .CLK(clknet_leaf_5_clk),
    .Q(\mult_u0.multiplicand[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._184_  (.D(\add_u0.b[2] ),
    .CLK(clknet_leaf_18_clk),
    .Q(\mult_u0.multiplicand[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._185_  (.D(\add_u0.b[3] ),
    .CLK(clknet_leaf_5_clk),
    .Q(\mult_u0.multiplicand[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._186_  (.D(\add_u0.b[4] ),
    .CLK(clknet_leaf_21_clk),
    .Q(\mult_u0.multiplicand[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._187_  (.D(\add_u0.b[5] ),
    .CLK(clknet_leaf_21_clk),
    .Q(\mult_u0.multiplicand[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._188_  (.D(\add_u0.b[6] ),
    .CLK(clknet_leaf_21_clk),
    .Q(\mult_u0.multiplicand[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 \mult_u0._189_  (.D(\add_u0.a[0] ),
    .CLK(clknet_leaf_0_clk),
    .Q(\mult_u0.multiplier[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._190_  (.D(\add_u0.a[1] ),
    .CLK(clknet_leaf_1_clk),
    .Q(\mult_u0.multiplier[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._191_  (.D(\add_u0.a[2] ),
    .CLK(clknet_leaf_5_clk),
    .Q(\mult_u0.multiplier[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._192_  (.D(\add_u0.a[3] ),
    .CLK(clknet_leaf_91_clk),
    .Q(\mult_u0.multiplier[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._193_  (.D(\add_u0.a[4] ),
    .CLK(clknet_leaf_90_clk),
    .Q(\mult_u0.multiplier[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._194_  (.D(\add_u0.a[5] ),
    .CLK(clknet_leaf_89_clk),
    .Q(\mult_u0.multiplier[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._195_  (.D(\add_u0.a[6] ),
    .CLK(clknet_leaf_89_clk),
    .Q(\mult_u0.multiplier[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._196_  (.D(\mult_u0.mul_sign ),
    .CLK(clknet_leaf_92_clk),
    .Q(\mult_u0.mul_sign_s1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._197_  (.D(\mult_u0.mul_sign_s1 ),
    .CLK(clknet_leaf_92_clk),
    .Q(\mult_u0.mul_sign_s2 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._198_  (.D(\mult_u0.mul_sign_s2 ),
    .CLK(clknet_leaf_92_clk),
    .Q(\mult_u0.mul_sign_s3 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._199_  (.D(\mult_u0.mul_sign_s3 ),
    .CLK(clknet_leaf_88_clk),
    .Q(\mult_u0.mul_sign_s4 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._200_  (.D(net147),
    .CLK(clknet_leaf_89_clk),
    .Q(\mult_u0.mul_sign_s5 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 \mult_u0._201_  (.D(\mult_u0.mul_sign_s5 ),
    .CLK(clknet_leaf_89_clk),
    .Q(\mult_u0.mul_sign_s6 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step1._09_  (.A1(net113),
    .A2(\mult_u0.multiplier[0] ),
    .Z(\mult_u0.step1._00_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_u0.step1._09__113  (.ZN(net113),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 \mult_u0.step1._10_  (.I(\mult_u0.step1._00_ ),
    .Z(\mult_u0.step1._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_u0.step1._11_  (.I0(net111),
    .I1(\mult_u0.step1.add_sub4_u0.ppa8_u0.S[6] ),
    .S(\mult_u0.step1._01_ ),
    .Z(\mult_u0.step1._02_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_u0.step1._11__111  (.ZN(net111),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1._12_  (.I(\mult_u0.step1._02_ ),
    .Z(\mult_u0.acc[1][6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_u0.step1._13_  (.I0(net91),
    .I1(\mult_u0.step1.add_sub4_u0.ppa8_u0.S[1] ),
    .S(\mult_u0.step1._01_ ),
    .Z(\mult_u0.step1._03_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_u0.step1._13__91  (.ZN(net91),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1._14_  (.I(\mult_u0.step1._03_ ),
    .Z(\mult_u0.acc[1][0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_u0.step1._15_  (.I0(net95),
    .I1(\mult_u0.step1.add_sub4_u0.ppa8_u0.S[2] ),
    .S(\mult_u0.step1._01_ ),
    .Z(\mult_u0.step1._04_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_u0.step1._15__95  (.ZN(net95),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1._16_  (.I(\mult_u0.step1._04_ ),
    .Z(\mult_u0.acc[1][1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_u0.step1._17_  (.I0(net99),
    .I1(\mult_u0.step1.add_sub4_u0.ppa8_u0.S[3] ),
    .S(\mult_u0.step1._01_ ),
    .Z(\mult_u0.step1._05_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_u0.step1._17__99  (.ZN(net99),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1._18_  (.I(\mult_u0.step1._05_ ),
    .Z(\mult_u0.acc[1][2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_u0.step1._19_  (.I0(net103),
    .I1(\mult_u0.step1.add_sub4_u0.ppa8_u0.S[4] ),
    .S(\mult_u0.step1._01_ ),
    .Z(\mult_u0.step1._06_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_u0.step1._19__103  (.ZN(net103),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1._20_  (.I(\mult_u0.step1._06_ ),
    .Z(\mult_u0.acc[1][3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_u0.step1._21_  (.I0(net107),
    .I1(\mult_u0.step1.add_sub4_u0.ppa8_u0.S[5] ),
    .S(\mult_u0.step1._01_ ),
    .Z(\mult_u0.step1._07_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_u0.step1._21__107  (.ZN(net107),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1._22_  (.I(\mult_u0.step1._07_ ),
    .Z(\mult_u0.acc[1][4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1._25_  (.I(\mult_u0.multiplier[1] ),
    .Z(\mult_u0.Q[0][0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1._26_  (.I(\mult_u0.multiplier[2] ),
    .Z(\mult_u0.Q[0][1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1._27_  (.I(\mult_u0.multiplier[3] ),
    .Z(\mult_u0.Q[0][2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1._28_  (.I(\mult_u0.multiplier[4] ),
    .Z(\mult_u0.Q[0][3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1._29_  (.I(\mult_u0.multiplier[5] ),
    .Z(\mult_u0.Q[0][4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1._30_  (.I(\mult_u0.multiplier[6] ),
    .Z(\mult_u0.Q[0][5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1._31_  (.I(\mult_u0.acc[1][6] ),
    .Z(\mult_u0.acc[1][5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1._32_  (.I(\mult_u0.multiplier[0] ),
    .Z(\mult_u0.q0[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.d1_0.a2._1_  (.A1(\mult_u0.multiplier[0] ),
    .A2(\mult_u0.step1.add_sub4_u0.ppa8_u0.d1_0.a2.in0 ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.d1_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.d1_0.a2._2_  (.I(\mult_u0.step1.add_sub4_u0.ppa8_u0.d1_0.a2._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.d1_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.d1_0.o2._1_  (.A1(\mult_u0.step1.add_sub4_u0.ppa8_u0.d1_0.g1 ),
    .A2(\mult_u0.step1.add_sub4_u0.ppa8_u0.d1_0.a2.out ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.d1_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.d1_0.o2._2_  (.I(\mult_u0.step1.add_sub4_u0.ppa8_u0.d1_0.o2._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.cg[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.d2_0.a2._1_  (.A1(\mult_u0.step1.add_sub4_u0.ppa8_u0.cg[0] ),
    .A2(\mult_u0.step1.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.d2_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.d2_0.a2._2_  (.I(\mult_u0.step1.add_sub4_u0.ppa8_u0.d2_0.a2._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.d2_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.d2_0.o2._1_  (.A1(\mult_u0.step1.add_sub4_u0.ppa8_u0.d2_0.g1 ),
    .A2(\mult_u0.step1.add_sub4_u0.ppa8_u0.d2_0.a2.out ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.d2_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.d2_0.o2._2_  (.I(\mult_u0.step1.add_sub4_u0.ppa8_u0.d2_0.o2._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.cg[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.d3_0.a1._1_  (.A1(\mult_u0.step1.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ),
    .A2(\mult_u0.step1.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.d3_0.a1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.d3_0.a1._2_  (.I(\mult_u0.step1.add_sub4_u0.ppa8_u0.d3_0.a1._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.cp21 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.d3_0.a2._1_  (.A1(\mult_u0.step1.add_sub4_u0.ppa8_u0.d2_0.g1 ),
    .A2(\mult_u0.step1.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.d3_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.d3_0.a2._2_  (.I(\mult_u0.step1.add_sub4_u0.ppa8_u0.d3_0.a2._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.d3_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.d3_0.o2._1_  (.A1(\mult_u0.step1.add_sub4_u0.ppa8_u0.d3_0.g1 ),
    .A2(\mult_u0.step1.add_sub4_u0.ppa8_u0.d3_0.a2.out ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.d3_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.d3_0.o2._2_  (.I(\mult_u0.step1.add_sub4_u0.ppa8_u0.d3_0.o2._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.cg21 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.d3_1.a2._1_  (.A1(\mult_u0.step1.add_sub4_u0.ppa8_u0.cg[0] ),
    .A2(\mult_u0.step1.add_sub4_u0.ppa8_u0.cp21 ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.d3_1.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.d3_1.a2._2_  (.I(\mult_u0.step1.add_sub4_u0.ppa8_u0.d3_1.a2._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.d3_1.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.d3_1.o2._1_  (.A1(\mult_u0.step1.add_sub4_u0.ppa8_u0.cg21 ),
    .A2(\mult_u0.step1.add_sub4_u0.ppa8_u0.d3_1.a2.out ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.d3_1.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.d3_1.o2._2_  (.I(\mult_u0.step1.add_sub4_u0.ppa8_u0.d3_1.o2._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.cg[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.d4_0.a2._1_  (.A1(\mult_u0.step1.add_sub4_u0.ppa8_u0.cg[2] ),
    .A2(\mult_u0.step1.add_sub4_u0.ppa8_u0.d4_0.a2.in0 ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.d4_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.d4_0.a2._2_  (.I(\mult_u0.step1.add_sub4_u0.ppa8_u0.d4_0.a2._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.d4_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.d4_0.o2._1_  (.A1(\mult_u0.step1.add_sub4_u0.ppa8_u0.d4_0.g1 ),
    .A2(\mult_u0.step1.add_sub4_u0.ppa8_u0.d4_0.a2.out ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.d4_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.d4_0.o2._2_  (.I(\mult_u0.step1.add_sub4_u0.ppa8_u0.d4_0.o2._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.cg[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.d5_0.a1._1_  (.A1(\mult_u0.step1.add_sub4_u0.ppa8_u0.d4_0.a2.in0 ),
    .A2(\mult_u0.step1.add_sub4_u0.ppa8_u0.d5_0.a1.in0 ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.d5_0.a1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.d5_0.a1._2_  (.I(\mult_u0.step1.add_sub4_u0.ppa8_u0.d5_0.a1._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.cp43 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.d5_0.a2._1_  (.A1(\mult_u0.step1.add_sub4_u0.ppa8_u0.d4_0.g1 ),
    .A2(\mult_u0.step1.add_sub4_u0.ppa8_u0.d5_0.a1.in0 ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.d5_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.d5_0.a2._2_  (.I(\mult_u0.step1.add_sub4_u0.ppa8_u0.d5_0.a2._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.d5_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.d5_0.o2._1_  (.A1(\mult_u0.step1.add_sub4_u0.ppa8_u0.d5_0.g1 ),
    .A2(\mult_u0.step1.add_sub4_u0.ppa8_u0.d5_0.a2.out ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.d5_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.d5_0.o2._2_  (.I(\mult_u0.step1.add_sub4_u0.ppa8_u0.d5_0.o2._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.cg43 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.d5_1.a2._1_  (.A1(\mult_u0.step1.add_sub4_u0.ppa8_u0.cg[2] ),
    .A2(\mult_u0.step1.add_sub4_u0.ppa8_u0.cp43 ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.d5_1.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.d5_1.a2._2_  (.I(\mult_u0.step1.add_sub4_u0.ppa8_u0.d5_1.a2._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.d5_1.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.d5_1.o2._1_  (.A1(\mult_u0.step1.add_sub4_u0.ppa8_u0.cg43 ),
    .A2(\mult_u0.step1.add_sub4_u0.ppa8_u0.d5_1.a2.out ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.d5_1.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.d5_1.o2._2_  (.I(\mult_u0.step1.add_sub4_u0.ppa8_u0.d5_1.o2._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.cg[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.d6_0.a1._1_  (.A1(\mult_u0.step1.add_sub4_u0.ppa8_u0.cp43 ),
    .A2(\mult_u0.step1.add_sub4_u0.ppa8_u0.d6_0.a1.in0 ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.d6_0.a1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.d6_0.a1._2_  (.I(\mult_u0.step1.add_sub4_u0.ppa8_u0.d6_0.a1._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.cp54 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.d6_0.a2._1_  (.A1(\mult_u0.step1.add_sub4_u0.ppa8_u0.cg43 ),
    .A2(\mult_u0.step1.add_sub4_u0.ppa8_u0.d6_0.a1.in0 ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.d6_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.d6_0.a2._2_  (.I(\mult_u0.step1.add_sub4_u0.ppa8_u0.d6_0.a2._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.d6_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.d6_0.o2._1_  (.A1(\mult_u0.step1.add_sub4_u0.ppa8_u0.d6_0.g1 ),
    .A2(\mult_u0.step1.add_sub4_u0.ppa8_u0.d6_0.a2.out ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.d6_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.d6_0.o2._2_  (.I(\mult_u0.step1.add_sub4_u0.ppa8_u0.d6_0.o2._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.cg54 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.d6_1.a2._1_  (.A1(\mult_u0.step1.add_sub4_u0.ppa8_u0.cg[2] ),
    .A2(\mult_u0.step1.add_sub4_u0.ppa8_u0.cp54 ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.d6_1.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.d6_1.a2._2_  (.I(\mult_u0.step1.add_sub4_u0.ppa8_u0.d6_1.a2._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.d6_1.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.d6_1.o2._1_  (.A1(\mult_u0.step1.add_sub4_u0.ppa8_u0.cg54 ),
    .A2(\mult_u0.step1.add_sub4_u0.ppa8_u0.d6_1.a2.out ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.d6_1.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.d6_1.o2._2_  (.I(\mult_u0.step1.add_sub4_u0.ppa8_u0.d6_1.o2._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.cg[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.p_0.a._1_  (.A1(\mult_u0.step1.add_sub4_u0.int_ip[0] ),
    .A2(net89),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.p_0.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_u0.step1.add_sub4_u0.ppa8_u0.p_0.a._1__89  (.ZN(net89),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.p_0.a._2_  (.I(\mult_u0.step1.add_sub4_u0.ppa8_u0.p_0.a._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.d1_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.p_0.o._1_  (.A1(\mult_u0.step1.add_sub4_u0.int_ip[0] ),
    .A2(net90),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.p_0.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_u0.step1.add_sub4_u0.ppa8_u0.p_0.o._1__90  (.ZN(net90),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.p_0.o._2_  (.I(\mult_u0.step1.add_sub4_u0.ppa8_u0.p_0.o._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.d1_0.a2.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.p_1.a._1_  (.A1(\mult_u0.step1.add_sub4_u0.int_ip[1] ),
    .A2(net92),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.p_1.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_u0.step1.add_sub4_u0.ppa8_u0.p_1.a._1__92  (.ZN(net92),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.p_1.a._2_  (.I(\mult_u0.step1.add_sub4_u0.ppa8_u0.p_1.a._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.d2_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.p_1.o._1_  (.A1(\mult_u0.step1.add_sub4_u0.int_ip[1] ),
    .A2(net93),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.p_1.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_u0.step1.add_sub4_u0.ppa8_u0.p_1.o._1__93  (.ZN(net93),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.p_1.o._2_  (.I(\mult_u0.step1.add_sub4_u0.ppa8_u0.p_1.o._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.p_2.a._1_  (.A1(\mult_u0.step1.add_sub4_u0.int_ip[2] ),
    .A2(net96),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.p_2.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_u0.step1.add_sub4_u0.ppa8_u0.p_2.a._1__96  (.ZN(net96),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.p_2.a._2_  (.I(\mult_u0.step1.add_sub4_u0.ppa8_u0.p_2.a._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.d3_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.p_2.o._1_  (.A1(\mult_u0.step1.add_sub4_u0.int_ip[2] ),
    .A2(net97),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.p_2.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_u0.step1.add_sub4_u0.ppa8_u0.p_2.o._1__97  (.ZN(net97),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.p_2.o._2_  (.I(\mult_u0.step1.add_sub4_u0.ppa8_u0.p_2.o._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.p_3.a._1_  (.A1(\mult_u0.step1.add_sub4_u0.int_ip[3] ),
    .A2(net100),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.p_3.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_u0.step1.add_sub4_u0.ppa8_u0.p_3.a._1__100  (.ZN(net100),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.p_3.a._2_  (.I(\mult_u0.step1.add_sub4_u0.ppa8_u0.p_3.a._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.d4_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.p_3.o._1_  (.A1(\mult_u0.step1.add_sub4_u0.int_ip[3] ),
    .A2(net101),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.p_3.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_u0.step1.add_sub4_u0.ppa8_u0.p_3.o._1__101  (.ZN(net101),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.p_3.o._2_  (.I(\mult_u0.step1.add_sub4_u0.ppa8_u0.p_3.o._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.d4_0.a2.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.p_4.a._1_  (.A1(\mult_u0.step1.add_sub4_u0.int_ip[4] ),
    .A2(net104),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.p_4.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_u0.step1.add_sub4_u0.ppa8_u0.p_4.a._1__104  (.ZN(net104),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.p_4.a._2_  (.I(\mult_u0.step1.add_sub4_u0.ppa8_u0.p_4.a._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.d5_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.p_4.o._1_  (.A1(\mult_u0.step1.add_sub4_u0.int_ip[4] ),
    .A2(net105),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.p_4.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_u0.step1.add_sub4_u0.ppa8_u0.p_4.o._1__105  (.ZN(net105),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.p_4.o._2_  (.I(\mult_u0.step1.add_sub4_u0.ppa8_u0.p_4.o._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.d5_0.a1.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.p_5.a._1_  (.A1(\mult_u0.step1.add_sub4_u0.int_ip[5] ),
    .A2(net108),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.p_5.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_u0.step1.add_sub4_u0.ppa8_u0.p_5.a._1__108  (.ZN(net108),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.p_5.a._2_  (.I(\mult_u0.step1.add_sub4_u0.ppa8_u0.p_5.a._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.d6_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.p_5.o._1_  (.A1(\mult_u0.step1.add_sub4_u0.int_ip[5] ),
    .A2(net109),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.p_5.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_u0.step1.add_sub4_u0.ppa8_u0.p_5.o._1__109  (.ZN(net109),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.p_5.o._2_  (.I(\mult_u0.step1.add_sub4_u0.ppa8_u0.p_5.o._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.d6_0.a1.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.s1.xor2_0._1_  (.A1(\mult_u0.step1.add_sub4_u0.int_ip[1] ),
    .A2(net94),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.s1.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_u0.step1.add_sub4_u0.ppa8_u0.s1.xor2_0._1__94  (.ZN(net94),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.s1.xor2_0._2_  (.I(\mult_u0.step1.add_sub4_u0.ppa8_u0.s1.xor2_0._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.s1.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.s1.xor2_1._1_  (.A1(\mult_u0.step1.add_sub4_u0.ppa8_u0.s1.temp ),
    .A2(\mult_u0.step1.add_sub4_u0.ppa8_u0.cg[0] ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.s1.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.s1.xor2_1._2_  (.I(\mult_u0.step1.add_sub4_u0.ppa8_u0.s1.xor2_1._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.S[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.s2.xor2_0._1_  (.A1(\mult_u0.step1.add_sub4_u0.int_ip[2] ),
    .A2(net98),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.s2.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_u0.step1.add_sub4_u0.ppa8_u0.s2.xor2_0._1__98  (.ZN(net98),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.s2.xor2_0._2_  (.I(\mult_u0.step1.add_sub4_u0.ppa8_u0.s2.xor2_0._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.s2.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.s2.xor2_1._1_  (.A1(\mult_u0.step1.add_sub4_u0.ppa8_u0.s2.temp ),
    .A2(\mult_u0.step1.add_sub4_u0.ppa8_u0.cg[1] ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.s2.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.s2.xor2_1._2_  (.I(\mult_u0.step1.add_sub4_u0.ppa8_u0.s2.xor2_1._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.S[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.s3.xor2_0._1_  (.A1(\mult_u0.step1.add_sub4_u0.int_ip[3] ),
    .A2(net102),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.s3.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_u0.step1.add_sub4_u0.ppa8_u0.s3.xor2_0._1__102  (.ZN(net102),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.s3.xor2_0._2_  (.I(\mult_u0.step1.add_sub4_u0.ppa8_u0.s3.xor2_0._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.s3.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.s3.xor2_1._1_  (.A1(\mult_u0.step1.add_sub4_u0.ppa8_u0.s3.temp ),
    .A2(\mult_u0.step1.add_sub4_u0.ppa8_u0.cg[2] ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.s3.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.s3.xor2_1._2_  (.I(\mult_u0.step1.add_sub4_u0.ppa8_u0.s3.xor2_1._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.S[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.s4.xor2_0._1_  (.A1(\mult_u0.step1.add_sub4_u0.int_ip[4] ),
    .A2(net106),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.s4.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_u0.step1.add_sub4_u0.ppa8_u0.s4.xor2_0._1__106  (.ZN(net106),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.s4.xor2_0._2_  (.I(\mult_u0.step1.add_sub4_u0.ppa8_u0.s4.xor2_0._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.s4.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.s4.xor2_1._1_  (.A1(\mult_u0.step1.add_sub4_u0.ppa8_u0.s4.temp ),
    .A2(\mult_u0.step1.add_sub4_u0.ppa8_u0.cg[3] ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.s4.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.s4.xor2_1._2_  (.I(\mult_u0.step1.add_sub4_u0.ppa8_u0.s4.xor2_1._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.S[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.s5.xor2_0._1_  (.A1(\mult_u0.step1.add_sub4_u0.int_ip[5] ),
    .A2(net110),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.s5.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_u0.step1.add_sub4_u0.ppa8_u0.s5.xor2_0._1__110  (.ZN(net110),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.s5.xor2_0._2_  (.I(\mult_u0.step1.add_sub4_u0.ppa8_u0.s5.xor2_0._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.s5.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.s5.xor2_1._1_  (.A1(\mult_u0.step1.add_sub4_u0.ppa8_u0.s5.temp ),
    .A2(\mult_u0.step1.add_sub4_u0.ppa8_u0.cg[4] ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.s5.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.s5.xor2_1._2_  (.I(\mult_u0.step1.add_sub4_u0.ppa8_u0.s5.xor2_1._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.S[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.s6.xor2_0._1_  (.A1(\mult_u0.step1.add_sub4_u0.int_ip[6] ),
    .A2(net112),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.s6.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \mult_u0.step1.add_sub4_u0.ppa8_u0.s6.xor2_0._1__112  (.ZN(net112),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.s6.xor2_0._2_  (.I(\mult_u0.step1.add_sub4_u0.ppa8_u0.s6.xor2_0._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.s6.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.s6.xor2_1._1_  (.A1(\mult_u0.step1.add_sub4_u0.ppa8_u0.s6.temp ),
    .A2(\mult_u0.step1.add_sub4_u0.ppa8_u0.cg[5] ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.s6.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1.add_sub4_u0.ppa8_u0.s6.xor2_1._2_  (.I(\mult_u0.step1.add_sub4_u0.ppa8_u0.s6.xor2_1._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.ppa8_u0.S[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step1.add_sub4_u0.x0._1_  (.A1(\mult_u0.multiplier[0] ),
    .A2(\mult_u0.multiplicand[0] ),
    .Z(\mult_u0.step1.add_sub4_u0.x0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1.add_sub4_u0.x0._2_  (.I(\mult_u0.step1.add_sub4_u0.x0._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.int_ip[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step1.add_sub4_u0.x1._1_  (.A1(\mult_u0.multiplier[0] ),
    .A2(\mult_u0.multiplicand[1] ),
    .Z(\mult_u0.step1.add_sub4_u0.x1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1.add_sub4_u0.x1._2_  (.I(\mult_u0.step1.add_sub4_u0.x1._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.int_ip[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step1.add_sub4_u0.x2._1_  (.A1(\mult_u0.multiplier[0] ),
    .A2(\mult_u0.multiplicand[2] ),
    .Z(\mult_u0.step1.add_sub4_u0.x2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1.add_sub4_u0.x2._2_  (.I(\mult_u0.step1.add_sub4_u0.x2._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.int_ip[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step1.add_sub4_u0.x3._1_  (.A1(\mult_u0.multiplier[0] ),
    .A2(\mult_u0.multiplicand[3] ),
    .Z(\mult_u0.step1.add_sub4_u0.x3._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1.add_sub4_u0.x3._2_  (.I(\mult_u0.step1.add_sub4_u0.x3._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.int_ip[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step1.add_sub4_u0.x4._1_  (.A1(\mult_u0.multiplier[0] ),
    .A2(\mult_u0.multiplicand[4] ),
    .Z(\mult_u0.step1.add_sub4_u0.x4._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1.add_sub4_u0.x4._2_  (.I(\mult_u0.step1.add_sub4_u0.x4._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.int_ip[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step1.add_sub4_u0.x5._1_  (.A1(\mult_u0.multiplier[0] ),
    .A2(\mult_u0.multiplicand[5] ),
    .Z(\mult_u0.step1.add_sub4_u0.x5._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1.add_sub4_u0.x5._2_  (.I(\mult_u0.step1.add_sub4_u0.x5._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.int_ip[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step1.add_sub4_u0.x6._1_  (.A1(\mult_u0.multiplier[0] ),
    .A2(\mult_u0.multiplicand[6] ),
    .Z(\mult_u0.step1.add_sub4_u0.x6._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step1.add_sub4_u0.x6._2_  (.I(\mult_u0.step1.add_sub4_u0.x6._0_ ),
    .Z(\mult_u0.step1.add_sub4_u0.int_ip[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step2._09_  (.A1(\mult_u0.q0_s1 ),
    .A2(\mult_u0.Q_s1[0] ),
    .Z(\mult_u0.step2._00_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 \mult_u0.step2._10_  (.I(\mult_u0.step2._00_ ),
    .Z(\mult_u0.step2._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_u0.step2._11_  (.I0(\mult_u0.acc_s1[6] ),
    .I1(\mult_u0.step2.add_sub4_u0.ppa8_u0.S[6] ),
    .S(\mult_u0.step2._01_ ),
    .Z(\mult_u0.step2._02_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2._12_  (.I(\mult_u0.step2._02_ ),
    .Z(\mult_u0.acc[2][6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_u0.step2._13_  (.I0(\mult_u0.acc_s1[1] ),
    .I1(\mult_u0.step2.add_sub4_u0.ppa8_u0.S[1] ),
    .S(\mult_u0.step2._01_ ),
    .Z(\mult_u0.step2._03_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2._14_  (.I(\mult_u0.step2._03_ ),
    .Z(\mult_u0.acc[2][0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_u0.step2._15_  (.I0(\mult_u0.acc_s1[2] ),
    .I1(\mult_u0.step2.add_sub4_u0.ppa8_u0.S[2] ),
    .S(\mult_u0.step2._01_ ),
    .Z(\mult_u0.step2._04_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2._16_  (.I(\mult_u0.step2._04_ ),
    .Z(\mult_u0.acc[2][1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_u0.step2._17_  (.I0(\mult_u0.acc_s1[3] ),
    .I1(\mult_u0.step2.add_sub4_u0.ppa8_u0.S[3] ),
    .S(\mult_u0.step2._01_ ),
    .Z(\mult_u0.step2._05_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2._18_  (.I(\mult_u0.step2._05_ ),
    .Z(\mult_u0.acc[2][2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_u0.step2._19_  (.I0(\mult_u0.acc_s1[4] ),
    .I1(\mult_u0.step2.add_sub4_u0.ppa8_u0.S[4] ),
    .S(\mult_u0.step2._01_ ),
    .Z(\mult_u0.step2._06_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2._20_  (.I(\mult_u0.step2._06_ ),
    .Z(\mult_u0.acc[2][3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_u0.step2._21_  (.I0(\mult_u0.acc_s1[5] ),
    .I1(\mult_u0.step2.add_sub4_u0.ppa8_u0.S[5] ),
    .S(\mult_u0.step2._01_ ),
    .Z(\mult_u0.step2._07_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2._22_  (.I(\mult_u0.step2._07_ ),
    .Z(\mult_u0.acc[2][4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2._25_  (.I(\mult_u0.Q_s1[1] ),
    .Z(\mult_u0.Q[1][0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2._26_  (.I(\mult_u0.Q_s1[2] ),
    .Z(\mult_u0.Q[1][1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2._27_  (.I(\mult_u0.Q_s1[3] ),
    .Z(\mult_u0.Q[1][2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2._28_  (.I(\mult_u0.Q_s1[4] ),
    .Z(\mult_u0.Q[1][3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2._29_  (.I(\mult_u0.Q_s1[5] ),
    .Z(\mult_u0.Q[1][4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2._31_  (.I(\mult_u0.acc[2][6] ),
    .Z(\mult_u0.acc[2][5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2._32_  (.I(\mult_u0.Q_s1[0] ),
    .Z(\mult_u0.q0[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.d1_0.a2._1_  (.A1(\mult_u0.Q_s1[0] ),
    .A2(\mult_u0.step2.add_sub4_u0.ppa8_u0.d1_0.a2.in0 ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.d1_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.d1_0.a2._2_  (.I(\mult_u0.step2.add_sub4_u0.ppa8_u0.d1_0.a2._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.d1_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.d1_0.o2._1_  (.A1(\mult_u0.step2.add_sub4_u0.ppa8_u0.d1_0.g1 ),
    .A2(\mult_u0.step2.add_sub4_u0.ppa8_u0.d1_0.a2.out ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.d1_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.d1_0.o2._2_  (.I(\mult_u0.step2.add_sub4_u0.ppa8_u0.d1_0.o2._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.cg[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.d2_0.a2._1_  (.A1(\mult_u0.step2.add_sub4_u0.ppa8_u0.cg[0] ),
    .A2(\mult_u0.step2.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.d2_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.d2_0.a2._2_  (.I(\mult_u0.step2.add_sub4_u0.ppa8_u0.d2_0.a2._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.d2_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.d2_0.o2._1_  (.A1(\mult_u0.step2.add_sub4_u0.ppa8_u0.d2_0.g1 ),
    .A2(\mult_u0.step2.add_sub4_u0.ppa8_u0.d2_0.a2.out ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.d2_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.d2_0.o2._2_  (.I(\mult_u0.step2.add_sub4_u0.ppa8_u0.d2_0.o2._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.cg[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.d3_0.a1._1_  (.A1(\mult_u0.step2.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ),
    .A2(\mult_u0.step2.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.d3_0.a1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.d3_0.a1._2_  (.I(\mult_u0.step2.add_sub4_u0.ppa8_u0.d3_0.a1._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.cp21 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.d3_0.a2._1_  (.A1(\mult_u0.step2.add_sub4_u0.ppa8_u0.d2_0.g1 ),
    .A2(\mult_u0.step2.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.d3_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.d3_0.a2._2_  (.I(\mult_u0.step2.add_sub4_u0.ppa8_u0.d3_0.a2._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.d3_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.d3_0.o2._1_  (.A1(\mult_u0.step2.add_sub4_u0.ppa8_u0.d3_0.g1 ),
    .A2(\mult_u0.step2.add_sub4_u0.ppa8_u0.d3_0.a2.out ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.d3_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.d3_0.o2._2_  (.I(\mult_u0.step2.add_sub4_u0.ppa8_u0.d3_0.o2._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.cg21 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.d3_1.a2._1_  (.A1(\mult_u0.step2.add_sub4_u0.ppa8_u0.cg[0] ),
    .A2(\mult_u0.step2.add_sub4_u0.ppa8_u0.cp21 ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.d3_1.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.d3_1.a2._2_  (.I(\mult_u0.step2.add_sub4_u0.ppa8_u0.d3_1.a2._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.d3_1.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.d3_1.o2._1_  (.A1(\mult_u0.step2.add_sub4_u0.ppa8_u0.cg21 ),
    .A2(\mult_u0.step2.add_sub4_u0.ppa8_u0.d3_1.a2.out ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.d3_1.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.d3_1.o2._2_  (.I(\mult_u0.step2.add_sub4_u0.ppa8_u0.d3_1.o2._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.cg[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.d4_0.a2._1_  (.A1(\mult_u0.step2.add_sub4_u0.ppa8_u0.cg[2] ),
    .A2(\mult_u0.step2.add_sub4_u0.ppa8_u0.d4_0.a2.in0 ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.d4_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.d4_0.a2._2_  (.I(\mult_u0.step2.add_sub4_u0.ppa8_u0.d4_0.a2._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.d4_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.d4_0.o2._1_  (.A1(\mult_u0.step2.add_sub4_u0.ppa8_u0.d4_0.g1 ),
    .A2(\mult_u0.step2.add_sub4_u0.ppa8_u0.d4_0.a2.out ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.d4_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.d4_0.o2._2_  (.I(\mult_u0.step2.add_sub4_u0.ppa8_u0.d4_0.o2._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.cg[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.d5_0.a1._1_  (.A1(\mult_u0.step2.add_sub4_u0.ppa8_u0.d4_0.a2.in0 ),
    .A2(\mult_u0.step2.add_sub4_u0.ppa8_u0.d5_0.a1.in0 ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.d5_0.a1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.d5_0.a1._2_  (.I(\mult_u0.step2.add_sub4_u0.ppa8_u0.d5_0.a1._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.cp43 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.d5_0.a2._1_  (.A1(\mult_u0.step2.add_sub4_u0.ppa8_u0.d4_0.g1 ),
    .A2(\mult_u0.step2.add_sub4_u0.ppa8_u0.d5_0.a1.in0 ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.d5_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.d5_0.a2._2_  (.I(\mult_u0.step2.add_sub4_u0.ppa8_u0.d5_0.a2._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.d5_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.d5_0.o2._1_  (.A1(\mult_u0.step2.add_sub4_u0.ppa8_u0.d5_0.g1 ),
    .A2(\mult_u0.step2.add_sub4_u0.ppa8_u0.d5_0.a2.out ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.d5_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.d5_0.o2._2_  (.I(\mult_u0.step2.add_sub4_u0.ppa8_u0.d5_0.o2._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.cg43 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.d5_1.a2._1_  (.A1(\mult_u0.step2.add_sub4_u0.ppa8_u0.cg[2] ),
    .A2(\mult_u0.step2.add_sub4_u0.ppa8_u0.cp43 ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.d5_1.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.d5_1.a2._2_  (.I(\mult_u0.step2.add_sub4_u0.ppa8_u0.d5_1.a2._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.d5_1.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.d5_1.o2._1_  (.A1(\mult_u0.step2.add_sub4_u0.ppa8_u0.cg43 ),
    .A2(\mult_u0.step2.add_sub4_u0.ppa8_u0.d5_1.a2.out ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.d5_1.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.d5_1.o2._2_  (.I(\mult_u0.step2.add_sub4_u0.ppa8_u0.d5_1.o2._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.cg[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.d6_0.a1._1_  (.A1(\mult_u0.step2.add_sub4_u0.ppa8_u0.cp43 ),
    .A2(\mult_u0.step2.add_sub4_u0.ppa8_u0.d6_0.a1.in0 ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.d6_0.a1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.d6_0.a1._2_  (.I(\mult_u0.step2.add_sub4_u0.ppa8_u0.d6_0.a1._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.cp54 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.d6_0.a2._1_  (.A1(\mult_u0.step2.add_sub4_u0.ppa8_u0.cg43 ),
    .A2(\mult_u0.step2.add_sub4_u0.ppa8_u0.d6_0.a1.in0 ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.d6_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.d6_0.a2._2_  (.I(\mult_u0.step2.add_sub4_u0.ppa8_u0.d6_0.a2._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.d6_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.d6_0.o2._1_  (.A1(\mult_u0.step2.add_sub4_u0.ppa8_u0.d6_0.g1 ),
    .A2(\mult_u0.step2.add_sub4_u0.ppa8_u0.d6_0.a2.out ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.d6_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.d6_0.o2._2_  (.I(\mult_u0.step2.add_sub4_u0.ppa8_u0.d6_0.o2._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.cg54 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.d6_1.a2._1_  (.A1(\mult_u0.step2.add_sub4_u0.ppa8_u0.cg[2] ),
    .A2(\mult_u0.step2.add_sub4_u0.ppa8_u0.cp54 ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.d6_1.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.d6_1.a2._2_  (.I(\mult_u0.step2.add_sub4_u0.ppa8_u0.d6_1.a2._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.d6_1.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.d6_1.o2._1_  (.A1(\mult_u0.step2.add_sub4_u0.ppa8_u0.cg54 ),
    .A2(\mult_u0.step2.add_sub4_u0.ppa8_u0.d6_1.a2.out ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.d6_1.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.d6_1.o2._2_  (.I(\mult_u0.step2.add_sub4_u0.ppa8_u0.d6_1.o2._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.cg[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.p_0.a._1_  (.A1(\mult_u0.step2.add_sub4_u0.int_ip[0] ),
    .A2(\mult_u0.acc_s1[0] ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.p_0.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.p_0.a._2_  (.I(\mult_u0.step2.add_sub4_u0.ppa8_u0.p_0.a._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.d1_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.p_0.o._1_  (.A1(\mult_u0.step2.add_sub4_u0.int_ip[0] ),
    .A2(\mult_u0.acc_s1[0] ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.p_0.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.p_0.o._2_  (.I(\mult_u0.step2.add_sub4_u0.ppa8_u0.p_0.o._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.d1_0.a2.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.p_1.a._1_  (.A1(\mult_u0.step2.add_sub4_u0.int_ip[1] ),
    .A2(\mult_u0.acc_s1[1] ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.p_1.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.p_1.a._2_  (.I(\mult_u0.step2.add_sub4_u0.ppa8_u0.p_1.a._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.d2_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.p_1.o._1_  (.A1(\mult_u0.step2.add_sub4_u0.int_ip[1] ),
    .A2(\mult_u0.acc_s1[1] ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.p_1.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.p_1.o._2_  (.I(\mult_u0.step2.add_sub4_u0.ppa8_u0.p_1.o._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.p_2.a._1_  (.A1(\mult_u0.step2.add_sub4_u0.int_ip[2] ),
    .A2(\mult_u0.acc_s1[2] ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.p_2.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.p_2.a._2_  (.I(\mult_u0.step2.add_sub4_u0.ppa8_u0.p_2.a._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.d3_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.p_2.o._1_  (.A1(\mult_u0.step2.add_sub4_u0.int_ip[2] ),
    .A2(\mult_u0.acc_s1[2] ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.p_2.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.p_2.o._2_  (.I(\mult_u0.step2.add_sub4_u0.ppa8_u0.p_2.o._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.p_3.a._1_  (.A1(\mult_u0.step2.add_sub4_u0.int_ip[3] ),
    .A2(\mult_u0.acc_s1[3] ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.p_3.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.p_3.a._2_  (.I(\mult_u0.step2.add_sub4_u0.ppa8_u0.p_3.a._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.d4_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.p_3.o._1_  (.A1(\mult_u0.step2.add_sub4_u0.int_ip[3] ),
    .A2(\mult_u0.acc_s1[3] ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.p_3.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.p_3.o._2_  (.I(\mult_u0.step2.add_sub4_u0.ppa8_u0.p_3.o._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.d4_0.a2.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.p_4.a._1_  (.A1(\mult_u0.step2.add_sub4_u0.int_ip[4] ),
    .A2(\mult_u0.acc_s1[4] ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.p_4.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.p_4.a._2_  (.I(\mult_u0.step2.add_sub4_u0.ppa8_u0.p_4.a._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.d5_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.p_4.o._1_  (.A1(\mult_u0.step2.add_sub4_u0.int_ip[4] ),
    .A2(\mult_u0.acc_s1[4] ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.p_4.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.p_4.o._2_  (.I(\mult_u0.step2.add_sub4_u0.ppa8_u0.p_4.o._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.d5_0.a1.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.p_5.a._1_  (.A1(\mult_u0.step2.add_sub4_u0.int_ip[5] ),
    .A2(\mult_u0.acc_s1[5] ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.p_5.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.p_5.a._2_  (.I(\mult_u0.step2.add_sub4_u0.ppa8_u0.p_5.a._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.d6_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.p_5.o._1_  (.A1(\mult_u0.step2.add_sub4_u0.int_ip[5] ),
    .A2(\mult_u0.acc_s1[5] ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.p_5.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.p_5.o._2_  (.I(\mult_u0.step2.add_sub4_u0.ppa8_u0.p_5.o._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.d6_0.a1.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.s1.xor2_0._1_  (.A1(\mult_u0.step2.add_sub4_u0.int_ip[1] ),
    .A2(\mult_u0.acc_s1[1] ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.s1.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.s1.xor2_0._2_  (.I(\mult_u0.step2.add_sub4_u0.ppa8_u0.s1.xor2_0._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.s1.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.s1.xor2_1._1_  (.A1(\mult_u0.step2.add_sub4_u0.ppa8_u0.s1.temp ),
    .A2(\mult_u0.step2.add_sub4_u0.ppa8_u0.cg[0] ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.s1.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.s1.xor2_1._2_  (.I(\mult_u0.step2.add_sub4_u0.ppa8_u0.s1.xor2_1._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.S[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.s2.xor2_0._1_  (.A1(\mult_u0.step2.add_sub4_u0.int_ip[2] ),
    .A2(\mult_u0.acc_s1[2] ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.s2.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.s2.xor2_0._2_  (.I(\mult_u0.step2.add_sub4_u0.ppa8_u0.s2.xor2_0._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.s2.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.s2.xor2_1._1_  (.A1(\mult_u0.step2.add_sub4_u0.ppa8_u0.s2.temp ),
    .A2(\mult_u0.step2.add_sub4_u0.ppa8_u0.cg[1] ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.s2.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.s2.xor2_1._2_  (.I(\mult_u0.step2.add_sub4_u0.ppa8_u0.s2.xor2_1._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.S[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.s3.xor2_0._1_  (.A1(\mult_u0.step2.add_sub4_u0.int_ip[3] ),
    .A2(\mult_u0.acc_s1[3] ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.s3.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.s3.xor2_0._2_  (.I(\mult_u0.step2.add_sub4_u0.ppa8_u0.s3.xor2_0._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.s3.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.s3.xor2_1._1_  (.A1(\mult_u0.step2.add_sub4_u0.ppa8_u0.s3.temp ),
    .A2(\mult_u0.step2.add_sub4_u0.ppa8_u0.cg[2] ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.s3.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.s3.xor2_1._2_  (.I(\mult_u0.step2.add_sub4_u0.ppa8_u0.s3.xor2_1._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.S[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.s4.xor2_0._1_  (.A1(\mult_u0.step2.add_sub4_u0.int_ip[4] ),
    .A2(\mult_u0.acc_s1[4] ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.s4.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.s4.xor2_0._2_  (.I(\mult_u0.step2.add_sub4_u0.ppa8_u0.s4.xor2_0._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.s4.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.s4.xor2_1._1_  (.A1(\mult_u0.step2.add_sub4_u0.ppa8_u0.s4.temp ),
    .A2(\mult_u0.step2.add_sub4_u0.ppa8_u0.cg[3] ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.s4.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.s4.xor2_1._2_  (.I(\mult_u0.step2.add_sub4_u0.ppa8_u0.s4.xor2_1._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.S[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.s5.xor2_0._1_  (.A1(\mult_u0.step2.add_sub4_u0.int_ip[5] ),
    .A2(\mult_u0.acc_s1[5] ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.s5.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.s5.xor2_0._2_  (.I(\mult_u0.step2.add_sub4_u0.ppa8_u0.s5.xor2_0._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.s5.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.s5.xor2_1._1_  (.A1(\mult_u0.step2.add_sub4_u0.ppa8_u0.s5.temp ),
    .A2(\mult_u0.step2.add_sub4_u0.ppa8_u0.cg[4] ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.s5.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.s5.xor2_1._2_  (.I(\mult_u0.step2.add_sub4_u0.ppa8_u0.s5.xor2_1._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.S[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.s6.xor2_0._1_  (.A1(\mult_u0.step2.add_sub4_u0.int_ip[6] ),
    .A2(\mult_u0.acc_s1[6] ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.s6.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.s6.xor2_0._2_  (.I(\mult_u0.step2.add_sub4_u0.ppa8_u0.s6.xor2_0._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.s6.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.s6.xor2_1._1_  (.A1(\mult_u0.step2.add_sub4_u0.ppa8_u0.s6.temp ),
    .A2(\mult_u0.step2.add_sub4_u0.ppa8_u0.cg[5] ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.s6.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.ppa8_u0.s6.xor2_1._2_  (.I(\mult_u0.step2.add_sub4_u0.ppa8_u0.s6.xor2_1._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.ppa8_u0.S[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step2.add_sub4_u0.x0._1_  (.A1(\mult_u0.Q_s1[0] ),
    .A2(\mult_u0.multiplicand_s1[0] ),
    .Z(\mult_u0.step2.add_sub4_u0.x0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.x0._2_  (.I(\mult_u0.step2.add_sub4_u0.x0._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.int_ip[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step2.add_sub4_u0.x1._1_  (.A1(\mult_u0.Q_s1[0] ),
    .A2(\mult_u0.multiplicand_s1[1] ),
    .Z(\mult_u0.step2.add_sub4_u0.x1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.x1._2_  (.I(\mult_u0.step2.add_sub4_u0.x1._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.int_ip[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step2.add_sub4_u0.x2._1_  (.A1(\mult_u0.Q_s1[0] ),
    .A2(\mult_u0.multiplicand_s1[2] ),
    .Z(\mult_u0.step2.add_sub4_u0.x2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.x2._2_  (.I(\mult_u0.step2.add_sub4_u0.x2._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.int_ip[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step2.add_sub4_u0.x3._1_  (.A1(\mult_u0.Q_s1[0] ),
    .A2(\mult_u0.multiplicand_s1[3] ),
    .Z(\mult_u0.step2.add_sub4_u0.x3._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.x3._2_  (.I(\mult_u0.step2.add_sub4_u0.x3._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.int_ip[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step2.add_sub4_u0.x4._1_  (.A1(\mult_u0.Q_s1[0] ),
    .A2(\mult_u0.multiplicand_s1[4] ),
    .Z(\mult_u0.step2.add_sub4_u0.x4._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.x4._2_  (.I(\mult_u0.step2.add_sub4_u0.x4._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.int_ip[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step2.add_sub4_u0.x5._1_  (.A1(\mult_u0.Q_s1[0] ),
    .A2(\mult_u0.multiplicand_s1[5] ),
    .Z(\mult_u0.step2.add_sub4_u0.x5._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.x5._2_  (.I(\mult_u0.step2.add_sub4_u0.x5._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.int_ip[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step2.add_sub4_u0.x6._1_  (.A1(\mult_u0.Q_s1[0] ),
    .A2(\mult_u0.multiplicand_s1[6] ),
    .Z(\mult_u0.step2.add_sub4_u0.x6._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step2.add_sub4_u0.x6._2_  (.I(\mult_u0.step2.add_sub4_u0.x6._0_ ),
    .Z(\mult_u0.step2.add_sub4_u0.int_ip[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step3._09_  (.A1(\mult_u0.q0_s2 ),
    .A2(\mult_u0.Q_s2[0] ),
    .Z(\mult_u0.step3._00_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 \mult_u0.step3._10_  (.I(\mult_u0.step3._00_ ),
    .Z(\mult_u0.step3._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_u0.step3._11_  (.I0(\mult_u0.acc_s2[6] ),
    .I1(\mult_u0.step3.add_sub4_u0.ppa8_u0.S[6] ),
    .S(\mult_u0.step3._01_ ),
    .Z(\mult_u0.step3._02_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3._12_  (.I(\mult_u0.step3._02_ ),
    .Z(\mult_u0.acc[3][6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_u0.step3._13_  (.I0(\mult_u0.acc_s2[1] ),
    .I1(\mult_u0.step3.add_sub4_u0.ppa8_u0.S[1] ),
    .S(\mult_u0.step3._01_ ),
    .Z(\mult_u0.step3._03_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3._14_  (.I(\mult_u0.step3._03_ ),
    .Z(\mult_u0.acc[3][0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_u0.step3._15_  (.I0(\mult_u0.acc_s2[2] ),
    .I1(\mult_u0.step3.add_sub4_u0.ppa8_u0.S[2] ),
    .S(\mult_u0.step3._01_ ),
    .Z(\mult_u0.step3._04_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3._16_  (.I(\mult_u0.step3._04_ ),
    .Z(\mult_u0.acc[3][1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_u0.step3._17_  (.I0(\mult_u0.acc_s2[3] ),
    .I1(\mult_u0.step3.add_sub4_u0.ppa8_u0.S[3] ),
    .S(\mult_u0.step3._01_ ),
    .Z(\mult_u0.step3._05_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3._18_  (.I(\mult_u0.step3._05_ ),
    .Z(\mult_u0.acc[3][2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_u0.step3._19_  (.I0(\mult_u0.acc_s2[4] ),
    .I1(\mult_u0.step3.add_sub4_u0.ppa8_u0.S[4] ),
    .S(\mult_u0.step3._01_ ),
    .Z(\mult_u0.step3._06_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3._20_  (.I(\mult_u0.step3._06_ ),
    .Z(\mult_u0.acc[3][3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_u0.step3._21_  (.I0(\mult_u0.acc_s2[5] ),
    .I1(\mult_u0.step3.add_sub4_u0.ppa8_u0.S[5] ),
    .S(\mult_u0.step3._01_ ),
    .Z(\mult_u0.step3._07_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3._22_  (.I(\mult_u0.step3._07_ ),
    .Z(\mult_u0.acc[3][4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3._25_  (.I(\mult_u0.Q_s2[1] ),
    .Z(\mult_u0.Q[2][0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3._26_  (.I(\mult_u0.Q_s2[2] ),
    .Z(\mult_u0.Q[2][1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3._27_  (.I(\mult_u0.Q_s2[3] ),
    .Z(\mult_u0.Q[2][2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3._28_  (.I(\mult_u0.Q_s2[4] ),
    .Z(\mult_u0.Q[2][3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3._31_  (.I(\mult_u0.acc[3][6] ),
    .Z(\mult_u0.acc[3][5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3._32_  (.I(\mult_u0.Q_s2[0] ),
    .Z(\mult_u0.q0[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.d1_0.a2._1_  (.A1(\mult_u0.Q_s2[0] ),
    .A2(\mult_u0.step3.add_sub4_u0.ppa8_u0.d1_0.a2.in0 ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.d1_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.d1_0.a2._2_  (.I(\mult_u0.step3.add_sub4_u0.ppa8_u0.d1_0.a2._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.d1_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.d1_0.o2._1_  (.A1(\mult_u0.step3.add_sub4_u0.ppa8_u0.d1_0.g1 ),
    .A2(\mult_u0.step3.add_sub4_u0.ppa8_u0.d1_0.a2.out ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.d1_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.d1_0.o2._2_  (.I(\mult_u0.step3.add_sub4_u0.ppa8_u0.d1_0.o2._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.cg[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.d2_0.a2._1_  (.A1(\mult_u0.step3.add_sub4_u0.ppa8_u0.cg[0] ),
    .A2(\mult_u0.step3.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.d2_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.d2_0.a2._2_  (.I(\mult_u0.step3.add_sub4_u0.ppa8_u0.d2_0.a2._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.d2_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.d2_0.o2._1_  (.A1(\mult_u0.step3.add_sub4_u0.ppa8_u0.d2_0.g1 ),
    .A2(\mult_u0.step3.add_sub4_u0.ppa8_u0.d2_0.a2.out ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.d2_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.d2_0.o2._2_  (.I(\mult_u0.step3.add_sub4_u0.ppa8_u0.d2_0.o2._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.cg[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.d3_0.a1._1_  (.A1(\mult_u0.step3.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ),
    .A2(\mult_u0.step3.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.d3_0.a1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.d3_0.a1._2_  (.I(\mult_u0.step3.add_sub4_u0.ppa8_u0.d3_0.a1._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.cp21 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.d3_0.a2._1_  (.A1(\mult_u0.step3.add_sub4_u0.ppa8_u0.d2_0.g1 ),
    .A2(\mult_u0.step3.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.d3_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.d3_0.a2._2_  (.I(\mult_u0.step3.add_sub4_u0.ppa8_u0.d3_0.a2._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.d3_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.d3_0.o2._1_  (.A1(\mult_u0.step3.add_sub4_u0.ppa8_u0.d3_0.g1 ),
    .A2(\mult_u0.step3.add_sub4_u0.ppa8_u0.d3_0.a2.out ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.d3_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.d3_0.o2._2_  (.I(\mult_u0.step3.add_sub4_u0.ppa8_u0.d3_0.o2._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.cg21 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.d3_1.a2._1_  (.A1(\mult_u0.step3.add_sub4_u0.ppa8_u0.cg[0] ),
    .A2(\mult_u0.step3.add_sub4_u0.ppa8_u0.cp21 ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.d3_1.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.d3_1.a2._2_  (.I(\mult_u0.step3.add_sub4_u0.ppa8_u0.d3_1.a2._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.d3_1.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.d3_1.o2._1_  (.A1(\mult_u0.step3.add_sub4_u0.ppa8_u0.cg21 ),
    .A2(\mult_u0.step3.add_sub4_u0.ppa8_u0.d3_1.a2.out ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.d3_1.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.d3_1.o2._2_  (.I(\mult_u0.step3.add_sub4_u0.ppa8_u0.d3_1.o2._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.cg[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.d4_0.a2._1_  (.A1(\mult_u0.step3.add_sub4_u0.ppa8_u0.cg[2] ),
    .A2(\mult_u0.step3.add_sub4_u0.ppa8_u0.d4_0.a2.in0 ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.d4_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.d4_0.a2._2_  (.I(\mult_u0.step3.add_sub4_u0.ppa8_u0.d4_0.a2._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.d4_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.d4_0.o2._1_  (.A1(\mult_u0.step3.add_sub4_u0.ppa8_u0.d4_0.g1 ),
    .A2(\mult_u0.step3.add_sub4_u0.ppa8_u0.d4_0.a2.out ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.d4_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.d4_0.o2._2_  (.I(\mult_u0.step3.add_sub4_u0.ppa8_u0.d4_0.o2._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.cg[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.d5_0.a1._1_  (.A1(\mult_u0.step3.add_sub4_u0.ppa8_u0.d4_0.a2.in0 ),
    .A2(\mult_u0.step3.add_sub4_u0.ppa8_u0.d5_0.a1.in0 ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.d5_0.a1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.d5_0.a1._2_  (.I(\mult_u0.step3.add_sub4_u0.ppa8_u0.d5_0.a1._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.cp43 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.d5_0.a2._1_  (.A1(\mult_u0.step3.add_sub4_u0.ppa8_u0.d4_0.g1 ),
    .A2(\mult_u0.step3.add_sub4_u0.ppa8_u0.d5_0.a1.in0 ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.d5_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.d5_0.a2._2_  (.I(\mult_u0.step3.add_sub4_u0.ppa8_u0.d5_0.a2._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.d5_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.d5_0.o2._1_  (.A1(\mult_u0.step3.add_sub4_u0.ppa8_u0.d5_0.g1 ),
    .A2(\mult_u0.step3.add_sub4_u0.ppa8_u0.d5_0.a2.out ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.d5_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.d5_0.o2._2_  (.I(\mult_u0.step3.add_sub4_u0.ppa8_u0.d5_0.o2._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.cg43 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.d5_1.a2._1_  (.A1(\mult_u0.step3.add_sub4_u0.ppa8_u0.cg[2] ),
    .A2(\mult_u0.step3.add_sub4_u0.ppa8_u0.cp43 ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.d5_1.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.d5_1.a2._2_  (.I(\mult_u0.step3.add_sub4_u0.ppa8_u0.d5_1.a2._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.d5_1.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.d5_1.o2._1_  (.A1(\mult_u0.step3.add_sub4_u0.ppa8_u0.cg43 ),
    .A2(\mult_u0.step3.add_sub4_u0.ppa8_u0.d5_1.a2.out ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.d5_1.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.d5_1.o2._2_  (.I(\mult_u0.step3.add_sub4_u0.ppa8_u0.d5_1.o2._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.cg[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.d6_0.a1._1_  (.A1(\mult_u0.step3.add_sub4_u0.ppa8_u0.cp43 ),
    .A2(\mult_u0.step3.add_sub4_u0.ppa8_u0.d6_0.a1.in0 ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.d6_0.a1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.d6_0.a1._2_  (.I(\mult_u0.step3.add_sub4_u0.ppa8_u0.d6_0.a1._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.cp54 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.d6_0.a2._1_  (.A1(\mult_u0.step3.add_sub4_u0.ppa8_u0.cg43 ),
    .A2(\mult_u0.step3.add_sub4_u0.ppa8_u0.d6_0.a1.in0 ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.d6_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.d6_0.a2._2_  (.I(\mult_u0.step3.add_sub4_u0.ppa8_u0.d6_0.a2._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.d6_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.d6_0.o2._1_  (.A1(\mult_u0.step3.add_sub4_u0.ppa8_u0.d6_0.g1 ),
    .A2(\mult_u0.step3.add_sub4_u0.ppa8_u0.d6_0.a2.out ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.d6_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.d6_0.o2._2_  (.I(\mult_u0.step3.add_sub4_u0.ppa8_u0.d6_0.o2._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.cg54 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.d6_1.a2._1_  (.A1(\mult_u0.step3.add_sub4_u0.ppa8_u0.cg[2] ),
    .A2(\mult_u0.step3.add_sub4_u0.ppa8_u0.cp54 ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.d6_1.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.d6_1.a2._2_  (.I(\mult_u0.step3.add_sub4_u0.ppa8_u0.d6_1.a2._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.d6_1.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.d6_1.o2._1_  (.A1(\mult_u0.step3.add_sub4_u0.ppa8_u0.cg54 ),
    .A2(\mult_u0.step3.add_sub4_u0.ppa8_u0.d6_1.a2.out ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.d6_1.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.d6_1.o2._2_  (.I(\mult_u0.step3.add_sub4_u0.ppa8_u0.d6_1.o2._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.cg[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.p_0.a._1_  (.A1(\mult_u0.step3.add_sub4_u0.int_ip[0] ),
    .A2(\mult_u0.acc_s2[0] ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.p_0.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.p_0.a._2_  (.I(\mult_u0.step3.add_sub4_u0.ppa8_u0.p_0.a._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.d1_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.p_0.o._1_  (.A1(\mult_u0.step3.add_sub4_u0.int_ip[0] ),
    .A2(\mult_u0.acc_s2[0] ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.p_0.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.p_0.o._2_  (.I(\mult_u0.step3.add_sub4_u0.ppa8_u0.p_0.o._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.d1_0.a2.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.p_1.a._1_  (.A1(\mult_u0.step3.add_sub4_u0.int_ip[1] ),
    .A2(\mult_u0.acc_s2[1] ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.p_1.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.p_1.a._2_  (.I(\mult_u0.step3.add_sub4_u0.ppa8_u0.p_1.a._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.d2_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.p_1.o._1_  (.A1(\mult_u0.step3.add_sub4_u0.int_ip[1] ),
    .A2(\mult_u0.acc_s2[1] ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.p_1.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.p_1.o._2_  (.I(\mult_u0.step3.add_sub4_u0.ppa8_u0.p_1.o._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.p_2.a._1_  (.A1(\mult_u0.step3.add_sub4_u0.int_ip[2] ),
    .A2(\mult_u0.acc_s2[2] ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.p_2.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.p_2.a._2_  (.I(\mult_u0.step3.add_sub4_u0.ppa8_u0.p_2.a._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.d3_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.p_2.o._1_  (.A1(\mult_u0.step3.add_sub4_u0.int_ip[2] ),
    .A2(\mult_u0.acc_s2[2] ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.p_2.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.p_2.o._2_  (.I(\mult_u0.step3.add_sub4_u0.ppa8_u0.p_2.o._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.p_3.a._1_  (.A1(\mult_u0.step3.add_sub4_u0.int_ip[3] ),
    .A2(\mult_u0.acc_s2[3] ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.p_3.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.p_3.a._2_  (.I(\mult_u0.step3.add_sub4_u0.ppa8_u0.p_3.a._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.d4_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.p_3.o._1_  (.A1(\mult_u0.step3.add_sub4_u0.int_ip[3] ),
    .A2(\mult_u0.acc_s2[3] ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.p_3.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.p_3.o._2_  (.I(\mult_u0.step3.add_sub4_u0.ppa8_u0.p_3.o._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.d4_0.a2.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.p_4.a._1_  (.A1(\mult_u0.step3.add_sub4_u0.int_ip[4] ),
    .A2(\mult_u0.acc_s2[4] ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.p_4.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.p_4.a._2_  (.I(\mult_u0.step3.add_sub4_u0.ppa8_u0.p_4.a._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.d5_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.p_4.o._1_  (.A1(\mult_u0.step3.add_sub4_u0.int_ip[4] ),
    .A2(\mult_u0.acc_s2[4] ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.p_4.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.p_4.o._2_  (.I(\mult_u0.step3.add_sub4_u0.ppa8_u0.p_4.o._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.d5_0.a1.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.p_5.a._1_  (.A1(\mult_u0.step3.add_sub4_u0.int_ip[5] ),
    .A2(\mult_u0.acc_s2[5] ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.p_5.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.p_5.a._2_  (.I(\mult_u0.step3.add_sub4_u0.ppa8_u0.p_5.a._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.d6_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.p_5.o._1_  (.A1(\mult_u0.step3.add_sub4_u0.int_ip[5] ),
    .A2(\mult_u0.acc_s2[5] ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.p_5.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.p_5.o._2_  (.I(\mult_u0.step3.add_sub4_u0.ppa8_u0.p_5.o._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.d6_0.a1.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.s1.xor2_0._1_  (.A1(\mult_u0.step3.add_sub4_u0.int_ip[1] ),
    .A2(\mult_u0.acc_s2[1] ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.s1.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.s1.xor2_0._2_  (.I(\mult_u0.step3.add_sub4_u0.ppa8_u0.s1.xor2_0._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.s1.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.s1.xor2_1._1_  (.A1(\mult_u0.step3.add_sub4_u0.ppa8_u0.s1.temp ),
    .A2(\mult_u0.step3.add_sub4_u0.ppa8_u0.cg[0] ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.s1.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.s1.xor2_1._2_  (.I(\mult_u0.step3.add_sub4_u0.ppa8_u0.s1.xor2_1._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.S[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.s2.xor2_0._1_  (.A1(\mult_u0.step3.add_sub4_u0.int_ip[2] ),
    .A2(\mult_u0.acc_s2[2] ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.s2.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.s2.xor2_0._2_  (.I(\mult_u0.step3.add_sub4_u0.ppa8_u0.s2.xor2_0._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.s2.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.s2.xor2_1._1_  (.A1(\mult_u0.step3.add_sub4_u0.ppa8_u0.s2.temp ),
    .A2(\mult_u0.step3.add_sub4_u0.ppa8_u0.cg[1] ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.s2.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.s2.xor2_1._2_  (.I(\mult_u0.step3.add_sub4_u0.ppa8_u0.s2.xor2_1._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.S[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.s3.xor2_0._1_  (.A1(\mult_u0.step3.add_sub4_u0.int_ip[3] ),
    .A2(\mult_u0.acc_s2[3] ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.s3.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.s3.xor2_0._2_  (.I(\mult_u0.step3.add_sub4_u0.ppa8_u0.s3.xor2_0._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.s3.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.s3.xor2_1._1_  (.A1(\mult_u0.step3.add_sub4_u0.ppa8_u0.s3.temp ),
    .A2(\mult_u0.step3.add_sub4_u0.ppa8_u0.cg[2] ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.s3.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.s3.xor2_1._2_  (.I(\mult_u0.step3.add_sub4_u0.ppa8_u0.s3.xor2_1._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.S[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.s4.xor2_0._1_  (.A1(\mult_u0.step3.add_sub4_u0.int_ip[4] ),
    .A2(\mult_u0.acc_s2[4] ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.s4.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.s4.xor2_0._2_  (.I(\mult_u0.step3.add_sub4_u0.ppa8_u0.s4.xor2_0._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.s4.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.s4.xor2_1._1_  (.A1(\mult_u0.step3.add_sub4_u0.ppa8_u0.s4.temp ),
    .A2(\mult_u0.step3.add_sub4_u0.ppa8_u0.cg[3] ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.s4.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.s4.xor2_1._2_  (.I(\mult_u0.step3.add_sub4_u0.ppa8_u0.s4.xor2_1._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.S[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.s5.xor2_0._1_  (.A1(\mult_u0.step3.add_sub4_u0.int_ip[5] ),
    .A2(\mult_u0.acc_s2[5] ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.s5.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.s5.xor2_0._2_  (.I(\mult_u0.step3.add_sub4_u0.ppa8_u0.s5.xor2_0._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.s5.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.s5.xor2_1._1_  (.A1(\mult_u0.step3.add_sub4_u0.ppa8_u0.s5.temp ),
    .A2(\mult_u0.step3.add_sub4_u0.ppa8_u0.cg[4] ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.s5.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.s5.xor2_1._2_  (.I(\mult_u0.step3.add_sub4_u0.ppa8_u0.s5.xor2_1._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.S[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.s6.xor2_0._1_  (.A1(\mult_u0.step3.add_sub4_u0.int_ip[6] ),
    .A2(\mult_u0.acc_s2[6] ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.s6.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.s6.xor2_0._2_  (.I(\mult_u0.step3.add_sub4_u0.ppa8_u0.s6.xor2_0._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.s6.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.s6.xor2_1._1_  (.A1(\mult_u0.step3.add_sub4_u0.ppa8_u0.s6.temp ),
    .A2(\mult_u0.step3.add_sub4_u0.ppa8_u0.cg[5] ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.s6.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.ppa8_u0.s6.xor2_1._2_  (.I(\mult_u0.step3.add_sub4_u0.ppa8_u0.s6.xor2_1._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.ppa8_u0.S[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step3.add_sub4_u0.x0._1_  (.A1(\mult_u0.Q_s2[0] ),
    .A2(\mult_u0.multiplicand_s2[0] ),
    .Z(\mult_u0.step3.add_sub4_u0.x0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.x0._2_  (.I(\mult_u0.step3.add_sub4_u0.x0._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.int_ip[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step3.add_sub4_u0.x1._1_  (.A1(\mult_u0.Q_s2[0] ),
    .A2(\mult_u0.multiplicand_s2[1] ),
    .Z(\mult_u0.step3.add_sub4_u0.x1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.x1._2_  (.I(\mult_u0.step3.add_sub4_u0.x1._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.int_ip[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step3.add_sub4_u0.x2._1_  (.A1(\mult_u0.Q_s2[0] ),
    .A2(\mult_u0.multiplicand_s2[2] ),
    .Z(\mult_u0.step3.add_sub4_u0.x2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.x2._2_  (.I(\mult_u0.step3.add_sub4_u0.x2._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.int_ip[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step3.add_sub4_u0.x3._1_  (.A1(\mult_u0.Q_s2[0] ),
    .A2(\mult_u0.multiplicand_s2[3] ),
    .Z(\mult_u0.step3.add_sub4_u0.x3._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.x3._2_  (.I(\mult_u0.step3.add_sub4_u0.x3._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.int_ip[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step3.add_sub4_u0.x4._1_  (.A1(\mult_u0.Q_s2[0] ),
    .A2(\mult_u0.multiplicand_s2[4] ),
    .Z(\mult_u0.step3.add_sub4_u0.x4._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.x4._2_  (.I(\mult_u0.step3.add_sub4_u0.x4._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.int_ip[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step3.add_sub4_u0.x5._1_  (.A1(\mult_u0.Q_s2[0] ),
    .A2(\mult_u0.multiplicand_s2[5] ),
    .Z(\mult_u0.step3.add_sub4_u0.x5._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.x5._2_  (.I(\mult_u0.step3.add_sub4_u0.x5._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.int_ip[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step3.add_sub4_u0.x6._1_  (.A1(\mult_u0.Q_s2[0] ),
    .A2(\mult_u0.multiplicand_s2[6] ),
    .Z(\mult_u0.step3.add_sub4_u0.x6._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step3.add_sub4_u0.x6._2_  (.I(\mult_u0.step3.add_sub4_u0.x6._0_ ),
    .Z(\mult_u0.step3.add_sub4_u0.int_ip[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step4._09_  (.A1(\mult_u0.q0_s3 ),
    .A2(\mult_u0.Q_s3[0] ),
    .Z(\mult_u0.step4._00_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 \mult_u0.step4._10_  (.I(\mult_u0.step4._00_ ),
    .Z(\mult_u0.step4._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_u0.step4._11_  (.I0(\mult_u0.acc_s3[6] ),
    .I1(\mult_u0.step4.add_sub4_u0.ppa8_u0.S[6] ),
    .S(\mult_u0.step4._01_ ),
    .Z(\mult_u0.step4._02_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4._12_  (.I(\mult_u0.step4._02_ ),
    .Z(\mult_u0.acc[4][6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_u0.step4._13_  (.I0(\mult_u0.acc_s3[1] ),
    .I1(\mult_u0.step4.add_sub4_u0.ppa8_u0.S[1] ),
    .S(\mult_u0.step4._01_ ),
    .Z(\mult_u0.step4._03_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4._14_  (.I(\mult_u0.step4._03_ ),
    .Z(\mult_u0.acc[4][0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_u0.step4._15_  (.I0(\mult_u0.acc_s3[2] ),
    .I1(\mult_u0.step4.add_sub4_u0.ppa8_u0.S[2] ),
    .S(\mult_u0.step4._01_ ),
    .Z(\mult_u0.step4._04_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4._16_  (.I(\mult_u0.step4._04_ ),
    .Z(\mult_u0.acc[4][1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_u0.step4._17_  (.I0(\mult_u0.acc_s3[3] ),
    .I1(\mult_u0.step4.add_sub4_u0.ppa8_u0.S[3] ),
    .S(\mult_u0.step4._01_ ),
    .Z(\mult_u0.step4._05_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4._18_  (.I(\mult_u0.step4._05_ ),
    .Z(\mult_u0.acc[4][2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_u0.step4._19_  (.I0(\mult_u0.acc_s3[4] ),
    .I1(\mult_u0.step4.add_sub4_u0.ppa8_u0.S[4] ),
    .S(\mult_u0.step4._01_ ),
    .Z(\mult_u0.step4._06_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4._20_  (.I(\mult_u0.step4._06_ ),
    .Z(\mult_u0.acc[4][3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_u0.step4._21_  (.I0(\mult_u0.acc_s3[5] ),
    .I1(\mult_u0.step4.add_sub4_u0.ppa8_u0.S[5] ),
    .S(\mult_u0.step4._01_ ),
    .Z(\mult_u0.step4._07_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4._22_  (.I(\mult_u0.step4._07_ ),
    .Z(\mult_u0.acc[4][4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_u0.step4._23_  (.I0(\mult_u0.acc_s3[0] ),
    .I1(\mult_u0.step4.add_sub4_u0.ppa8_u0.S[0] ),
    .S(\mult_u0.step4._01_ ),
    .Z(\mult_u0.step4._08_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4._24_  (.I(\mult_u0.step4._08_ ),
    .Z(\mult_u0.Q[3][6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4._25_  (.I(\mult_u0.Q_s3[1] ),
    .Z(\mult_u0.Q[3][0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4._26_  (.I(\mult_u0.Q_s3[2] ),
    .Z(\mult_u0.Q[3][1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4._27_  (.I(\mult_u0.Q_s3[3] ),
    .Z(\mult_u0.Q[3][2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4._31_  (.I(\mult_u0.acc[4][6] ),
    .Z(\mult_u0.acc[4][5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4._32_  (.I(\mult_u0.Q_s3[0] ),
    .Z(\mult_u0.q0[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.d1_0.a2._1_  (.A1(\mult_u0.Q_s3[0] ),
    .A2(\mult_u0.step4.add_sub4_u0.ppa8_u0.d1_0.a2.in0 ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.d1_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.d1_0.a2._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.d1_0.a2._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.d1_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.d1_0.o2._1_  (.A1(\mult_u0.step4.add_sub4_u0.ppa8_u0.d1_0.g1 ),
    .A2(\mult_u0.step4.add_sub4_u0.ppa8_u0.d1_0.a2.out ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.d1_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.d1_0.o2._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.d1_0.o2._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.cg[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.d2_0.a2._1_  (.A1(\mult_u0.step4.add_sub4_u0.ppa8_u0.cg[0] ),
    .A2(\mult_u0.step4.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.d2_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.d2_0.a2._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.d2_0.a2._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.d2_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.d2_0.o2._1_  (.A1(\mult_u0.step4.add_sub4_u0.ppa8_u0.d2_0.g1 ),
    .A2(\mult_u0.step4.add_sub4_u0.ppa8_u0.d2_0.a2.out ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.d2_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.d2_0.o2._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.d2_0.o2._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.cg[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.d3_0.a1._1_  (.A1(\mult_u0.step4.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ),
    .A2(\mult_u0.step4.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.d3_0.a1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.d3_0.a1._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.d3_0.a1._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.cp21 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.d3_0.a2._1_  (.A1(\mult_u0.step4.add_sub4_u0.ppa8_u0.d2_0.g1 ),
    .A2(\mult_u0.step4.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.d3_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.d3_0.a2._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.d3_0.a2._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.d3_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.d3_0.o2._1_  (.A1(\mult_u0.step4.add_sub4_u0.ppa8_u0.d3_0.g1 ),
    .A2(\mult_u0.step4.add_sub4_u0.ppa8_u0.d3_0.a2.out ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.d3_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.d3_0.o2._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.d3_0.o2._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.cg21 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.d3_1.a2._1_  (.A1(\mult_u0.step4.add_sub4_u0.ppa8_u0.cg[0] ),
    .A2(\mult_u0.step4.add_sub4_u0.ppa8_u0.cp21 ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.d3_1.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.d3_1.a2._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.d3_1.a2._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.d3_1.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.d3_1.o2._1_  (.A1(\mult_u0.step4.add_sub4_u0.ppa8_u0.cg21 ),
    .A2(\mult_u0.step4.add_sub4_u0.ppa8_u0.d3_1.a2.out ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.d3_1.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.d3_1.o2._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.d3_1.o2._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.cg[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.d4_0.a2._1_  (.A1(\mult_u0.step4.add_sub4_u0.ppa8_u0.cg[2] ),
    .A2(\mult_u0.step4.add_sub4_u0.ppa8_u0.d4_0.a2.in0 ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.d4_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.d4_0.a2._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.d4_0.a2._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.d4_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.d4_0.o2._1_  (.A1(\mult_u0.step4.add_sub4_u0.ppa8_u0.d4_0.g1 ),
    .A2(\mult_u0.step4.add_sub4_u0.ppa8_u0.d4_0.a2.out ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.d4_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.d4_0.o2._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.d4_0.o2._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.cg[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.d5_0.a1._1_  (.A1(\mult_u0.step4.add_sub4_u0.ppa8_u0.d4_0.a2.in0 ),
    .A2(\mult_u0.step4.add_sub4_u0.ppa8_u0.d5_0.a1.in0 ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.d5_0.a1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.d5_0.a1._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.d5_0.a1._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.cp43 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.d5_0.a2._1_  (.A1(\mult_u0.step4.add_sub4_u0.ppa8_u0.d4_0.g1 ),
    .A2(\mult_u0.step4.add_sub4_u0.ppa8_u0.d5_0.a1.in0 ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.d5_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.d5_0.a2._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.d5_0.a2._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.d5_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.d5_0.o2._1_  (.A1(\mult_u0.step4.add_sub4_u0.ppa8_u0.d5_0.g1 ),
    .A2(\mult_u0.step4.add_sub4_u0.ppa8_u0.d5_0.a2.out ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.d5_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.d5_0.o2._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.d5_0.o2._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.cg43 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.d5_1.a2._1_  (.A1(\mult_u0.step4.add_sub4_u0.ppa8_u0.cg[2] ),
    .A2(\mult_u0.step4.add_sub4_u0.ppa8_u0.cp43 ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.d5_1.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.d5_1.a2._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.d5_1.a2._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.d5_1.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.d5_1.o2._1_  (.A1(\mult_u0.step4.add_sub4_u0.ppa8_u0.cg43 ),
    .A2(\mult_u0.step4.add_sub4_u0.ppa8_u0.d5_1.a2.out ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.d5_1.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.d5_1.o2._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.d5_1.o2._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.cg[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.d6_0.a1._1_  (.A1(\mult_u0.step4.add_sub4_u0.ppa8_u0.cp43 ),
    .A2(\mult_u0.step4.add_sub4_u0.ppa8_u0.d6_0.a1.in0 ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.d6_0.a1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.d6_0.a1._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.d6_0.a1._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.cp54 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.d6_0.a2._1_  (.A1(\mult_u0.step4.add_sub4_u0.ppa8_u0.cg43 ),
    .A2(\mult_u0.step4.add_sub4_u0.ppa8_u0.d6_0.a1.in0 ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.d6_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.d6_0.a2._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.d6_0.a2._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.d6_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.d6_0.o2._1_  (.A1(\mult_u0.step4.add_sub4_u0.ppa8_u0.d6_0.g1 ),
    .A2(\mult_u0.step4.add_sub4_u0.ppa8_u0.d6_0.a2.out ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.d6_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.d6_0.o2._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.d6_0.o2._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.cg54 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.d6_1.a2._1_  (.A1(\mult_u0.step4.add_sub4_u0.ppa8_u0.cg[2] ),
    .A2(\mult_u0.step4.add_sub4_u0.ppa8_u0.cp54 ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.d6_1.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.d6_1.a2._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.d6_1.a2._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.d6_1.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.d6_1.o2._1_  (.A1(\mult_u0.step4.add_sub4_u0.ppa8_u0.cg54 ),
    .A2(\mult_u0.step4.add_sub4_u0.ppa8_u0.d6_1.a2.out ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.d6_1.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.d6_1.o2._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.d6_1.o2._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.cg[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.p_0.a._1_  (.A1(\mult_u0.step4.add_sub4_u0.int_ip[0] ),
    .A2(\mult_u0.acc_s3[0] ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.p_0.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.p_0.a._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.p_0.a._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.d1_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.p_0.o._1_  (.A1(\mult_u0.step4.add_sub4_u0.int_ip[0] ),
    .A2(\mult_u0.acc_s3[0] ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.p_0.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.p_0.o._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.p_0.o._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.d1_0.a2.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.p_1.a._1_  (.A1(\mult_u0.step4.add_sub4_u0.int_ip[1] ),
    .A2(\mult_u0.acc_s3[1] ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.p_1.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.p_1.a._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.p_1.a._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.d2_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.p_1.o._1_  (.A1(\mult_u0.step4.add_sub4_u0.int_ip[1] ),
    .A2(\mult_u0.acc_s3[1] ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.p_1.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.p_1.o._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.p_1.o._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.p_2.a._1_  (.A1(\mult_u0.step4.add_sub4_u0.int_ip[2] ),
    .A2(\mult_u0.acc_s3[2] ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.p_2.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.p_2.a._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.p_2.a._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.d3_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.p_2.o._1_  (.A1(\mult_u0.step4.add_sub4_u0.int_ip[2] ),
    .A2(\mult_u0.acc_s3[2] ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.p_2.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.p_2.o._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.p_2.o._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.p_3.a._1_  (.A1(\mult_u0.step4.add_sub4_u0.int_ip[3] ),
    .A2(\mult_u0.acc_s3[3] ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.p_3.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.p_3.a._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.p_3.a._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.d4_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.p_3.o._1_  (.A1(\mult_u0.step4.add_sub4_u0.int_ip[3] ),
    .A2(\mult_u0.acc_s3[3] ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.p_3.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.p_3.o._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.p_3.o._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.d4_0.a2.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.p_4.a._1_  (.A1(\mult_u0.step4.add_sub4_u0.int_ip[4] ),
    .A2(\mult_u0.acc_s3[4] ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.p_4.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.p_4.a._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.p_4.a._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.d5_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.p_4.o._1_  (.A1(\mult_u0.step4.add_sub4_u0.int_ip[4] ),
    .A2(\mult_u0.acc_s3[4] ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.p_4.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.p_4.o._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.p_4.o._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.d5_0.a1.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.p_5.a._1_  (.A1(\mult_u0.step4.add_sub4_u0.int_ip[5] ),
    .A2(\mult_u0.acc_s3[5] ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.p_5.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.p_5.a._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.p_5.a._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.d6_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.p_5.o._1_  (.A1(\mult_u0.step4.add_sub4_u0.int_ip[5] ),
    .A2(\mult_u0.acc_s3[5] ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.p_5.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.p_5.o._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.p_5.o._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.d6_0.a1.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.s0.xor2_0._1_  (.A1(\mult_u0.step4.add_sub4_u0.int_ip[0] ),
    .A2(\mult_u0.acc_s3[0] ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.s0.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.s0.xor2_0._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.s0.xor2_0._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.s0.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.s0.xor2_1._1_  (.A1(\mult_u0.step4.add_sub4_u0.ppa8_u0.s0.temp ),
    .A2(\mult_u0.Q_s3[0] ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.s0.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.s0.xor2_1._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.s0.xor2_1._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.S[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.s1.xor2_0._1_  (.A1(\mult_u0.step4.add_sub4_u0.int_ip[1] ),
    .A2(\mult_u0.acc_s3[1] ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.s1.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.s1.xor2_0._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.s1.xor2_0._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.s1.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.s1.xor2_1._1_  (.A1(\mult_u0.step4.add_sub4_u0.ppa8_u0.s1.temp ),
    .A2(\mult_u0.step4.add_sub4_u0.ppa8_u0.cg[0] ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.s1.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.s1.xor2_1._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.s1.xor2_1._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.S[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.s2.xor2_0._1_  (.A1(\mult_u0.step4.add_sub4_u0.int_ip[2] ),
    .A2(\mult_u0.acc_s3[2] ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.s2.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.s2.xor2_0._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.s2.xor2_0._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.s2.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.s2.xor2_1._1_  (.A1(\mult_u0.step4.add_sub4_u0.ppa8_u0.s2.temp ),
    .A2(\mult_u0.step4.add_sub4_u0.ppa8_u0.cg[1] ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.s2.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.s2.xor2_1._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.s2.xor2_1._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.S[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.s3.xor2_0._1_  (.A1(\mult_u0.step4.add_sub4_u0.int_ip[3] ),
    .A2(\mult_u0.acc_s3[3] ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.s3.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.s3.xor2_0._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.s3.xor2_0._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.s3.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.s3.xor2_1._1_  (.A1(\mult_u0.step4.add_sub4_u0.ppa8_u0.s3.temp ),
    .A2(\mult_u0.step4.add_sub4_u0.ppa8_u0.cg[2] ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.s3.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.s3.xor2_1._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.s3.xor2_1._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.S[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.s4.xor2_0._1_  (.A1(\mult_u0.step4.add_sub4_u0.int_ip[4] ),
    .A2(\mult_u0.acc_s3[4] ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.s4.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.s4.xor2_0._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.s4.xor2_0._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.s4.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.s4.xor2_1._1_  (.A1(\mult_u0.step4.add_sub4_u0.ppa8_u0.s4.temp ),
    .A2(\mult_u0.step4.add_sub4_u0.ppa8_u0.cg[3] ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.s4.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.s4.xor2_1._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.s4.xor2_1._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.S[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.s5.xor2_0._1_  (.A1(\mult_u0.step4.add_sub4_u0.int_ip[5] ),
    .A2(\mult_u0.acc_s3[5] ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.s5.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.s5.xor2_0._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.s5.xor2_0._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.s5.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.s5.xor2_1._1_  (.A1(\mult_u0.step4.add_sub4_u0.ppa8_u0.s5.temp ),
    .A2(\mult_u0.step4.add_sub4_u0.ppa8_u0.cg[4] ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.s5.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.s5.xor2_1._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.s5.xor2_1._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.S[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.s6.xor2_0._1_  (.A1(\mult_u0.step4.add_sub4_u0.int_ip[6] ),
    .A2(\mult_u0.acc_s3[6] ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.s6.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.s6.xor2_0._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.s6.xor2_0._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.s6.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.s6.xor2_1._1_  (.A1(\mult_u0.step4.add_sub4_u0.ppa8_u0.s6.temp ),
    .A2(\mult_u0.step4.add_sub4_u0.ppa8_u0.cg[5] ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.s6.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.ppa8_u0.s6.xor2_1._2_  (.I(\mult_u0.step4.add_sub4_u0.ppa8_u0.s6.xor2_1._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.ppa8_u0.S[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step4.add_sub4_u0.x0._1_  (.A1(\mult_u0.Q_s3[0] ),
    .A2(\mult_u0.multiplicand_s3[0] ),
    .Z(\mult_u0.step4.add_sub4_u0.x0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.x0._2_  (.I(\mult_u0.step4.add_sub4_u0.x0._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.int_ip[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step4.add_sub4_u0.x1._1_  (.A1(\mult_u0.Q_s3[0] ),
    .A2(\mult_u0.multiplicand_s3[1] ),
    .Z(\mult_u0.step4.add_sub4_u0.x1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.x1._2_  (.I(\mult_u0.step4.add_sub4_u0.x1._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.int_ip[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step4.add_sub4_u0.x2._1_  (.A1(\mult_u0.Q_s3[0] ),
    .A2(\mult_u0.multiplicand_s3[2] ),
    .Z(\mult_u0.step4.add_sub4_u0.x2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.x2._2_  (.I(\mult_u0.step4.add_sub4_u0.x2._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.int_ip[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step4.add_sub4_u0.x3._1_  (.A1(\mult_u0.Q_s3[0] ),
    .A2(\mult_u0.multiplicand_s3[3] ),
    .Z(\mult_u0.step4.add_sub4_u0.x3._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.x3._2_  (.I(\mult_u0.step4.add_sub4_u0.x3._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.int_ip[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step4.add_sub4_u0.x4._1_  (.A1(\mult_u0.Q_s3[0] ),
    .A2(\mult_u0.multiplicand_s3[4] ),
    .Z(\mult_u0.step4.add_sub4_u0.x4._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.x4._2_  (.I(\mult_u0.step4.add_sub4_u0.x4._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.int_ip[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step4.add_sub4_u0.x5._1_  (.A1(\mult_u0.Q_s3[0] ),
    .A2(\mult_u0.multiplicand_s3[5] ),
    .Z(\mult_u0.step4.add_sub4_u0.x5._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.x5._2_  (.I(\mult_u0.step4.add_sub4_u0.x5._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.int_ip[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step4.add_sub4_u0.x6._1_  (.A1(\mult_u0.Q_s3[0] ),
    .A2(\mult_u0.multiplicand_s3[6] ),
    .Z(\mult_u0.step4.add_sub4_u0.x6._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step4.add_sub4_u0.x6._2_  (.I(\mult_u0.step4.add_sub4_u0.x6._0_ ),
    .Z(\mult_u0.step4.add_sub4_u0.int_ip[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step5._09_  (.A1(\mult_u0.q0_s4 ),
    .A2(\mult_u0.Q_s4[0] ),
    .Z(\mult_u0.step5._00_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 \mult_u0.step5._10_  (.I(\mult_u0.step5._00_ ),
    .Z(\mult_u0.step5._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_u0.step5._13_  (.I0(\mult_u0.acc_s4[1] ),
    .I1(\mult_u0.step5.add_sub4_u0.ppa8_u0.S[1] ),
    .S(\mult_u0.step5._01_ ),
    .Z(\mult_u0.step5._03_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5._14_  (.I(\mult_u0.step5._03_ ),
    .Z(\mult_u0.acc[5][0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_u0.step5._15_  (.I0(\mult_u0.acc_s4[2] ),
    .I1(\mult_u0.step5.add_sub4_u0.ppa8_u0.S[2] ),
    .S(\mult_u0.step5._01_ ),
    .Z(\mult_u0.step5._04_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5._16_  (.I(\mult_u0.step5._04_ ),
    .Z(\mult_u0.acc[5][1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_u0.step5._17_  (.I0(\mult_u0.acc_s4[3] ),
    .I1(\mult_u0.step5.add_sub4_u0.ppa8_u0.S[3] ),
    .S(\mult_u0.step5._01_ ),
    .Z(\mult_u0.step5._05_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5._18_  (.I(\mult_u0.step5._05_ ),
    .Z(\mult_u0.acc[5][2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_u0.step5._19_  (.I0(\mult_u0.acc_s4[4] ),
    .I1(\mult_u0.step5.add_sub4_u0.ppa8_u0.S[4] ),
    .S(\mult_u0.step5._01_ ),
    .Z(\mult_u0.step5._06_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5._20_  (.I(\mult_u0.step5._06_ ),
    .Z(\mult_u0.acc[5][3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_u0.step5._21_  (.I0(\mult_u0.acc_s4[5] ),
    .I1(\mult_u0.step5.add_sub4_u0.ppa8_u0.S[5] ),
    .S(\mult_u0.step5._01_ ),
    .Z(\mult_u0.step5._07_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5._22_  (.I(\mult_u0.step5._07_ ),
    .Z(\mult_u0.acc[5][4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_u0.step5._23_  (.I0(\mult_u0.acc_s4[0] ),
    .I1(\mult_u0.step5.add_sub4_u0.ppa8_u0.S[0] ),
    .S(\mult_u0.step5._01_ ),
    .Z(\mult_u0.step5._08_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5._24_  (.I(\mult_u0.step5._08_ ),
    .Z(\mult_u0.Q[4][6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5._25_  (.I(\mult_u0.Q_s4[1] ),
    .Z(\mult_u0.Q[4][0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5._26_  (.I(\mult_u0.Q_s4[2] ),
    .Z(\mult_u0.Q[4][1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5._30_  (.I(\mult_u0.Q_s4[6] ),
    .Z(\mult_u0.Q[4][5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5._32_  (.I(\mult_u0.Q_s4[0] ),
    .Z(\mult_u0.q0[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.d1_0.a2._1_  (.A1(\mult_u0.Q_s4[0] ),
    .A2(\mult_u0.step5.add_sub4_u0.ppa8_u0.d1_0.a2.in0 ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.d1_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.d1_0.a2._2_  (.I(\mult_u0.step5.add_sub4_u0.ppa8_u0.d1_0.a2._0_ ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.d1_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.d1_0.o2._1_  (.A1(\mult_u0.step5.add_sub4_u0.ppa8_u0.d1_0.g1 ),
    .A2(\mult_u0.step5.add_sub4_u0.ppa8_u0.d1_0.a2.out ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.d1_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.d1_0.o2._2_  (.I(\mult_u0.step5.add_sub4_u0.ppa8_u0.d1_0.o2._0_ ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.cg[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.d2_0.a2._1_  (.A1(\mult_u0.step5.add_sub4_u0.ppa8_u0.cg[0] ),
    .A2(\mult_u0.step5.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.d2_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.d2_0.a2._2_  (.I(\mult_u0.step5.add_sub4_u0.ppa8_u0.d2_0.a2._0_ ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.d2_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.d2_0.o2._1_  (.A1(\mult_u0.step5.add_sub4_u0.ppa8_u0.d2_0.g1 ),
    .A2(\mult_u0.step5.add_sub4_u0.ppa8_u0.d2_0.a2.out ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.d2_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.d2_0.o2._2_  (.I(\mult_u0.step5.add_sub4_u0.ppa8_u0.d2_0.o2._0_ ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.cg[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.d3_0.a1._1_  (.A1(\mult_u0.step5.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ),
    .A2(\mult_u0.step5.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.d3_0.a1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.d3_0.a1._2_  (.I(\mult_u0.step5.add_sub4_u0.ppa8_u0.d3_0.a1._0_ ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.cp21 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.d3_0.a2._1_  (.A1(\mult_u0.step5.add_sub4_u0.ppa8_u0.d2_0.g1 ),
    .A2(\mult_u0.step5.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.d3_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.d3_0.a2._2_  (.I(\mult_u0.step5.add_sub4_u0.ppa8_u0.d3_0.a2._0_ ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.d3_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.d3_0.o2._1_  (.A1(\mult_u0.step5.add_sub4_u0.ppa8_u0.d3_0.g1 ),
    .A2(\mult_u0.step5.add_sub4_u0.ppa8_u0.d3_0.a2.out ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.d3_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.d3_0.o2._2_  (.I(\mult_u0.step5.add_sub4_u0.ppa8_u0.d3_0.o2._0_ ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.cg21 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.d3_1.a2._1_  (.A1(\mult_u0.step5.add_sub4_u0.ppa8_u0.cg[0] ),
    .A2(\mult_u0.step5.add_sub4_u0.ppa8_u0.cp21 ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.d3_1.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.d3_1.a2._2_  (.I(\mult_u0.step5.add_sub4_u0.ppa8_u0.d3_1.a2._0_ ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.d3_1.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.d3_1.o2._1_  (.A1(\mult_u0.step5.add_sub4_u0.ppa8_u0.cg21 ),
    .A2(\mult_u0.step5.add_sub4_u0.ppa8_u0.d3_1.a2.out ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.d3_1.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.d3_1.o2._2_  (.I(\mult_u0.step5.add_sub4_u0.ppa8_u0.d3_1.o2._0_ ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.cg[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.d4_0.a2._1_  (.A1(\mult_u0.step5.add_sub4_u0.ppa8_u0.cg[2] ),
    .A2(\mult_u0.step5.add_sub4_u0.ppa8_u0.d4_0.a2.in0 ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.d4_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.d4_0.a2._2_  (.I(\mult_u0.step5.add_sub4_u0.ppa8_u0.d4_0.a2._0_ ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.d4_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.d4_0.o2._1_  (.A1(\mult_u0.step5.add_sub4_u0.ppa8_u0.d4_0.g1 ),
    .A2(\mult_u0.step5.add_sub4_u0.ppa8_u0.d4_0.a2.out ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.d4_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.d4_0.o2._2_  (.I(\mult_u0.step5.add_sub4_u0.ppa8_u0.d4_0.o2._0_ ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.cg[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.d5_0.a1._1_  (.A1(\mult_u0.step5.add_sub4_u0.ppa8_u0.d4_0.a2.in0 ),
    .A2(\mult_u0.step5.add_sub4_u0.ppa8_u0.d5_0.a1.in0 ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.d5_0.a1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.d5_0.a1._2_  (.I(\mult_u0.step5.add_sub4_u0.ppa8_u0.d5_0.a1._0_ ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.cp43 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.d5_0.a2._1_  (.A1(\mult_u0.step5.add_sub4_u0.ppa8_u0.d4_0.g1 ),
    .A2(\mult_u0.step5.add_sub4_u0.ppa8_u0.d5_0.a1.in0 ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.d5_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.d5_0.a2._2_  (.I(\mult_u0.step5.add_sub4_u0.ppa8_u0.d5_0.a2._0_ ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.d5_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.d5_0.o2._1_  (.A1(\mult_u0.step5.add_sub4_u0.ppa8_u0.d5_0.g1 ),
    .A2(\mult_u0.step5.add_sub4_u0.ppa8_u0.d5_0.a2.out ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.d5_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.d5_0.o2._2_  (.I(\mult_u0.step5.add_sub4_u0.ppa8_u0.d5_0.o2._0_ ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.cg43 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.d5_1.a2._1_  (.A1(\mult_u0.step5.add_sub4_u0.ppa8_u0.cg[2] ),
    .A2(\mult_u0.step5.add_sub4_u0.ppa8_u0.cp43 ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.d5_1.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.d5_1.a2._2_  (.I(\mult_u0.step5.add_sub4_u0.ppa8_u0.d5_1.a2._0_ ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.d5_1.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.d5_1.o2._1_  (.A1(\mult_u0.step5.add_sub4_u0.ppa8_u0.cg43 ),
    .A2(\mult_u0.step5.add_sub4_u0.ppa8_u0.d5_1.a2.out ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.d5_1.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.d5_1.o2._2_  (.I(\mult_u0.step5.add_sub4_u0.ppa8_u0.d5_1.o2._0_ ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.cg[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.p_0.a._1_  (.A1(\mult_u0.step5.add_sub4_u0.int_ip[0] ),
    .A2(\mult_u0.acc_s4[0] ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.p_0.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.p_0.a._2_  (.I(\mult_u0.step5.add_sub4_u0.ppa8_u0.p_0.a._0_ ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.d1_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.p_0.o._1_  (.A1(\mult_u0.step5.add_sub4_u0.int_ip[0] ),
    .A2(\mult_u0.acc_s4[0] ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.p_0.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.p_0.o._2_  (.I(\mult_u0.step5.add_sub4_u0.ppa8_u0.p_0.o._0_ ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.d1_0.a2.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.p_1.a._1_  (.A1(\mult_u0.step5.add_sub4_u0.int_ip[1] ),
    .A2(\mult_u0.acc_s4[1] ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.p_1.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.p_1.a._2_  (.I(\mult_u0.step5.add_sub4_u0.ppa8_u0.p_1.a._0_ ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.d2_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.p_1.o._1_  (.A1(\mult_u0.step5.add_sub4_u0.int_ip[1] ),
    .A2(\mult_u0.acc_s4[1] ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.p_1.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.p_1.o._2_  (.I(\mult_u0.step5.add_sub4_u0.ppa8_u0.p_1.o._0_ ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.p_2.a._1_  (.A1(\mult_u0.step5.add_sub4_u0.int_ip[2] ),
    .A2(\mult_u0.acc_s4[2] ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.p_2.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.p_2.a._2_  (.I(\mult_u0.step5.add_sub4_u0.ppa8_u0.p_2.a._0_ ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.d3_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.p_2.o._1_  (.A1(\mult_u0.step5.add_sub4_u0.int_ip[2] ),
    .A2(\mult_u0.acc_s4[2] ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.p_2.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.p_2.o._2_  (.I(\mult_u0.step5.add_sub4_u0.ppa8_u0.p_2.o._0_ ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.p_3.a._1_  (.A1(\mult_u0.step5.add_sub4_u0.int_ip[3] ),
    .A2(\mult_u0.acc_s4[3] ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.p_3.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.p_3.a._2_  (.I(\mult_u0.step5.add_sub4_u0.ppa8_u0.p_3.a._0_ ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.d4_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.p_3.o._1_  (.A1(\mult_u0.step5.add_sub4_u0.int_ip[3] ),
    .A2(\mult_u0.acc_s4[3] ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.p_3.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.p_3.o._2_  (.I(\mult_u0.step5.add_sub4_u0.ppa8_u0.p_3.o._0_ ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.d4_0.a2.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.p_4.a._1_  (.A1(\mult_u0.step5.add_sub4_u0.int_ip[4] ),
    .A2(\mult_u0.acc_s4[4] ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.p_4.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.p_4.a._2_  (.I(\mult_u0.step5.add_sub4_u0.ppa8_u0.p_4.a._0_ ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.d5_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.p_4.o._1_  (.A1(\mult_u0.step5.add_sub4_u0.int_ip[4] ),
    .A2(\mult_u0.acc_s4[4] ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.p_4.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.p_4.o._2_  (.I(\mult_u0.step5.add_sub4_u0.ppa8_u0.p_4.o._0_ ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.d5_0.a1.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.s0.xor2_0._1_  (.A1(\mult_u0.step5.add_sub4_u0.int_ip[0] ),
    .A2(\mult_u0.acc_s4[0] ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.s0.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.s0.xor2_0._2_  (.I(\mult_u0.step5.add_sub4_u0.ppa8_u0.s0.xor2_0._0_ ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.s0.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.s0.xor2_1._1_  (.A1(\mult_u0.step5.add_sub4_u0.ppa8_u0.s0.temp ),
    .A2(\mult_u0.Q_s4[0] ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.s0.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.s0.xor2_1._2_  (.I(\mult_u0.step5.add_sub4_u0.ppa8_u0.s0.xor2_1._0_ ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.S[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.s1.xor2_0._1_  (.A1(\mult_u0.step5.add_sub4_u0.int_ip[1] ),
    .A2(\mult_u0.acc_s4[1] ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.s1.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.s1.xor2_0._2_  (.I(\mult_u0.step5.add_sub4_u0.ppa8_u0.s1.xor2_0._0_ ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.s1.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.s1.xor2_1._1_  (.A1(\mult_u0.step5.add_sub4_u0.ppa8_u0.s1.temp ),
    .A2(\mult_u0.step5.add_sub4_u0.ppa8_u0.cg[0] ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.s1.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.s1.xor2_1._2_  (.I(\mult_u0.step5.add_sub4_u0.ppa8_u0.s1.xor2_1._0_ ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.S[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.s2.xor2_0._1_  (.A1(\mult_u0.step5.add_sub4_u0.int_ip[2] ),
    .A2(\mult_u0.acc_s4[2] ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.s2.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.s2.xor2_0._2_  (.I(\mult_u0.step5.add_sub4_u0.ppa8_u0.s2.xor2_0._0_ ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.s2.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.s2.xor2_1._1_  (.A1(\mult_u0.step5.add_sub4_u0.ppa8_u0.s2.temp ),
    .A2(\mult_u0.step5.add_sub4_u0.ppa8_u0.cg[1] ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.s2.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.s2.xor2_1._2_  (.I(\mult_u0.step5.add_sub4_u0.ppa8_u0.s2.xor2_1._0_ ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.S[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.s3.xor2_0._1_  (.A1(\mult_u0.step5.add_sub4_u0.int_ip[3] ),
    .A2(\mult_u0.acc_s4[3] ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.s3.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.s3.xor2_0._2_  (.I(\mult_u0.step5.add_sub4_u0.ppa8_u0.s3.xor2_0._0_ ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.s3.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.s3.xor2_1._1_  (.A1(\mult_u0.step5.add_sub4_u0.ppa8_u0.s3.temp ),
    .A2(\mult_u0.step5.add_sub4_u0.ppa8_u0.cg[2] ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.s3.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.s3.xor2_1._2_  (.I(\mult_u0.step5.add_sub4_u0.ppa8_u0.s3.xor2_1._0_ ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.S[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.s4.xor2_0._1_  (.A1(\mult_u0.step5.add_sub4_u0.int_ip[4] ),
    .A2(\mult_u0.acc_s4[4] ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.s4.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.s4.xor2_0._2_  (.I(\mult_u0.step5.add_sub4_u0.ppa8_u0.s4.xor2_0._0_ ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.s4.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.s4.xor2_1._1_  (.A1(\mult_u0.step5.add_sub4_u0.ppa8_u0.s4.temp ),
    .A2(\mult_u0.step5.add_sub4_u0.ppa8_u0.cg[3] ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.s4.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.s4.xor2_1._2_  (.I(\mult_u0.step5.add_sub4_u0.ppa8_u0.s4.xor2_1._0_ ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.S[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.s5.xor2_0._1_  (.A1(\mult_u0.step5.add_sub4_u0.int_ip[5] ),
    .A2(\mult_u0.acc_s4[5] ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.s5.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.s5.xor2_0._2_  (.I(\mult_u0.step5.add_sub4_u0.ppa8_u0.s5.xor2_0._0_ ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.s5.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.s5.xor2_1._1_  (.A1(\mult_u0.step5.add_sub4_u0.ppa8_u0.s5.temp ),
    .A2(\mult_u0.step5.add_sub4_u0.ppa8_u0.cg[4] ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.s5.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5.add_sub4_u0.ppa8_u0.s5.xor2_1._2_  (.I(\mult_u0.step5.add_sub4_u0.ppa8_u0.s5.xor2_1._0_ ),
    .Z(\mult_u0.step5.add_sub4_u0.ppa8_u0.S[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step5.add_sub4_u0.x0._1_  (.A1(\mult_u0.Q_s4[0] ),
    .A2(\mult_u0.multiplicand_s4[0] ),
    .Z(\mult_u0.step5.add_sub4_u0.x0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5.add_sub4_u0.x0._2_  (.I(\mult_u0.step5.add_sub4_u0.x0._0_ ),
    .Z(\mult_u0.step5.add_sub4_u0.int_ip[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step5.add_sub4_u0.x1._1_  (.A1(\mult_u0.Q_s4[0] ),
    .A2(\mult_u0.multiplicand_s4[1] ),
    .Z(\mult_u0.step5.add_sub4_u0.x1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5.add_sub4_u0.x1._2_  (.I(\mult_u0.step5.add_sub4_u0.x1._0_ ),
    .Z(\mult_u0.step5.add_sub4_u0.int_ip[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step5.add_sub4_u0.x2._1_  (.A1(\mult_u0.Q_s4[0] ),
    .A2(\mult_u0.multiplicand_s4[2] ),
    .Z(\mult_u0.step5.add_sub4_u0.x2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5.add_sub4_u0.x2._2_  (.I(\mult_u0.step5.add_sub4_u0.x2._0_ ),
    .Z(\mult_u0.step5.add_sub4_u0.int_ip[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step5.add_sub4_u0.x3._1_  (.A1(\mult_u0.Q_s4[0] ),
    .A2(\mult_u0.multiplicand_s4[3] ),
    .Z(\mult_u0.step5.add_sub4_u0.x3._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5.add_sub4_u0.x3._2_  (.I(\mult_u0.step5.add_sub4_u0.x3._0_ ),
    .Z(\mult_u0.step5.add_sub4_u0.int_ip[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step5.add_sub4_u0.x4._1_  (.A1(\mult_u0.Q_s4[0] ),
    .A2(\mult_u0.multiplicand_s4[4] ),
    .Z(\mult_u0.step5.add_sub4_u0.x4._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5.add_sub4_u0.x4._2_  (.I(\mult_u0.step5.add_sub4_u0.x4._0_ ),
    .Z(\mult_u0.step5.add_sub4_u0.int_ip[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step5.add_sub4_u0.x5._1_  (.A1(\mult_u0.Q_s4[0] ),
    .A2(\mult_u0.multiplicand_s4[5] ),
    .Z(\mult_u0.step5.add_sub4_u0.x5._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step5.add_sub4_u0.x5._2_  (.I(\mult_u0.step5.add_sub4_u0.x5._0_ ),
    .Z(\mult_u0.step5.add_sub4_u0.int_ip[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step6._09_  (.A1(\mult_u0.q0_s5 ),
    .A2(\mult_u0.Q_s5[0] ),
    .Z(\mult_u0.step6._00_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 \mult_u0.step6._10_  (.I(\mult_u0.step6._00_ ),
    .Z(\mult_u0.step6._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_u0.step6._13_  (.I0(\mult_u0.acc_s5[1] ),
    .I1(\mult_u0.step6.add_sub4_u0.ppa8_u0.S[1] ),
    .S(\mult_u0.step6._01_ ),
    .Z(\mult_u0.step6._03_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step6._14_  (.I(\mult_u0.step6._03_ ),
    .Z(\mult_u0.acc[6][0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_u0.step6._15_  (.I0(\mult_u0.acc_s5[2] ),
    .I1(\mult_u0.step6.add_sub4_u0.ppa8_u0.S[2] ),
    .S(\mult_u0.step6._01_ ),
    .Z(\mult_u0.step6._04_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step6._16_  (.I(\mult_u0.step6._04_ ),
    .Z(\mult_u0.acc[6][1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_u0.step6._17_  (.I0(\mult_u0.acc_s5[3] ),
    .I1(\mult_u0.step6.add_sub4_u0.ppa8_u0.S[3] ),
    .S(\mult_u0.step6._01_ ),
    .Z(\mult_u0.step6._05_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step6._18_  (.I(\mult_u0.step6._05_ ),
    .Z(\mult_u0.acc[6][2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_u0.step6._19_  (.I0(\mult_u0.acc_s5[4] ),
    .I1(\mult_u0.step6.add_sub4_u0.ppa8_u0.S[4] ),
    .S(\mult_u0.step6._01_ ),
    .Z(\mult_u0.step6._06_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step6._20_  (.I(\mult_u0.step6._06_ ),
    .Z(\mult_u0.acc[6][3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_u0.step6._23_  (.I0(\mult_u0.acc_s5[0] ),
    .I1(\mult_u0.step6.add_sub4_u0.ppa8_u0.S[0] ),
    .S(\mult_u0.step6._01_ ),
    .Z(\mult_u0.step6._08_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step6._24_  (.I(\mult_u0.step6._08_ ),
    .Z(\mult_u0.Q[5][6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step6._25_  (.I(\mult_u0.Q_s5[1] ),
    .Z(\mult_u0.Q[5][0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step6._29_  (.I(\mult_u0.Q_s5[5] ),
    .Z(\mult_u0.Q[5][4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step6._30_  (.I(\mult_u0.Q_s5[6] ),
    .Z(\mult_u0.Q[5][5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step6._32_  (.I(\mult_u0.Q_s5[0] ),
    .Z(\mult_u0.q0[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.d1_0.a2._1_  (.A1(\mult_u0.Q_s5[0] ),
    .A2(\mult_u0.step6.add_sub4_u0.ppa8_u0.d1_0.a2.in0 ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.d1_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.d1_0.a2._2_  (.I(\mult_u0.step6.add_sub4_u0.ppa8_u0.d1_0.a2._0_ ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.d1_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.d1_0.o2._1_  (.A1(\mult_u0.step6.add_sub4_u0.ppa8_u0.d1_0.g1 ),
    .A2(\mult_u0.step6.add_sub4_u0.ppa8_u0.d1_0.a2.out ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.d1_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.d1_0.o2._2_  (.I(\mult_u0.step6.add_sub4_u0.ppa8_u0.d1_0.o2._0_ ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.cg[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.d2_0.a2._1_  (.A1(\mult_u0.step6.add_sub4_u0.ppa8_u0.cg[0] ),
    .A2(\mult_u0.step6.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.d2_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.d2_0.a2._2_  (.I(\mult_u0.step6.add_sub4_u0.ppa8_u0.d2_0.a2._0_ ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.d2_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.d2_0.o2._1_  (.A1(\mult_u0.step6.add_sub4_u0.ppa8_u0.d2_0.g1 ),
    .A2(\mult_u0.step6.add_sub4_u0.ppa8_u0.d2_0.a2.out ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.d2_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.d2_0.o2._2_  (.I(\mult_u0.step6.add_sub4_u0.ppa8_u0.d2_0.o2._0_ ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.cg[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.d3_0.a1._1_  (.A1(\mult_u0.step6.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ),
    .A2(\mult_u0.step6.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.d3_0.a1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.d3_0.a1._2_  (.I(\mult_u0.step6.add_sub4_u0.ppa8_u0.d3_0.a1._0_ ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.cp21 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.d3_0.a2._1_  (.A1(\mult_u0.step6.add_sub4_u0.ppa8_u0.d2_0.g1 ),
    .A2(\mult_u0.step6.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.d3_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.d3_0.a2._2_  (.I(\mult_u0.step6.add_sub4_u0.ppa8_u0.d3_0.a2._0_ ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.d3_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.d3_0.o2._1_  (.A1(\mult_u0.step6.add_sub4_u0.ppa8_u0.d3_0.g1 ),
    .A2(\mult_u0.step6.add_sub4_u0.ppa8_u0.d3_0.a2.out ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.d3_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.d3_0.o2._2_  (.I(\mult_u0.step6.add_sub4_u0.ppa8_u0.d3_0.o2._0_ ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.cg21 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.d3_1.a2._1_  (.A1(\mult_u0.step6.add_sub4_u0.ppa8_u0.cg[0] ),
    .A2(\mult_u0.step6.add_sub4_u0.ppa8_u0.cp21 ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.d3_1.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.d3_1.a2._2_  (.I(\mult_u0.step6.add_sub4_u0.ppa8_u0.d3_1.a2._0_ ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.d3_1.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.d3_1.o2._1_  (.A1(\mult_u0.step6.add_sub4_u0.ppa8_u0.cg21 ),
    .A2(\mult_u0.step6.add_sub4_u0.ppa8_u0.d3_1.a2.out ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.d3_1.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.d3_1.o2._2_  (.I(\mult_u0.step6.add_sub4_u0.ppa8_u0.d3_1.o2._0_ ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.cg[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.d4_0.a2._1_  (.A1(\mult_u0.step6.add_sub4_u0.ppa8_u0.cg[2] ),
    .A2(\mult_u0.step6.add_sub4_u0.ppa8_u0.d4_0.a2.in0 ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.d4_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.d4_0.a2._2_  (.I(\mult_u0.step6.add_sub4_u0.ppa8_u0.d4_0.a2._0_ ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.d4_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.d4_0.o2._1_  (.A1(\mult_u0.step6.add_sub4_u0.ppa8_u0.d4_0.g1 ),
    .A2(\mult_u0.step6.add_sub4_u0.ppa8_u0.d4_0.a2.out ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.d4_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.d4_0.o2._2_  (.I(\mult_u0.step6.add_sub4_u0.ppa8_u0.d4_0.o2._0_ ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.cg[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.p_0.a._1_  (.A1(\mult_u0.step6.add_sub4_u0.int_ip[0] ),
    .A2(\mult_u0.acc_s5[0] ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.p_0.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.p_0.a._2_  (.I(\mult_u0.step6.add_sub4_u0.ppa8_u0.p_0.a._0_ ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.d1_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.p_0.o._1_  (.A1(\mult_u0.step6.add_sub4_u0.int_ip[0] ),
    .A2(\mult_u0.acc_s5[0] ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.p_0.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.p_0.o._2_  (.I(\mult_u0.step6.add_sub4_u0.ppa8_u0.p_0.o._0_ ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.d1_0.a2.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.p_1.a._1_  (.A1(\mult_u0.step6.add_sub4_u0.int_ip[1] ),
    .A2(\mult_u0.acc_s5[1] ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.p_1.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.p_1.a._2_  (.I(\mult_u0.step6.add_sub4_u0.ppa8_u0.p_1.a._0_ ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.d2_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.p_1.o._1_  (.A1(\mult_u0.step6.add_sub4_u0.int_ip[1] ),
    .A2(\mult_u0.acc_s5[1] ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.p_1.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.p_1.o._2_  (.I(\mult_u0.step6.add_sub4_u0.ppa8_u0.p_1.o._0_ ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.p_2.a._1_  (.A1(\mult_u0.step6.add_sub4_u0.int_ip[2] ),
    .A2(\mult_u0.acc_s5[2] ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.p_2.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.p_2.a._2_  (.I(\mult_u0.step6.add_sub4_u0.ppa8_u0.p_2.a._0_ ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.d3_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.p_2.o._1_  (.A1(\mult_u0.step6.add_sub4_u0.int_ip[2] ),
    .A2(\mult_u0.acc_s5[2] ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.p_2.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.p_2.o._2_  (.I(\mult_u0.step6.add_sub4_u0.ppa8_u0.p_2.o._0_ ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.p_3.a._1_  (.A1(\mult_u0.step6.add_sub4_u0.int_ip[3] ),
    .A2(\mult_u0.acc_s5[3] ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.p_3.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.p_3.a._2_  (.I(\mult_u0.step6.add_sub4_u0.ppa8_u0.p_3.a._0_ ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.d4_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.p_3.o._1_  (.A1(\mult_u0.step6.add_sub4_u0.int_ip[3] ),
    .A2(\mult_u0.acc_s5[3] ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.p_3.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.p_3.o._2_  (.I(\mult_u0.step6.add_sub4_u0.ppa8_u0.p_3.o._0_ ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.d4_0.a2.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.s0.xor2_0._1_  (.A1(\mult_u0.step6.add_sub4_u0.int_ip[0] ),
    .A2(\mult_u0.acc_s5[0] ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.s0.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.s0.xor2_0._2_  (.I(\mult_u0.step6.add_sub4_u0.ppa8_u0.s0.xor2_0._0_ ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.s0.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.s0.xor2_1._1_  (.A1(\mult_u0.step6.add_sub4_u0.ppa8_u0.s0.temp ),
    .A2(\mult_u0.Q_s5[0] ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.s0.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.s0.xor2_1._2_  (.I(\mult_u0.step6.add_sub4_u0.ppa8_u0.s0.xor2_1._0_ ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.S[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.s1.xor2_0._1_  (.A1(\mult_u0.step6.add_sub4_u0.int_ip[1] ),
    .A2(\mult_u0.acc_s5[1] ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.s1.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.s1.xor2_0._2_  (.I(\mult_u0.step6.add_sub4_u0.ppa8_u0.s1.xor2_0._0_ ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.s1.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.s1.xor2_1._1_  (.A1(\mult_u0.step6.add_sub4_u0.ppa8_u0.s1.temp ),
    .A2(\mult_u0.step6.add_sub4_u0.ppa8_u0.cg[0] ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.s1.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.s1.xor2_1._2_  (.I(\mult_u0.step6.add_sub4_u0.ppa8_u0.s1.xor2_1._0_ ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.S[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.s2.xor2_0._1_  (.A1(\mult_u0.step6.add_sub4_u0.int_ip[2] ),
    .A2(\mult_u0.acc_s5[2] ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.s2.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.s2.xor2_0._2_  (.I(\mult_u0.step6.add_sub4_u0.ppa8_u0.s2.xor2_0._0_ ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.s2.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.s2.xor2_1._1_  (.A1(\mult_u0.step6.add_sub4_u0.ppa8_u0.s2.temp ),
    .A2(\mult_u0.step6.add_sub4_u0.ppa8_u0.cg[1] ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.s2.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.s2.xor2_1._2_  (.I(\mult_u0.step6.add_sub4_u0.ppa8_u0.s2.xor2_1._0_ ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.S[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.s3.xor2_0._1_  (.A1(\mult_u0.step6.add_sub4_u0.int_ip[3] ),
    .A2(\mult_u0.acc_s5[3] ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.s3.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.s3.xor2_0._2_  (.I(\mult_u0.step6.add_sub4_u0.ppa8_u0.s3.xor2_0._0_ ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.s3.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.s3.xor2_1._1_  (.A1(\mult_u0.step6.add_sub4_u0.ppa8_u0.s3.temp ),
    .A2(\mult_u0.step6.add_sub4_u0.ppa8_u0.cg[2] ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.s3.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.s3.xor2_1._2_  (.I(\mult_u0.step6.add_sub4_u0.ppa8_u0.s3.xor2_1._0_ ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.S[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.s4.xor2_0._1_  (.A1(\mult_u0.step6.add_sub4_u0.int_ip[4] ),
    .A2(\mult_u0.acc_s5[4] ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.s4.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.s4.xor2_0._2_  (.I(\mult_u0.step6.add_sub4_u0.ppa8_u0.s4.xor2_0._0_ ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.s4.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.s4.xor2_1._1_  (.A1(\mult_u0.step6.add_sub4_u0.ppa8_u0.s4.temp ),
    .A2(\mult_u0.step6.add_sub4_u0.ppa8_u0.cg[3] ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.s4.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step6.add_sub4_u0.ppa8_u0.s4.xor2_1._2_  (.I(\mult_u0.step6.add_sub4_u0.ppa8_u0.s4.xor2_1._0_ ),
    .Z(\mult_u0.step6.add_sub4_u0.ppa8_u0.S[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step6.add_sub4_u0.x0._1_  (.A1(\mult_u0.Q_s5[0] ),
    .A2(\mult_u0.multiplicand_s5[0] ),
    .Z(\mult_u0.step6.add_sub4_u0.x0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step6.add_sub4_u0.x0._2_  (.I(\mult_u0.step6.add_sub4_u0.x0._0_ ),
    .Z(\mult_u0.step6.add_sub4_u0.int_ip[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step6.add_sub4_u0.x1._1_  (.A1(\mult_u0.Q_s5[0] ),
    .A2(\mult_u0.multiplicand_s5[1] ),
    .Z(\mult_u0.step6.add_sub4_u0.x1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step6.add_sub4_u0.x1._2_  (.I(\mult_u0.step6.add_sub4_u0.x1._0_ ),
    .Z(\mult_u0.step6.add_sub4_u0.int_ip[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step6.add_sub4_u0.x2._1_  (.A1(\mult_u0.Q_s5[0] ),
    .A2(\mult_u0.multiplicand_s5[2] ),
    .Z(\mult_u0.step6.add_sub4_u0.x2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step6.add_sub4_u0.x2._2_  (.I(\mult_u0.step6.add_sub4_u0.x2._0_ ),
    .Z(\mult_u0.step6.add_sub4_u0.int_ip[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step6.add_sub4_u0.x3._1_  (.A1(\mult_u0.Q_s5[0] ),
    .A2(\mult_u0.multiplicand_s5[3] ),
    .Z(\mult_u0.step6.add_sub4_u0.x3._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step6.add_sub4_u0.x3._2_  (.I(\mult_u0.step6.add_sub4_u0.x3._0_ ),
    .Z(\mult_u0.step6.add_sub4_u0.int_ip[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step6.add_sub4_u0.x4._1_  (.A1(\mult_u0.Q_s5[0] ),
    .A2(\mult_u0.multiplicand_s5[4] ),
    .Z(\mult_u0.step6.add_sub4_u0.x4._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step6.add_sub4_u0.x4._2_  (.I(\mult_u0.step6.add_sub4_u0.x4._0_ ),
    .Z(\mult_u0.step6.add_sub4_u0.int_ip[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step7._09_  (.A1(\mult_u0.q0_s6 ),
    .A2(\mult_u0.Q_s6[0] ),
    .Z(\mult_u0.step7._00_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \mult_u0.step7._10_  (.I(\mult_u0.step7._00_ ),
    .Z(\mult_u0.step7._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_u0.step7._13_  (.I0(\mult_u0.acc_s6[1] ),
    .I1(\mult_u0.step7.add_sub4_u0.ppa8_u0.S[1] ),
    .S(\mult_u0.step7._01_ ),
    .Z(\mult_u0.step7._03_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step7._14_  (.I(\mult_u0.step7._03_ ),
    .Z(\mult_u0.step7.next_acc[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_u0.step7._15_  (.I0(\mult_u0.acc_s6[2] ),
    .I1(\mult_u0.step7.add_sub4_u0.ppa8_u0.S[2] ),
    .S(\mult_u0.step7._01_ ),
    .Z(\mult_u0.step7._04_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step7._16_  (.I(\mult_u0.step7._04_ ),
    .Z(\mult_u0.step7.next_acc[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_u0.step7._17_  (.I0(\mult_u0.acc_s6[3] ),
    .I1(\mult_u0.step7.add_sub4_u0.ppa8_u0.S[3] ),
    .S(\mult_u0.step7._01_ ),
    .Z(\mult_u0.step7._05_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step7._18_  (.I(\mult_u0.step7._05_ ),
    .Z(\mult_u0.step7.next_acc[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 \mult_u0.step7._23_  (.I0(\mult_u0.acc_s6[0] ),
    .I1(\mult_u0.step7.add_sub4_u0.ppa8_u0.S[0] ),
    .S(\mult_u0.step7._01_ ),
    .Z(\mult_u0.step7._08_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step7._24_  (.I(\mult_u0.step7._08_ ),
    .Z(\mult_u0.product[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step7._28_  (.I(\mult_u0.Q_s6[4] ),
    .Z(\mult_u0.product[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step7._29_  (.I(\mult_u0.Q_s6[5] ),
    .Z(\mult_u0.product[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step7._30_  (.I(\mult_u0.Q_s6[6] ),
    .Z(\mult_u0.product[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step7.add_sub4_u0.ppa8_u0.d1_0.a2._1_  (.A1(\mult_u0.Q_s6[0] ),
    .A2(\mult_u0.step7.add_sub4_u0.ppa8_u0.d1_0.a2.in0 ),
    .Z(\mult_u0.step7.add_sub4_u0.ppa8_u0.d1_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step7.add_sub4_u0.ppa8_u0.d1_0.a2._2_  (.I(\mult_u0.step7.add_sub4_u0.ppa8_u0.d1_0.a2._0_ ),
    .Z(\mult_u0.step7.add_sub4_u0.ppa8_u0.d1_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step7.add_sub4_u0.ppa8_u0.d1_0.o2._1_  (.A1(\mult_u0.step7.add_sub4_u0.ppa8_u0.d1_0.g1 ),
    .A2(\mult_u0.step7.add_sub4_u0.ppa8_u0.d1_0.a2.out ),
    .Z(\mult_u0.step7.add_sub4_u0.ppa8_u0.d1_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step7.add_sub4_u0.ppa8_u0.d1_0.o2._2_  (.I(\mult_u0.step7.add_sub4_u0.ppa8_u0.d1_0.o2._0_ ),
    .Z(\mult_u0.step7.add_sub4_u0.ppa8_u0.cg[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step7.add_sub4_u0.ppa8_u0.d2_0.a2._1_  (.A1(\mult_u0.step7.add_sub4_u0.ppa8_u0.cg[0] ),
    .A2(\mult_u0.step7.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ),
    .Z(\mult_u0.step7.add_sub4_u0.ppa8_u0.d2_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step7.add_sub4_u0.ppa8_u0.d2_0.a2._2_  (.I(\mult_u0.step7.add_sub4_u0.ppa8_u0.d2_0.a2._0_ ),
    .Z(\mult_u0.step7.add_sub4_u0.ppa8_u0.d2_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step7.add_sub4_u0.ppa8_u0.d2_0.o2._1_  (.A1(\mult_u0.step7.add_sub4_u0.ppa8_u0.d2_0.g1 ),
    .A2(\mult_u0.step7.add_sub4_u0.ppa8_u0.d2_0.a2.out ),
    .Z(\mult_u0.step7.add_sub4_u0.ppa8_u0.d2_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step7.add_sub4_u0.ppa8_u0.d2_0.o2._2_  (.I(\mult_u0.step7.add_sub4_u0.ppa8_u0.d2_0.o2._0_ ),
    .Z(\mult_u0.step7.add_sub4_u0.ppa8_u0.cg[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step7.add_sub4_u0.ppa8_u0.d3_0.a1._1_  (.A1(\mult_u0.step7.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ),
    .A2(\mult_u0.step7.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ),
    .Z(\mult_u0.step7.add_sub4_u0.ppa8_u0.d3_0.a1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step7.add_sub4_u0.ppa8_u0.d3_0.a1._2_  (.I(\mult_u0.step7.add_sub4_u0.ppa8_u0.d3_0.a1._0_ ),
    .Z(\mult_u0.step7.add_sub4_u0.ppa8_u0.cp21 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step7.add_sub4_u0.ppa8_u0.d3_0.a2._1_  (.A1(\mult_u0.step7.add_sub4_u0.ppa8_u0.d2_0.g1 ),
    .A2(\mult_u0.step7.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ),
    .Z(\mult_u0.step7.add_sub4_u0.ppa8_u0.d3_0.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step7.add_sub4_u0.ppa8_u0.d3_0.a2._2_  (.I(\mult_u0.step7.add_sub4_u0.ppa8_u0.d3_0.a2._0_ ),
    .Z(\mult_u0.step7.add_sub4_u0.ppa8_u0.d3_0.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step7.add_sub4_u0.ppa8_u0.d3_0.o2._1_  (.A1(\mult_u0.step7.add_sub4_u0.ppa8_u0.d3_0.g1 ),
    .A2(\mult_u0.step7.add_sub4_u0.ppa8_u0.d3_0.a2.out ),
    .Z(\mult_u0.step7.add_sub4_u0.ppa8_u0.d3_0.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step7.add_sub4_u0.ppa8_u0.d3_0.o2._2_  (.I(\mult_u0.step7.add_sub4_u0.ppa8_u0.d3_0.o2._0_ ),
    .Z(\mult_u0.step7.add_sub4_u0.ppa8_u0.cg21 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step7.add_sub4_u0.ppa8_u0.d3_1.a2._1_  (.A1(\mult_u0.step7.add_sub4_u0.ppa8_u0.cg[0] ),
    .A2(\mult_u0.step7.add_sub4_u0.ppa8_u0.cp21 ),
    .Z(\mult_u0.step7.add_sub4_u0.ppa8_u0.d3_1.a2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step7.add_sub4_u0.ppa8_u0.d3_1.a2._2_  (.I(\mult_u0.step7.add_sub4_u0.ppa8_u0.d3_1.a2._0_ ),
    .Z(\mult_u0.step7.add_sub4_u0.ppa8_u0.d3_1.a2.out ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step7.add_sub4_u0.ppa8_u0.d3_1.o2._1_  (.A1(\mult_u0.step7.add_sub4_u0.ppa8_u0.cg21 ),
    .A2(\mult_u0.step7.add_sub4_u0.ppa8_u0.d3_1.a2.out ),
    .Z(\mult_u0.step7.add_sub4_u0.ppa8_u0.d3_1.o2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step7.add_sub4_u0.ppa8_u0.d3_1.o2._2_  (.I(\mult_u0.step7.add_sub4_u0.ppa8_u0.d3_1.o2._0_ ),
    .Z(\mult_u0.step7.add_sub4_u0.ppa8_u0.cg[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step7.add_sub4_u0.ppa8_u0.p_0.a._1_  (.A1(\mult_u0.step7.add_sub4_u0.int_ip[0] ),
    .A2(\mult_u0.acc_s6[0] ),
    .Z(\mult_u0.step7.add_sub4_u0.ppa8_u0.p_0.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step7.add_sub4_u0.ppa8_u0.p_0.a._2_  (.I(\mult_u0.step7.add_sub4_u0.ppa8_u0.p_0.a._0_ ),
    .Z(\mult_u0.step7.add_sub4_u0.ppa8_u0.d1_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step7.add_sub4_u0.ppa8_u0.p_0.o._1_  (.A1(\mult_u0.step7.add_sub4_u0.int_ip[0] ),
    .A2(\mult_u0.acc_s6[0] ),
    .Z(\mult_u0.step7.add_sub4_u0.ppa8_u0.p_0.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step7.add_sub4_u0.ppa8_u0.p_0.o._2_  (.I(\mult_u0.step7.add_sub4_u0.ppa8_u0.p_0.o._0_ ),
    .Z(\mult_u0.step7.add_sub4_u0.ppa8_u0.d1_0.a2.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step7.add_sub4_u0.ppa8_u0.p_1.a._1_  (.A1(\mult_u0.step7.add_sub4_u0.int_ip[1] ),
    .A2(\mult_u0.acc_s6[1] ),
    .Z(\mult_u0.step7.add_sub4_u0.ppa8_u0.p_1.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step7.add_sub4_u0.ppa8_u0.p_1.a._2_  (.I(\mult_u0.step7.add_sub4_u0.ppa8_u0.p_1.a._0_ ),
    .Z(\mult_u0.step7.add_sub4_u0.ppa8_u0.d2_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step7.add_sub4_u0.ppa8_u0.p_1.o._1_  (.A1(\mult_u0.step7.add_sub4_u0.int_ip[1] ),
    .A2(\mult_u0.acc_s6[1] ),
    .Z(\mult_u0.step7.add_sub4_u0.ppa8_u0.p_1.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step7.add_sub4_u0.ppa8_u0.p_1.o._2_  (.I(\mult_u0.step7.add_sub4_u0.ppa8_u0.p_1.o._0_ ),
    .Z(\mult_u0.step7.add_sub4_u0.ppa8_u0.d2_0.a2.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \mult_u0.step7.add_sub4_u0.ppa8_u0.p_2.a._1_  (.A1(\mult_u0.step7.add_sub4_u0.int_ip[2] ),
    .A2(\mult_u0.acc_s6[2] ),
    .Z(\mult_u0.step7.add_sub4_u0.ppa8_u0.p_2.a._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step7.add_sub4_u0.ppa8_u0.p_2.a._2_  (.I(\mult_u0.step7.add_sub4_u0.ppa8_u0.p_2.a._0_ ),
    .Z(\mult_u0.step7.add_sub4_u0.ppa8_u0.d3_0.g1 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \mult_u0.step7.add_sub4_u0.ppa8_u0.p_2.o._1_  (.A1(\mult_u0.step7.add_sub4_u0.int_ip[2] ),
    .A2(\mult_u0.acc_s6[2] ),
    .Z(\mult_u0.step7.add_sub4_u0.ppa8_u0.p_2.o._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step7.add_sub4_u0.ppa8_u0.p_2.o._2_  (.I(\mult_u0.step7.add_sub4_u0.ppa8_u0.p_2.o._0_ ),
    .Z(\mult_u0.step7.add_sub4_u0.ppa8_u0.d3_0.a1.in0 ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step7.add_sub4_u0.ppa8_u0.s0.xor2_0._1_  (.A1(\mult_u0.step7.add_sub4_u0.int_ip[0] ),
    .A2(\mult_u0.acc_s6[0] ),
    .Z(\mult_u0.step7.add_sub4_u0.ppa8_u0.s0.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step7.add_sub4_u0.ppa8_u0.s0.xor2_0._2_  (.I(\mult_u0.step7.add_sub4_u0.ppa8_u0.s0.xor2_0._0_ ),
    .Z(\mult_u0.step7.add_sub4_u0.ppa8_u0.s0.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step7.add_sub4_u0.ppa8_u0.s0.xor2_1._1_  (.A1(\mult_u0.step7.add_sub4_u0.ppa8_u0.s0.temp ),
    .A2(\mult_u0.Q_s6[0] ),
    .Z(\mult_u0.step7.add_sub4_u0.ppa8_u0.s0.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step7.add_sub4_u0.ppa8_u0.s0.xor2_1._2_  (.I(\mult_u0.step7.add_sub4_u0.ppa8_u0.s0.xor2_1._0_ ),
    .Z(\mult_u0.step7.add_sub4_u0.ppa8_u0.S[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step7.add_sub4_u0.ppa8_u0.s1.xor2_0._1_  (.A1(\mult_u0.step7.add_sub4_u0.int_ip[1] ),
    .A2(\mult_u0.acc_s6[1] ),
    .Z(\mult_u0.step7.add_sub4_u0.ppa8_u0.s1.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step7.add_sub4_u0.ppa8_u0.s1.xor2_0._2_  (.I(\mult_u0.step7.add_sub4_u0.ppa8_u0.s1.xor2_0._0_ ),
    .Z(\mult_u0.step7.add_sub4_u0.ppa8_u0.s1.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step7.add_sub4_u0.ppa8_u0.s1.xor2_1._1_  (.A1(\mult_u0.step7.add_sub4_u0.ppa8_u0.s1.temp ),
    .A2(\mult_u0.step7.add_sub4_u0.ppa8_u0.cg[0] ),
    .Z(\mult_u0.step7.add_sub4_u0.ppa8_u0.s1.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step7.add_sub4_u0.ppa8_u0.s1.xor2_1._2_  (.I(\mult_u0.step7.add_sub4_u0.ppa8_u0.s1.xor2_1._0_ ),
    .Z(\mult_u0.step7.add_sub4_u0.ppa8_u0.S[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step7.add_sub4_u0.ppa8_u0.s2.xor2_0._1_  (.A1(\mult_u0.step7.add_sub4_u0.int_ip[2] ),
    .A2(\mult_u0.acc_s6[2] ),
    .Z(\mult_u0.step7.add_sub4_u0.ppa8_u0.s2.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step7.add_sub4_u0.ppa8_u0.s2.xor2_0._2_  (.I(\mult_u0.step7.add_sub4_u0.ppa8_u0.s2.xor2_0._0_ ),
    .Z(\mult_u0.step7.add_sub4_u0.ppa8_u0.s2.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step7.add_sub4_u0.ppa8_u0.s2.xor2_1._1_  (.A1(\mult_u0.step7.add_sub4_u0.ppa8_u0.s2.temp ),
    .A2(\mult_u0.step7.add_sub4_u0.ppa8_u0.cg[1] ),
    .Z(\mult_u0.step7.add_sub4_u0.ppa8_u0.s2.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step7.add_sub4_u0.ppa8_u0.s2.xor2_1._2_  (.I(\mult_u0.step7.add_sub4_u0.ppa8_u0.s2.xor2_1._0_ ),
    .Z(\mult_u0.step7.add_sub4_u0.ppa8_u0.S[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step7.add_sub4_u0.ppa8_u0.s3.xor2_0._1_  (.A1(\mult_u0.step7.add_sub4_u0.int_ip[3] ),
    .A2(\mult_u0.acc_s6[3] ),
    .Z(\mult_u0.step7.add_sub4_u0.ppa8_u0.s3.xor2_0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step7.add_sub4_u0.ppa8_u0.s3.xor2_0._2_  (.I(\mult_u0.step7.add_sub4_u0.ppa8_u0.s3.xor2_0._0_ ),
    .Z(\mult_u0.step7.add_sub4_u0.ppa8_u0.s3.temp ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step7.add_sub4_u0.ppa8_u0.s3.xor2_1._1_  (.A1(\mult_u0.step7.add_sub4_u0.ppa8_u0.s3.temp ),
    .A2(\mult_u0.step7.add_sub4_u0.ppa8_u0.cg[2] ),
    .Z(\mult_u0.step7.add_sub4_u0.ppa8_u0.s3.xor2_1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step7.add_sub4_u0.ppa8_u0.s3.xor2_1._2_  (.I(\mult_u0.step7.add_sub4_u0.ppa8_u0.s3.xor2_1._0_ ),
    .Z(\mult_u0.step7.add_sub4_u0.ppa8_u0.S[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step7.add_sub4_u0.x0._1_  (.A1(\mult_u0.Q_s6[0] ),
    .A2(\mult_u0.multiplicand_s6[0] ),
    .Z(\mult_u0.step7.add_sub4_u0.x0._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step7.add_sub4_u0.x0._2_  (.I(\mult_u0.step7.add_sub4_u0.x0._0_ ),
    .Z(\mult_u0.step7.add_sub4_u0.int_ip[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step7.add_sub4_u0.x1._1_  (.A1(\mult_u0.Q_s6[0] ),
    .A2(\mult_u0.multiplicand_s6[1] ),
    .Z(\mult_u0.step7.add_sub4_u0.x1._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step7.add_sub4_u0.x1._2_  (.I(\mult_u0.step7.add_sub4_u0.x1._0_ ),
    .Z(\mult_u0.step7.add_sub4_u0.int_ip[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step7.add_sub4_u0.x2._1_  (.A1(\mult_u0.Q_s6[0] ),
    .A2(\mult_u0.multiplicand_s6[2] ),
    .Z(\mult_u0.step7.add_sub4_u0.x2._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step7.add_sub4_u0.x2._2_  (.I(\mult_u0.step7.add_sub4_u0.x2._0_ ),
    .Z(\mult_u0.step7.add_sub4_u0.int_ip[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.step7.add_sub4_u0.x3._1_  (.A1(\mult_u0.Q_s6[0] ),
    .A2(\mult_u0.multiplicand_s6[3] ),
    .Z(\mult_u0.step7.add_sub4_u0.x3._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.step7.add_sub4_u0.x3._2_  (.I(\mult_u0.step7.add_sub4_u0.x3._0_ ),
    .Z(\mult_u0.step7.add_sub4_u0.int_ip[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \mult_u0.x_sign._1_  (.A1(\add_u0.b[7] ),
    .A2(\add_u0.a[7] ),
    .Z(\mult_u0.x_sign._0_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \mult_u0.x_sign._2_  (.I(\mult_u0.x_sign._0_ ),
    .Z(\mult_u0.mul_sign ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 wire1 (.I(clk),
    .Z(net114),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 assign o_wb_stall = net63;
endmodule
