VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO uart_i2c_usb_spi_top
  CLASS BLOCK ;
  FOREIGN uart_i2c_usb_spi_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 1000.000 BY 900.000 ;
  PIN app_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 973.280 0.000 973.840 4.000 ;
    END
  END app_clk
  PIN i2c_rstn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 209.440 896.000 210.000 900.000 ;
    END
  END i2c_rstn
  PIN i2cm_intr_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 473.760 1000.000 474.320 ;
    END
  END i2cm_intr_o
  PIN reg_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 879.200 4.000 879.760 ;
    END
  END reg_ack
  PIN reg_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 227.360 0.000 227.920 4.000 ;
    END
  END reg_addr[0]
  PIN reg_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 207.200 0.000 207.760 4.000 ;
    END
  END reg_addr[1]
  PIN reg_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 187.040 0.000 187.600 4.000 ;
    END
  END reg_addr[2]
  PIN reg_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 166.880 0.000 167.440 4.000 ;
    END
  END reg_addr[3]
  PIN reg_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 146.720 0.000 147.280 4.000 ;
    END
  END reg_addr[4]
  PIN reg_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 126.560 0.000 127.120 4.000 ;
    END
  END reg_addr[5]
  PIN reg_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 106.400 0.000 106.960 4.000 ;
    END
  END reg_addr[6]
  PIN reg_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 86.240 0.000 86.800 4.000 ;
    END
  END reg_addr[7]
  PIN reg_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 66.080 0.000 66.640 4.000 ;
    END
  END reg_addr[8]
  PIN reg_be[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 308.000 0.000 308.560 4.000 ;
    END
  END reg_be[0]
  PIN reg_be[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 287.840 0.000 288.400 4.000 ;
    END
  END reg_be[1]
  PIN reg_be[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 267.680 0.000 268.240 4.000 ;
    END
  END reg_be[2]
  PIN reg_be[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 247.520 0.000 248.080 4.000 ;
    END
  END reg_be[3]
  PIN reg_cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 25.760 0.000 26.320 4.000 ;
    END
  END reg_cs
  PIN reg_rdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 852.320 4.000 852.880 ;
    END
  END reg_rdata[0]
  PIN reg_rdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 583.520 4.000 584.080 ;
    END
  END reg_rdata[10]
  PIN reg_rdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 556.640 4.000 557.200 ;
    END
  END reg_rdata[11]
  PIN reg_rdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 529.760 4.000 530.320 ;
    END
  END reg_rdata[12]
  PIN reg_rdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 502.880 4.000 503.440 ;
    END
  END reg_rdata[13]
  PIN reg_rdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 476.000 4.000 476.560 ;
    END
  END reg_rdata[14]
  PIN reg_rdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 449.120 4.000 449.680 ;
    END
  END reg_rdata[15]
  PIN reg_rdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 422.240 4.000 422.800 ;
    END
  END reg_rdata[16]
  PIN reg_rdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 395.360 4.000 395.920 ;
    END
  END reg_rdata[17]
  PIN reg_rdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 368.480 4.000 369.040 ;
    END
  END reg_rdata[18]
  PIN reg_rdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 341.600 4.000 342.160 ;
    END
  END reg_rdata[19]
  PIN reg_rdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 825.440 4.000 826.000 ;
    END
  END reg_rdata[1]
  PIN reg_rdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 314.720 4.000 315.280 ;
    END
  END reg_rdata[20]
  PIN reg_rdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 287.840 4.000 288.400 ;
    END
  END reg_rdata[21]
  PIN reg_rdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 260.960 4.000 261.520 ;
    END
  END reg_rdata[22]
  PIN reg_rdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 234.080 4.000 234.640 ;
    END
  END reg_rdata[23]
  PIN reg_rdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 207.200 4.000 207.760 ;
    END
  END reg_rdata[24]
  PIN reg_rdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 180.320 4.000 180.880 ;
    END
  END reg_rdata[25]
  PIN reg_rdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 153.440 4.000 154.000 ;
    END
  END reg_rdata[26]
  PIN reg_rdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 126.560 4.000 127.120 ;
    END
  END reg_rdata[27]
  PIN reg_rdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 99.680 4.000 100.240 ;
    END
  END reg_rdata[28]
  PIN reg_rdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 72.800 4.000 73.360 ;
    END
  END reg_rdata[29]
  PIN reg_rdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 798.560 4.000 799.120 ;
    END
  END reg_rdata[2]
  PIN reg_rdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 45.920 4.000 46.480 ;
    END
  END reg_rdata[30]
  PIN reg_rdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 19.040 4.000 19.600 ;
    END
  END reg_rdata[31]
  PIN reg_rdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 771.680 4.000 772.240 ;
    END
  END reg_rdata[3]
  PIN reg_rdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 744.800 4.000 745.360 ;
    END
  END reg_rdata[4]
  PIN reg_rdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 717.920 4.000 718.480 ;
    END
  END reg_rdata[5]
  PIN reg_rdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 691.040 4.000 691.600 ;
    END
  END reg_rdata[6]
  PIN reg_rdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 664.160 4.000 664.720 ;
    END
  END reg_rdata[7]
  PIN reg_rdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 637.280 4.000 637.840 ;
    END
  END reg_rdata[8]
  PIN reg_rdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 610.400 4.000 610.960 ;
    END
  END reg_rdata[9]
  PIN reg_wdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 953.120 0.000 953.680 4.000 ;
    END
  END reg_wdata[0]
  PIN reg_wdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 751.520 0.000 752.080 4.000 ;
    END
  END reg_wdata[10]
  PIN reg_wdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 731.360 0.000 731.920 4.000 ;
    END
  END reg_wdata[11]
  PIN reg_wdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 711.200 0.000 711.760 4.000 ;
    END
  END reg_wdata[12]
  PIN reg_wdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 691.040 0.000 691.600 4.000 ;
    END
  END reg_wdata[13]
  PIN reg_wdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 670.880 0.000 671.440 4.000 ;
    END
  END reg_wdata[14]
  PIN reg_wdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 650.720 0.000 651.280 4.000 ;
    END
  END reg_wdata[15]
  PIN reg_wdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 630.560 0.000 631.120 4.000 ;
    END
  END reg_wdata[16]
  PIN reg_wdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 610.400 0.000 610.960 4.000 ;
    END
  END reg_wdata[17]
  PIN reg_wdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 590.240 0.000 590.800 4.000 ;
    END
  END reg_wdata[18]
  PIN reg_wdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 570.080 0.000 570.640 4.000 ;
    END
  END reg_wdata[19]
  PIN reg_wdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 932.960 0.000 933.520 4.000 ;
    END
  END reg_wdata[1]
  PIN reg_wdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 549.920 0.000 550.480 4.000 ;
    END
  END reg_wdata[20]
  PIN reg_wdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 529.760 0.000 530.320 4.000 ;
    END
  END reg_wdata[21]
  PIN reg_wdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 509.600 0.000 510.160 4.000 ;
    END
  END reg_wdata[22]
  PIN reg_wdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 489.440 0.000 490.000 4.000 ;
    END
  END reg_wdata[23]
  PIN reg_wdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 469.280 0.000 469.840 4.000 ;
    END
  END reg_wdata[24]
  PIN reg_wdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 449.120 0.000 449.680 4.000 ;
    END
  END reg_wdata[25]
  PIN reg_wdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 428.960 0.000 429.520 4.000 ;
    END
  END reg_wdata[26]
  PIN reg_wdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 408.800 0.000 409.360 4.000 ;
    END
  END reg_wdata[27]
  PIN reg_wdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 388.640 0.000 389.200 4.000 ;
    END
  END reg_wdata[28]
  PIN reg_wdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 368.480 0.000 369.040 4.000 ;
    END
  END reg_wdata[29]
  PIN reg_wdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 912.800 0.000 913.360 4.000 ;
    END
  END reg_wdata[2]
  PIN reg_wdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 348.320 0.000 348.880 4.000 ;
    END
  END reg_wdata[30]
  PIN reg_wdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 328.160 0.000 328.720 4.000 ;
    END
  END reg_wdata[31]
  PIN reg_wdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 892.640 0.000 893.200 4.000 ;
    END
  END reg_wdata[3]
  PIN reg_wdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 872.480 0.000 873.040 4.000 ;
    END
  END reg_wdata[4]
  PIN reg_wdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 852.320 0.000 852.880 4.000 ;
    END
  END reg_wdata[5]
  PIN reg_wdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 832.160 0.000 832.720 4.000 ;
    END
  END reg_wdata[6]
  PIN reg_wdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 812.000 0.000 812.560 4.000 ;
    END
  END reg_wdata[7]
  PIN reg_wdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 791.840 0.000 792.400 4.000 ;
    END
  END reg_wdata[8]
  PIN reg_wdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 771.680 0.000 772.240 4.000 ;
    END
  END reg_wdata[9]
  PIN reg_wr
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 45.920 0.000 46.480 4.000 ;
    END
  END reg_wr
  PIN scl_pad_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 540.960 896.000 541.520 900.000 ;
    END
  END scl_pad_i
  PIN scl_pad_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 623.840 896.000 624.400 900.000 ;
    END
  END scl_pad_o
  PIN scl_pad_oen_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 706.720 896.000 707.280 900.000 ;
    END
  END scl_pad_oen_o
  PIN sda_pad_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 789.600 896.000 790.160 900.000 ;
    END
  END sda_pad_i
  PIN sda_pad_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 872.480 896.000 873.040 900.000 ;
    END
  END sda_pad_o
  PIN sda_padoen_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 955.360 896.000 955.920 900.000 ;
    END
  END sda_padoen_o
  PIN spi_rstn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 375.200 896.000 375.760 900.000 ;
    END
  END spi_rstn
  PIN sspim_sck
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 572.320 1000.000 572.880 ;
    END
  END sspim_sck
  PIN sspim_si
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 621.600 1000.000 622.160 ;
    END
  END sspim_si
  PIN sspim_so
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 670.880 1000.000 671.440 ;
    END
  END sspim_so
  PIN sspim_ssn[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 868.000 1000.000 868.560 ;
    END
  END sspim_ssn[0]
  PIN sspim_ssn[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 818.720 1000.000 819.280 ;
    END
  END sspim_ssn[1]
  PIN sspim_ssn[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 769.440 1000.000 770.000 ;
    END
  END sspim_ssn[2]
  PIN sspim_ssn[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 720.160 1000.000 720.720 ;
    END
  END sspim_ssn[3]
  PIN uart_rstn[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 126.560 896.000 127.120 900.000 ;
    END
  END uart_rstn[0]
  PIN uart_rstn[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 43.680 896.000 44.240 900.000 ;
    END
  END uart_rstn[1]
  PIN uart_rxd[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 30.240 1000.000 30.800 ;
    END
  END uart_rxd[0]
  PIN uart_rxd[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 128.800 1000.000 129.360 ;
    END
  END uart_rxd[1]
  PIN uart_txd[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 79.520 1000.000 80.080 ;
    END
  END uart_txd[0]
  PIN uart_txd[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 178.080 1000.000 178.640 ;
    END
  END uart_txd[1]
  PIN usb_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 458.080 896.000 458.640 900.000 ;
    END
  END usb_clk
  PIN usb_in_dn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 276.640 1000.000 277.200 ;
    END
  END usb_in_dn
  PIN usb_in_dp
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 227.360 1000.000 227.920 ;
    END
  END usb_in_dp
  PIN usb_intr_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 523.040 1000.000 523.600 ;
    END
  END usb_intr_o
  PIN usb_out_dn
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 375.200 1000.000 375.760 ;
    END
  END usb_out_dn
  PIN usb_out_dp
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 325.920 1000.000 326.480 ;
    END
  END usb_out_dp
  PIN usb_out_tx_oen
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 424.480 1000.000 425.040 ;
    END
  END usb_out_tx_oen
  PIN usb_rstn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 292.320 896.000 292.880 900.000 ;
    END
  END usb_rstn
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 19.940 15.380 26.140 882.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 119.940 15.380 126.140 882.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 219.940 15.380 226.140 882.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 319.940 15.380 326.140 882.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 419.940 15.380 426.140 882.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 519.940 15.380 526.140 882.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 619.940 15.380 626.140 882.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 719.940 15.380 726.140 882.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 819.940 15.380 826.140 882.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 919.940 15.380 926.140 882.300 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 69.940 15.380 76.140 882.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 169.940 15.380 176.140 882.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 269.940 15.380 276.140 882.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 369.940 15.380 376.140 882.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 469.940 15.380 476.140 882.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 569.940 15.380 576.140 882.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 669.940 15.380 676.140 882.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 769.940 15.380 776.140 882.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 869.940 15.380 876.140 882.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 969.940 15.380 976.140 882.300 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 14.710 992.880 882.300 ;
      LAYER Metal2 ;
        RECT 7.980 895.700 43.380 896.420 ;
        RECT 44.540 895.700 126.260 896.420 ;
        RECT 127.420 895.700 209.140 896.420 ;
        RECT 210.300 895.700 292.020 896.420 ;
        RECT 293.180 895.700 374.900 896.420 ;
        RECT 376.060 895.700 457.780 896.420 ;
        RECT 458.940 895.700 540.660 896.420 ;
        RECT 541.820 895.700 623.540 896.420 ;
        RECT 624.700 895.700 706.420 896.420 ;
        RECT 707.580 895.700 789.300 896.420 ;
        RECT 790.460 895.700 872.180 896.420 ;
        RECT 873.340 895.700 955.060 896.420 ;
        RECT 956.220 895.700 992.180 896.420 ;
        RECT 7.980 4.300 992.180 895.700 ;
        RECT 7.980 3.500 25.460 4.300 ;
        RECT 26.620 3.500 45.620 4.300 ;
        RECT 46.780 3.500 65.780 4.300 ;
        RECT 66.940 3.500 85.940 4.300 ;
        RECT 87.100 3.500 106.100 4.300 ;
        RECT 107.260 3.500 126.260 4.300 ;
        RECT 127.420 3.500 146.420 4.300 ;
        RECT 147.580 3.500 166.580 4.300 ;
        RECT 167.740 3.500 186.740 4.300 ;
        RECT 187.900 3.500 206.900 4.300 ;
        RECT 208.060 3.500 227.060 4.300 ;
        RECT 228.220 3.500 247.220 4.300 ;
        RECT 248.380 3.500 267.380 4.300 ;
        RECT 268.540 3.500 287.540 4.300 ;
        RECT 288.700 3.500 307.700 4.300 ;
        RECT 308.860 3.500 327.860 4.300 ;
        RECT 329.020 3.500 348.020 4.300 ;
        RECT 349.180 3.500 368.180 4.300 ;
        RECT 369.340 3.500 388.340 4.300 ;
        RECT 389.500 3.500 408.500 4.300 ;
        RECT 409.660 3.500 428.660 4.300 ;
        RECT 429.820 3.500 448.820 4.300 ;
        RECT 449.980 3.500 468.980 4.300 ;
        RECT 470.140 3.500 489.140 4.300 ;
        RECT 490.300 3.500 509.300 4.300 ;
        RECT 510.460 3.500 529.460 4.300 ;
        RECT 530.620 3.500 549.620 4.300 ;
        RECT 550.780 3.500 569.780 4.300 ;
        RECT 570.940 3.500 589.940 4.300 ;
        RECT 591.100 3.500 610.100 4.300 ;
        RECT 611.260 3.500 630.260 4.300 ;
        RECT 631.420 3.500 650.420 4.300 ;
        RECT 651.580 3.500 670.580 4.300 ;
        RECT 671.740 3.500 690.740 4.300 ;
        RECT 691.900 3.500 710.900 4.300 ;
        RECT 712.060 3.500 731.060 4.300 ;
        RECT 732.220 3.500 751.220 4.300 ;
        RECT 752.380 3.500 771.380 4.300 ;
        RECT 772.540 3.500 791.540 4.300 ;
        RECT 792.700 3.500 811.700 4.300 ;
        RECT 812.860 3.500 831.860 4.300 ;
        RECT 833.020 3.500 852.020 4.300 ;
        RECT 853.180 3.500 872.180 4.300 ;
        RECT 873.340 3.500 892.340 4.300 ;
        RECT 893.500 3.500 912.500 4.300 ;
        RECT 913.660 3.500 932.660 4.300 ;
        RECT 933.820 3.500 952.820 4.300 ;
        RECT 953.980 3.500 972.980 4.300 ;
        RECT 974.140 3.500 992.180 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 880.060 996.000 882.140 ;
        RECT 4.300 878.900 996.000 880.060 ;
        RECT 4.000 868.860 996.000 878.900 ;
        RECT 4.000 867.700 995.700 868.860 ;
        RECT 4.000 853.180 996.000 867.700 ;
        RECT 4.300 852.020 996.000 853.180 ;
        RECT 4.000 826.300 996.000 852.020 ;
        RECT 4.300 825.140 996.000 826.300 ;
        RECT 4.000 819.580 996.000 825.140 ;
        RECT 4.000 818.420 995.700 819.580 ;
        RECT 4.000 799.420 996.000 818.420 ;
        RECT 4.300 798.260 996.000 799.420 ;
        RECT 4.000 772.540 996.000 798.260 ;
        RECT 4.300 771.380 996.000 772.540 ;
        RECT 4.000 770.300 996.000 771.380 ;
        RECT 4.000 769.140 995.700 770.300 ;
        RECT 4.000 745.660 996.000 769.140 ;
        RECT 4.300 744.500 996.000 745.660 ;
        RECT 4.000 721.020 996.000 744.500 ;
        RECT 4.000 719.860 995.700 721.020 ;
        RECT 4.000 718.780 996.000 719.860 ;
        RECT 4.300 717.620 996.000 718.780 ;
        RECT 4.000 691.900 996.000 717.620 ;
        RECT 4.300 690.740 996.000 691.900 ;
        RECT 4.000 671.740 996.000 690.740 ;
        RECT 4.000 670.580 995.700 671.740 ;
        RECT 4.000 665.020 996.000 670.580 ;
        RECT 4.300 663.860 996.000 665.020 ;
        RECT 4.000 638.140 996.000 663.860 ;
        RECT 4.300 636.980 996.000 638.140 ;
        RECT 4.000 622.460 996.000 636.980 ;
        RECT 4.000 621.300 995.700 622.460 ;
        RECT 4.000 611.260 996.000 621.300 ;
        RECT 4.300 610.100 996.000 611.260 ;
        RECT 4.000 584.380 996.000 610.100 ;
        RECT 4.300 583.220 996.000 584.380 ;
        RECT 4.000 573.180 996.000 583.220 ;
        RECT 4.000 572.020 995.700 573.180 ;
        RECT 4.000 557.500 996.000 572.020 ;
        RECT 4.300 556.340 996.000 557.500 ;
        RECT 4.000 530.620 996.000 556.340 ;
        RECT 4.300 529.460 996.000 530.620 ;
        RECT 4.000 523.900 996.000 529.460 ;
        RECT 4.000 522.740 995.700 523.900 ;
        RECT 4.000 503.740 996.000 522.740 ;
        RECT 4.300 502.580 996.000 503.740 ;
        RECT 4.000 476.860 996.000 502.580 ;
        RECT 4.300 475.700 996.000 476.860 ;
        RECT 4.000 474.620 996.000 475.700 ;
        RECT 4.000 473.460 995.700 474.620 ;
        RECT 4.000 449.980 996.000 473.460 ;
        RECT 4.300 448.820 996.000 449.980 ;
        RECT 4.000 425.340 996.000 448.820 ;
        RECT 4.000 424.180 995.700 425.340 ;
        RECT 4.000 423.100 996.000 424.180 ;
        RECT 4.300 421.940 996.000 423.100 ;
        RECT 4.000 396.220 996.000 421.940 ;
        RECT 4.300 395.060 996.000 396.220 ;
        RECT 4.000 376.060 996.000 395.060 ;
        RECT 4.000 374.900 995.700 376.060 ;
        RECT 4.000 369.340 996.000 374.900 ;
        RECT 4.300 368.180 996.000 369.340 ;
        RECT 4.000 342.460 996.000 368.180 ;
        RECT 4.300 341.300 996.000 342.460 ;
        RECT 4.000 326.780 996.000 341.300 ;
        RECT 4.000 325.620 995.700 326.780 ;
        RECT 4.000 315.580 996.000 325.620 ;
        RECT 4.300 314.420 996.000 315.580 ;
        RECT 4.000 288.700 996.000 314.420 ;
        RECT 4.300 287.540 996.000 288.700 ;
        RECT 4.000 277.500 996.000 287.540 ;
        RECT 4.000 276.340 995.700 277.500 ;
        RECT 4.000 261.820 996.000 276.340 ;
        RECT 4.300 260.660 996.000 261.820 ;
        RECT 4.000 234.940 996.000 260.660 ;
        RECT 4.300 233.780 996.000 234.940 ;
        RECT 4.000 228.220 996.000 233.780 ;
        RECT 4.000 227.060 995.700 228.220 ;
        RECT 4.000 208.060 996.000 227.060 ;
        RECT 4.300 206.900 996.000 208.060 ;
        RECT 4.000 181.180 996.000 206.900 ;
        RECT 4.300 180.020 996.000 181.180 ;
        RECT 4.000 178.940 996.000 180.020 ;
        RECT 4.000 177.780 995.700 178.940 ;
        RECT 4.000 154.300 996.000 177.780 ;
        RECT 4.300 153.140 996.000 154.300 ;
        RECT 4.000 129.660 996.000 153.140 ;
        RECT 4.000 128.500 995.700 129.660 ;
        RECT 4.000 127.420 996.000 128.500 ;
        RECT 4.300 126.260 996.000 127.420 ;
        RECT 4.000 100.540 996.000 126.260 ;
        RECT 4.300 99.380 996.000 100.540 ;
        RECT 4.000 80.380 996.000 99.380 ;
        RECT 4.000 79.220 995.700 80.380 ;
        RECT 4.000 73.660 996.000 79.220 ;
        RECT 4.300 72.500 996.000 73.660 ;
        RECT 4.000 46.780 996.000 72.500 ;
        RECT 4.300 45.620 996.000 46.780 ;
        RECT 4.000 31.100 996.000 45.620 ;
        RECT 4.000 29.940 995.700 31.100 ;
        RECT 4.000 19.900 996.000 29.940 ;
        RECT 4.300 18.740 996.000 19.900 ;
        RECT 4.000 12.460 996.000 18.740 ;
      LAYER Metal4 ;
        RECT 14.700 16.890 19.640 879.110 ;
        RECT 26.440 16.890 69.640 879.110 ;
        RECT 76.440 16.890 119.640 879.110 ;
        RECT 126.440 16.890 169.640 879.110 ;
        RECT 176.440 16.890 219.640 879.110 ;
        RECT 226.440 16.890 269.640 879.110 ;
        RECT 276.440 16.890 319.640 879.110 ;
        RECT 326.440 16.890 369.640 879.110 ;
        RECT 376.440 16.890 419.640 879.110 ;
        RECT 426.440 16.890 469.640 879.110 ;
        RECT 476.440 16.890 519.640 879.110 ;
        RECT 526.440 16.890 569.640 879.110 ;
        RECT 576.440 16.890 619.640 879.110 ;
        RECT 626.440 16.890 669.640 879.110 ;
        RECT 676.440 16.890 719.640 879.110 ;
        RECT 726.440 16.890 769.640 879.110 ;
        RECT 776.440 16.890 819.640 879.110 ;
        RECT 826.440 16.890 869.640 879.110 ;
        RECT 876.440 16.890 919.640 879.110 ;
        RECT 926.440 16.890 969.640 879.110 ;
        RECT 976.440 16.890 988.260 879.110 ;
      LAYER Metal5 ;
        RECT 14.620 17.330 966.500 781.870 ;
  END
END uart_i2c_usb_spi_top
END LIBRARY

