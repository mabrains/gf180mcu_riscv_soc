* NGSPICE file created from wb_buttons_leds.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VNW VPW VSS
.ends

.subckt wb_buttons_leds VDD VSS buttons[0] buttons[1] clk i_wb_addr[0] i_wb_addr[10]
+ i_wb_addr[11] i_wb_addr[12] i_wb_addr[13] i_wb_addr[14] i_wb_addr[15] i_wb_addr[16]
+ i_wb_addr[17] i_wb_addr[18] i_wb_addr[19] i_wb_addr[1] i_wb_addr[20] i_wb_addr[21]
+ i_wb_addr[22] i_wb_addr[23] i_wb_addr[24] i_wb_addr[25] i_wb_addr[26] i_wb_addr[27]
+ i_wb_addr[28] i_wb_addr[29] i_wb_addr[2] i_wb_addr[30] i_wb_addr[31] i_wb_addr[3]
+ i_wb_addr[4] i_wb_addr[5] i_wb_addr[6] i_wb_addr[7] i_wb_addr[8] i_wb_addr[9] i_wb_cyc
+ i_wb_data[0] i_wb_data[1] i_wb_stb i_wb_we leds[0] leds[1] o_wb_ack o_wb_data[0]
+ o_wb_data[15] o_wb_data[1] o_wb_data[20] o_wb_data[21] o_wb_data[22] o_wb_data[23]
+ o_wb_data[5] o_wb_stall reset o_wb_data[4] o_wb_data[14] o_wb_data[3] o_wb_data[25]
+ o_wb_data[13] o_wb_data[2] o_wb_data[24] o_wb_data[12] o_wb_data[11] o_wb_data[10]
+ o_wb_data[31] o_wb_data[9] o_wb_data[19] o_wb_data[30] o_wb_data[8] o_wb_data[29]
+ o_wb_data[18] o_wb_data[7] o_wb_data[28] o_wb_data[6] o_wb_data[17] o_wb_data[27]
+ o_wb_data[16] o_wb_data[26]
XFILLER_0_2_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_062_ _025_ _026_ _000_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input36_I i_wb_data[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_8_Left_25 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
Xwb_buttons_leds_63 o_wb_data[19] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__tiel
X_045_ net34 net33 net5 net4 _010_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xwb_buttons_leds_52 o_wb_data[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__tiel
Xwb_buttons_leds_74 o_wb_data[30] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_16_95 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_84 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput42 net42 leds[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_1_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input29_I i_wb_addr[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_83 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_12_Right_12 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_061_ net38 _008_ _026_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xwb_buttons_leds_53 o_wb_data[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__tiel
X_044_ net7 net6 net9 net8 _009_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xwb_buttons_leds_75 o_wb_data[31] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__tiel
Xwb_buttons_leds_64 o_wb_data[20] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_5_46 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input11_I i_wb_addr[17] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_6_Right_6 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_15_66 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput43 net43 o_wb_ack VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_input3_I i_wb_addr[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_129 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_060_ _022_ _024_ _025_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_10_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwb_buttons_leds_76 o_wb_stall VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__tiel
Xwb_buttons_leds_54 o_wb_data[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__tiel
Xwb_buttons_leds_65 o_wb_data[21] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_TAPCELL_ROW_5_47 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_043_ net40 _008_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_16_119 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_108 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_67 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput44 net44 o_wb_data[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_7_62 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_144 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input34_I i_wb_addr[9] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xwb_buttons_leds_66 o_wb_data[22] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__tiel
X_042_ net25 _007_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xwb_buttons_leds_55 o_wb_data[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_15_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_123 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput45 net45 o_wb_data[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_4_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input27_I i_wb_addr[31] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xwb_buttons_leds_67 o_wb_data[23] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__tiel
Xwb_buttons_leds_56 o_wb_data[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__tiel
X_041_ net36 _006_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_12_Left_29 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_15_Left_32 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input1_I buttons[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_0_Left_17 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwb_buttons_leds_68 o_wb_data[24] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__tiel
Xwb_buttons_leds_46 o_wb_data[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__tiel
Xwb_buttons_leds_57 o_wb_data[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__tiel
XPHY_EDGE_ROW_3_Left_20 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_040_ net37 _005_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_15_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_89 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_99 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xwb_buttons_leds_47 o_wb_data[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__tiel
Xwb_buttons_leds_69 o_wb_data[25] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__tiel
Xwb_buttons_leds_58 o_wb_data[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA_input32_I i_wb_addr[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_1_Right_1 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_7_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_70 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xwb_buttons_leds_48 o_wb_data[4] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__tiel
Xwb_buttons_leds_59 o_wb_data[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_15_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input25_I i_wb_addr[2] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_47 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_121 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_0_clk clk clknet_0_clk VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_15_Right_15 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_7_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_16_71 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_48 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xwb_buttons_leds_49 o_wb_data[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_11_81 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input18_I i_wb_addr[23] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_7_Left_24 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_59 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_117 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_42 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_62 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_079_ _005_ _037_ _039_ _004_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_input30_I i_wb_addr[5] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_5_Right_5 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_3_43 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_13_63 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_078_ net42 _037_ _008_ _039_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input23_I i_wb_addr[28] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_11_Right_11 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_4_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_34 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_54 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_077_ _006_ _037_ _038_ _003_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_input16_I i_wb_addr[21] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input8_I i_wb_addr[14] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_35 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_55 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput1 buttons[0] net1 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_11_Left_28 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_076_ net41 _037_ _008_ _038_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_0_clk_I clk VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_059_ _012_ _015_ _018_ _023_ _024_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XPHY_EDGE_ROW_9_Right_9 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_14_Left_31 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_14_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_36 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input39_I i_wb_we VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_64 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput2 buttons[1] net2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_10_56 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_075_ _015_ _018_ _031_ _036_ _037_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_058_ net25 _019_ _023_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input21_I i_wb_addr[26] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_37 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_109 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput3 i_wb_addr[0] net3 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_10_57 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_074_ net35 net38 net39 _036_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_7_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_057_ _012_ _015_ _018_ _021_ _022_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_3_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input14_I i_wb_addr[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_0_Right_0 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input6_I i_wb_addr[12] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput4 i_wb_addr[10] net4 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_11_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_48 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_073_ _033_ _034_ _035_ _002_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_2_97 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_056_ _007_ _019_ _021_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_16_68 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput40 reset net40 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_14_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput5 i_wb_addr[11] net5 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input37_I i_wb_data[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_49 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_072_ net45 _028_ _008_ _035_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_055_ net14 net3 net28 net25 _020_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XPHY_EDGE_ROW_6_Left_23 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_16_69 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput30 i_wb_addr[5] net30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_46 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput6 i_wb_addr[12] net6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_14_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_071_ net42 _022_ _034_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_14_Right_14 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_2_44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput31 i_wb_addr[6] net31 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput20 i_wb_addr[25] net20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_054_ net14 net3 net28 _019_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor3_1
XPHY_EDGE_ROW_4_Right_4 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input12_I i_wb_addr[18] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input4_I i_wb_addr[10] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput7 i_wb_addr[13] net7 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_070_ net2 _024_ _027_ net39 _033_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_053_ net24 net23 _016_ _017_ _018_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_TAPCELL_ROW_7_50 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput32 i_wb_addr[7] net32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput21 i_wb_addr[26] net21 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput10 i_wb_addr[16] net10 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput8 i_wb_addr[14] net8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_14_147 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input35_I i_wb_cyc VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_052_ net20 net19 net22 net21 _017_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xinput11 i_wb_addr[17] net11 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput33 i_wb_addr[8] net33 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_136 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_7_51 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput22 i_wb_addr[27] net22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_1_0__f_clk clknet_0_clk clknet_1_0__leaf_clk VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_8_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput9 i_wb_addr[15] net9 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_11_38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_10_Right_10 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input28_I i_wb_addr[3] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_051_ net27 net26 _016_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xinput12 i_wb_addr[18] net12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput34 i_wb_addr[9] net34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput23 i_wb_addr[28] net23 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_10_Left_27 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_8_Right_8 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input10_I i_wb_addr[16] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_13_Left_30 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_5_69 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input2_I buttons[1] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
X_050_ _013_ _014_ _015_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_4
Xinput13 i_wb_addr[19] net13 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput24 i_wb_addr[29] net24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput35 i_wb_cyc net35 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input40_I reset VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_70 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_150 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_131 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput25 i_wb_addr[2] net25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput14 i_wb_addr[1] net14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput36 i_wb_data[0] net36 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input33_I i_wb_addr[8] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_4_44 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_64 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_2_39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput15 i_wb_addr[20] net15 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput26 i_wb_addr[30] net26 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput37 i_wb_data[1] net37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input26_I i_wb_addr[30] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_45 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_65 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_2_Left_19 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_13_130 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput16 i_wb_addr[21] net16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput27 i_wb_addr[31] net27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput38 i_wb_stb net38 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input19_I i_wb_addr[24] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_5_Left_22 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_61 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput17 i_wb_addr[22] net17 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput28 i_wb_addr[3] net28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput39 i_wb_we net39 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input31_I i_wb_addr[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_3_Right_3 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_9_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_1_1__f_clk clknet_0_clk clknet_1_1__leaf_clk VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_6_118 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput18 i_wb_addr[23] net18 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput29 i_wb_addr[4] net29 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_85 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input24_I i_wb_addr[29] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_13_Right_13 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_1_38 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_30 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_103 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_58 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput19 i_wb_addr[24] net19 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2_122 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_20 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input17_I i_wb_addr[22] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_9_Left_26 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input9_I i_wb_addr[15] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_63 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_74 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_77 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_1_39 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_53 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_139 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_59 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_142 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_134 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_76 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_069_ _029_ _030_ _032_ _001_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_7_Right_7 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_12_68 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_068_ net44 _028_ _008_ _032_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input22_I i_wb_addr[27] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_32 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_133 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_22 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_141 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_2 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_114 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_2_40 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_60 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_084_ _004_ clknet_1_0__leaf_clk net42 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_067_ _009_ _010_ _011_ _020_ _031_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA_input15_I i_wb_addr[20] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input7_I i_wb_addr[13] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_101 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_6_34 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_41 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_115 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_24 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_79 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_61 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_083_ _003_ clknet_1_0__leaf_clk net41 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_25 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_12 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_066_ net41 _022_ _030_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xwb_buttons_leds_70 o_wb_data[26] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__tiel
X_049_ net11 net10 net13 net12 _014_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_16_146 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_135 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_113 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_80 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_16_Left_33 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_13_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_143 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_1_Left_18 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_2_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input38_I i_wb_stb VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
X_082_ _002_ clknet_1_1__leaf_clk net45 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_8_52 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_4_Left_21 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
X_065_ net1 _024_ _027_ net39 _029_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xwb_buttons_leds_60 o_wb_data[16] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__tiel
Xwb_buttons_leds_71 o_wb_data[27] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_16_125 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_048_ net16 net15 net18 net17 _013_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA_input20_I i_wb_addr[25] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_14 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_8 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_28 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_128 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_081_ _001_ clknet_1_1__leaf_clk net44 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_16_Right_16 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_8_53 VDD VSS gf180mcu_fd_sc_mcu7t5v0__filltie
X_064_ net39 _027_ _028_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_0_27 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_104 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xwb_buttons_leds_61 o_wb_data[17] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__tiel
Xwb_buttons_leds_72 o_wb_data[28] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__tiel
X_047_ _009_ _010_ _011_ _012_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand3_4
Xwb_buttons_leds_50 o_wb_data[6] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA_input13_I i_wb_addr[19] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_2_Right_2 VDD VSS gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_6_37 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input5_I i_wb_addr[11] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_6 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_5_137 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_148 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_107 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_16 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_151 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fill_1
X_080_ _000_ clknet_1_1__leaf_clk net43 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_72 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_063_ net35 net38 _027_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xwb_buttons_leds_51 o_wb_data[7] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__tiel
Xwb_buttons_leds_73 o_wb_data[29] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__tiel
X_046_ net30 net29 net32 net31 _011_ VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__nor4_4
Xwb_buttons_leds_62 o_wb_data[18] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_16_138 VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput41 net41 leds[0] VDD VDD VSS VSS gf180mcu_fd_sc_mcu7t5v0__buf_3
.ends

