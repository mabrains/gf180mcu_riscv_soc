`ifndef USER_PARMS
`define USER_PARMS


// ---- DEFINES ----
`define SEL_I2C   3'b001  // 0x3000_0040 --> 00110000000000000000000[001]000000
`define SEL_USB   3'b010  // 0x3000_0080 --> 00110000000000000000000[010]000000
`define SEL_SPI   3'b011  // 0x3000_00C0 --> 00110000000000000000000[011]000000
`define SEL_UART0 3'b100  // 0x3000_0100 --> 00110000000000000000000[100]000000
`define SEL_UART1 3'b111  // 0x3000_01C0 --> 00110000000000000000000[111]000000

//----------------------------------------------------------------------------
// Pinumux/Peri Reg Map - 0x3000_0600 --> 0011000000000000000000[10000]00000
//                      : 0x3000_06FF --> 0011000000000000000000[10111]11111

`define SEL_GLBL    5'b10000   // GLOBAL REGISTER
`define SEL_GPIO    5'b10001   // GPIO REGISTER
`define SEL_PWM     5'b10010   // PWM REGISTER
`define SEL_TIMER   5'b10011   // TIMER REGISTER
`define SEL_PERI    1'b1       // Peripheral
`define SEL_RTC     5'b10100   // RTC REGISTER

// ----- WB-Testing -----
`define LED_ADDRESS     32'h3000_0000   // BASE ADR
`define BUTTON_ADDRESS  32'h3000_0004   // BASE ADR + 4

// ---- Analog-TEMP-SENSOR ----
`define TEMP_SENS_ADDRESS     32'h3000_0008   // BASE ADR + 8

`endif // USER_PARMS
