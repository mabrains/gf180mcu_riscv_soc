magic
tech gf180mcuD
magscale 1 10
timestamp 1698594339
<< metal1 >>
rect 1344 96458 38640 96492
rect 1344 96406 4478 96458
rect 4530 96406 4582 96458
rect 4634 96406 4686 96458
rect 4738 96406 35198 96458
rect 35250 96406 35302 96458
rect 35354 96406 35406 96458
rect 35458 96406 38640 96458
rect 1344 96372 38640 96406
rect 3614 95954 3666 95966
rect 3614 95890 3666 95902
rect 1344 95674 38640 95708
rect 1344 95622 19838 95674
rect 19890 95622 19942 95674
rect 19994 95622 20046 95674
rect 20098 95622 38640 95674
rect 1344 95588 38640 95622
rect 1344 94890 38640 94924
rect 1344 94838 4478 94890
rect 4530 94838 4582 94890
rect 4634 94838 4686 94890
rect 4738 94838 35198 94890
rect 35250 94838 35302 94890
rect 35354 94838 35406 94890
rect 35458 94838 38640 94890
rect 1344 94804 38640 94838
rect 1344 94106 38640 94140
rect 1344 94054 19838 94106
rect 19890 94054 19942 94106
rect 19994 94054 20046 94106
rect 20098 94054 38640 94106
rect 1344 94020 38640 94054
rect 1344 93322 38640 93356
rect 1344 93270 4478 93322
rect 4530 93270 4582 93322
rect 4634 93270 4686 93322
rect 4738 93270 35198 93322
rect 35250 93270 35302 93322
rect 35354 93270 35406 93322
rect 35458 93270 38640 93322
rect 1344 93236 38640 93270
rect 1344 92538 38640 92572
rect 1344 92486 19838 92538
rect 19890 92486 19942 92538
rect 19994 92486 20046 92538
rect 20098 92486 38640 92538
rect 1344 92452 38640 92486
rect 1344 91754 38640 91788
rect 1344 91702 4478 91754
rect 4530 91702 4582 91754
rect 4634 91702 4686 91754
rect 4738 91702 35198 91754
rect 35250 91702 35302 91754
rect 35354 91702 35406 91754
rect 35458 91702 38640 91754
rect 1344 91668 38640 91702
rect 1344 90970 38640 91004
rect 1344 90918 19838 90970
rect 19890 90918 19942 90970
rect 19994 90918 20046 90970
rect 20098 90918 38640 90970
rect 1344 90884 38640 90918
rect 1344 90186 38640 90220
rect 1344 90134 4478 90186
rect 4530 90134 4582 90186
rect 4634 90134 4686 90186
rect 4738 90134 35198 90186
rect 35250 90134 35302 90186
rect 35354 90134 35406 90186
rect 35458 90134 38640 90186
rect 1344 90100 38640 90134
rect 1344 89402 38640 89436
rect 1344 89350 19838 89402
rect 19890 89350 19942 89402
rect 19994 89350 20046 89402
rect 20098 89350 38640 89402
rect 1344 89316 38640 89350
rect 1344 88618 38640 88652
rect 1344 88566 4478 88618
rect 4530 88566 4582 88618
rect 4634 88566 4686 88618
rect 4738 88566 35198 88618
rect 35250 88566 35302 88618
rect 35354 88566 35406 88618
rect 35458 88566 38640 88618
rect 1344 88532 38640 88566
rect 1344 87834 38640 87868
rect 1344 87782 19838 87834
rect 19890 87782 19942 87834
rect 19994 87782 20046 87834
rect 20098 87782 38640 87834
rect 1344 87748 38640 87782
rect 1344 87050 38640 87084
rect 1344 86998 4478 87050
rect 4530 86998 4582 87050
rect 4634 86998 4686 87050
rect 4738 86998 35198 87050
rect 35250 86998 35302 87050
rect 35354 86998 35406 87050
rect 35458 86998 38640 87050
rect 1344 86964 38640 86998
rect 1344 86266 38640 86300
rect 1344 86214 19838 86266
rect 19890 86214 19942 86266
rect 19994 86214 20046 86266
rect 20098 86214 38640 86266
rect 1344 86180 38640 86214
rect 1344 85482 38640 85516
rect 1344 85430 4478 85482
rect 4530 85430 4582 85482
rect 4634 85430 4686 85482
rect 4738 85430 35198 85482
rect 35250 85430 35302 85482
rect 35354 85430 35406 85482
rect 35458 85430 38640 85482
rect 1344 85396 38640 85430
rect 1344 84698 38640 84732
rect 1344 84646 19838 84698
rect 19890 84646 19942 84698
rect 19994 84646 20046 84698
rect 20098 84646 38640 84698
rect 1344 84612 38640 84646
rect 1344 83914 38640 83948
rect 1344 83862 4478 83914
rect 4530 83862 4582 83914
rect 4634 83862 4686 83914
rect 4738 83862 35198 83914
rect 35250 83862 35302 83914
rect 35354 83862 35406 83914
rect 35458 83862 38640 83914
rect 1344 83828 38640 83862
rect 1344 83130 38640 83164
rect 1344 83078 19838 83130
rect 19890 83078 19942 83130
rect 19994 83078 20046 83130
rect 20098 83078 38640 83130
rect 1344 83044 38640 83078
rect 1344 82346 38640 82380
rect 1344 82294 4478 82346
rect 4530 82294 4582 82346
rect 4634 82294 4686 82346
rect 4738 82294 35198 82346
rect 35250 82294 35302 82346
rect 35354 82294 35406 82346
rect 35458 82294 38640 82346
rect 1344 82260 38640 82294
rect 1344 81562 38640 81596
rect 1344 81510 19838 81562
rect 19890 81510 19942 81562
rect 19994 81510 20046 81562
rect 20098 81510 38640 81562
rect 1344 81476 38640 81510
rect 1344 80778 38640 80812
rect 1344 80726 4478 80778
rect 4530 80726 4582 80778
rect 4634 80726 4686 80778
rect 4738 80726 35198 80778
rect 35250 80726 35302 80778
rect 35354 80726 35406 80778
rect 35458 80726 38640 80778
rect 1344 80692 38640 80726
rect 1344 79994 38640 80028
rect 1344 79942 19838 79994
rect 19890 79942 19942 79994
rect 19994 79942 20046 79994
rect 20098 79942 38640 79994
rect 1344 79908 38640 79942
rect 1344 79210 38640 79244
rect 1344 79158 4478 79210
rect 4530 79158 4582 79210
rect 4634 79158 4686 79210
rect 4738 79158 35198 79210
rect 35250 79158 35302 79210
rect 35354 79158 35406 79210
rect 35458 79158 38640 79210
rect 1344 79124 38640 79158
rect 1344 78426 38640 78460
rect 1344 78374 19838 78426
rect 19890 78374 19942 78426
rect 19994 78374 20046 78426
rect 20098 78374 38640 78426
rect 1344 78340 38640 78374
rect 1344 77642 38640 77676
rect 1344 77590 4478 77642
rect 4530 77590 4582 77642
rect 4634 77590 4686 77642
rect 4738 77590 35198 77642
rect 35250 77590 35302 77642
rect 35354 77590 35406 77642
rect 35458 77590 38640 77642
rect 1344 77556 38640 77590
rect 1344 76858 38640 76892
rect 1344 76806 19838 76858
rect 19890 76806 19942 76858
rect 19994 76806 20046 76858
rect 20098 76806 38640 76858
rect 1344 76772 38640 76806
rect 1344 76074 38640 76108
rect 1344 76022 4478 76074
rect 4530 76022 4582 76074
rect 4634 76022 4686 76074
rect 4738 76022 35198 76074
rect 35250 76022 35302 76074
rect 35354 76022 35406 76074
rect 35458 76022 38640 76074
rect 1344 75988 38640 76022
rect 1344 75290 38640 75324
rect 1344 75238 19838 75290
rect 19890 75238 19942 75290
rect 19994 75238 20046 75290
rect 20098 75238 38640 75290
rect 1344 75204 38640 75238
rect 1344 74506 38640 74540
rect 1344 74454 4478 74506
rect 4530 74454 4582 74506
rect 4634 74454 4686 74506
rect 4738 74454 35198 74506
rect 35250 74454 35302 74506
rect 35354 74454 35406 74506
rect 35458 74454 38640 74506
rect 1344 74420 38640 74454
rect 1344 73722 38640 73756
rect 1344 73670 19838 73722
rect 19890 73670 19942 73722
rect 19994 73670 20046 73722
rect 20098 73670 38640 73722
rect 1344 73636 38640 73670
rect 1344 72938 38640 72972
rect 1344 72886 4478 72938
rect 4530 72886 4582 72938
rect 4634 72886 4686 72938
rect 4738 72886 35198 72938
rect 35250 72886 35302 72938
rect 35354 72886 35406 72938
rect 35458 72886 38640 72938
rect 1344 72852 38640 72886
rect 1344 72154 38640 72188
rect 1344 72102 19838 72154
rect 19890 72102 19942 72154
rect 19994 72102 20046 72154
rect 20098 72102 38640 72154
rect 1344 72068 38640 72102
rect 1344 71370 38640 71404
rect 1344 71318 4478 71370
rect 4530 71318 4582 71370
rect 4634 71318 4686 71370
rect 4738 71318 35198 71370
rect 35250 71318 35302 71370
rect 35354 71318 35406 71370
rect 35458 71318 38640 71370
rect 1344 71284 38640 71318
rect 1344 70586 38640 70620
rect 1344 70534 19838 70586
rect 19890 70534 19942 70586
rect 19994 70534 20046 70586
rect 20098 70534 38640 70586
rect 1344 70500 38640 70534
rect 25342 70306 25394 70318
rect 25342 70242 25394 70254
rect 20078 70194 20130 70206
rect 17938 70142 17950 70194
rect 18002 70142 18014 70194
rect 19842 70142 19854 70194
rect 19906 70142 19918 70194
rect 20078 70130 20130 70142
rect 20190 70194 20242 70206
rect 20190 70130 20242 70142
rect 25566 70082 25618 70094
rect 25566 70018 25618 70030
rect 26126 70082 26178 70094
rect 26126 70018 26178 70030
rect 18174 69970 18226 69982
rect 18174 69906 18226 69918
rect 18398 69970 18450 69982
rect 18398 69906 18450 69918
rect 18510 69970 18562 69982
rect 25230 69970 25282 69982
rect 20626 69918 20638 69970
rect 20690 69918 20702 69970
rect 18510 69906 18562 69918
rect 25230 69906 25282 69918
rect 1344 69802 38640 69836
rect 1344 69750 4478 69802
rect 4530 69750 4582 69802
rect 4634 69750 4686 69802
rect 4738 69750 35198 69802
rect 35250 69750 35302 69802
rect 35354 69750 35406 69802
rect 35458 69750 38640 69802
rect 1344 69716 38640 69750
rect 20638 69634 20690 69646
rect 20638 69570 20690 69582
rect 20414 69522 20466 69534
rect 22306 69470 22318 69522
rect 22370 69470 22382 69522
rect 24434 69470 24446 69522
rect 24498 69470 24510 69522
rect 20414 69458 20466 69470
rect 15262 69410 15314 69422
rect 18398 69410 18450 69422
rect 16594 69358 16606 69410
rect 16658 69358 16670 69410
rect 17826 69358 17838 69410
rect 17890 69358 17902 69410
rect 19058 69358 19070 69410
rect 19122 69358 19134 69410
rect 20178 69358 20190 69410
rect 20242 69358 20254 69410
rect 25218 69358 25230 69410
rect 25282 69358 25294 69410
rect 25554 69358 25566 69410
rect 25618 69358 25630 69410
rect 15262 69346 15314 69358
rect 18398 69346 18450 69358
rect 20750 69298 20802 69310
rect 19618 69246 19630 69298
rect 19682 69246 19694 69298
rect 20750 69234 20802 69246
rect 25790 69298 25842 69310
rect 25790 69234 25842 69246
rect 25902 69298 25954 69310
rect 25902 69234 25954 69246
rect 15822 69186 15874 69198
rect 15822 69122 15874 69134
rect 16830 69186 16882 69198
rect 26338 69134 26350 69186
rect 26402 69134 26414 69186
rect 16830 69122 16882 69134
rect 1344 69018 38640 69052
rect 1344 68966 19838 69018
rect 19890 68966 19942 69018
rect 19994 68966 20046 69018
rect 20098 68966 38640 69018
rect 1344 68932 38640 68966
rect 17614 68850 17666 68862
rect 17614 68786 17666 68798
rect 2046 68738 2098 68750
rect 2046 68674 2098 68686
rect 9662 68738 9714 68750
rect 9662 68674 9714 68686
rect 9774 68738 9826 68750
rect 9774 68674 9826 68686
rect 17390 68738 17442 68750
rect 25230 68738 25282 68750
rect 24658 68686 24670 68738
rect 24722 68686 24734 68738
rect 17390 68674 17442 68686
rect 25230 68674 25282 68686
rect 25790 68738 25842 68750
rect 25790 68674 25842 68686
rect 1710 68626 1762 68638
rect 18958 68626 19010 68638
rect 24334 68626 24386 68638
rect 10322 68574 10334 68626
rect 10386 68574 10398 68626
rect 13682 68574 13694 68626
rect 13746 68574 13758 68626
rect 18498 68574 18510 68626
rect 18562 68574 18574 68626
rect 19618 68574 19630 68626
rect 19682 68574 19694 68626
rect 23986 68574 23998 68626
rect 24050 68574 24062 68626
rect 1710 68562 1762 68574
rect 18958 68562 19010 68574
rect 24334 68562 24386 68574
rect 25454 68626 25506 68638
rect 28914 68574 28926 68626
rect 28978 68574 28990 68626
rect 25454 68562 25506 68574
rect 2494 68514 2546 68526
rect 25678 68514 25730 68526
rect 10994 68462 11006 68514
rect 11058 68462 11070 68514
rect 13234 68462 13246 68514
rect 13298 68462 13310 68514
rect 14466 68462 14478 68514
rect 14530 68462 14542 68514
rect 16594 68462 16606 68514
rect 16658 68462 16670 68514
rect 17714 68462 17726 68514
rect 17778 68462 17790 68514
rect 21074 68462 21086 68514
rect 21138 68462 21150 68514
rect 23202 68462 23214 68514
rect 23266 68462 23278 68514
rect 26114 68462 26126 68514
rect 26178 68462 26190 68514
rect 28242 68462 28254 68514
rect 28306 68462 28318 68514
rect 2494 68450 2546 68462
rect 25678 68450 25730 68462
rect 9774 68402 9826 68414
rect 20178 68350 20190 68402
rect 20242 68350 20254 68402
rect 9774 68338 9826 68350
rect 1344 68234 38640 68268
rect 1344 68182 4478 68234
rect 4530 68182 4582 68234
rect 4634 68182 4686 68234
rect 4738 68182 35198 68234
rect 35250 68182 35302 68234
rect 35354 68182 35406 68234
rect 35458 68182 38640 68234
rect 1344 68148 38640 68182
rect 7646 67954 7698 67966
rect 7646 67890 7698 67902
rect 11006 67954 11058 67966
rect 11006 67890 11058 67902
rect 19630 67954 19682 67966
rect 20514 67902 20526 67954
rect 20578 67902 20590 67954
rect 24546 67902 24558 67954
rect 24610 67902 24622 67954
rect 28578 67902 28590 67954
rect 28642 67902 28654 67954
rect 19630 67890 19682 67902
rect 10782 67842 10834 67854
rect 10546 67790 10558 67842
rect 10610 67790 10622 67842
rect 10782 67778 10834 67790
rect 11790 67842 11842 67854
rect 11790 67778 11842 67790
rect 12126 67842 12178 67854
rect 12126 67778 12178 67790
rect 12574 67842 12626 67854
rect 23550 67842 23602 67854
rect 14130 67790 14142 67842
rect 14194 67790 14206 67842
rect 15474 67790 15486 67842
rect 15538 67790 15550 67842
rect 17714 67790 17726 67842
rect 17778 67790 17790 67842
rect 20066 67790 20078 67842
rect 20130 67790 20142 67842
rect 24658 67790 24670 67842
rect 24722 67790 24734 67842
rect 25778 67790 25790 67842
rect 25842 67790 25854 67842
rect 12574 67778 12626 67790
rect 23550 67778 23602 67790
rect 1710 67730 1762 67742
rect 11230 67730 11282 67742
rect 9762 67678 9774 67730
rect 9826 67678 9838 67730
rect 1710 67666 1762 67678
rect 11230 67666 11282 67678
rect 11454 67730 11506 67742
rect 11454 67666 11506 67678
rect 12350 67730 12402 67742
rect 12350 67666 12402 67678
rect 12910 67730 12962 67742
rect 12910 67666 12962 67678
rect 16718 67730 16770 67742
rect 16718 67666 16770 67678
rect 18174 67730 18226 67742
rect 24222 67730 24274 67742
rect 23874 67678 23886 67730
rect 23938 67678 23950 67730
rect 26450 67678 26462 67730
rect 26514 67678 26526 67730
rect 18174 67666 18226 67678
rect 24222 67666 24274 67678
rect 2046 67618 2098 67630
rect 2046 67554 2098 67566
rect 2494 67618 2546 67630
rect 2494 67554 2546 67566
rect 11902 67618 11954 67630
rect 11902 67554 11954 67566
rect 12798 67618 12850 67630
rect 12798 67554 12850 67566
rect 13582 67618 13634 67630
rect 13582 67554 13634 67566
rect 14478 67618 14530 67630
rect 14478 67554 14530 67566
rect 16270 67618 16322 67630
rect 16270 67554 16322 67566
rect 1344 67450 38640 67484
rect 1344 67398 19838 67450
rect 19890 67398 19942 67450
rect 19994 67398 20046 67450
rect 20098 67398 38640 67450
rect 1344 67364 38640 67398
rect 9774 67282 9826 67294
rect 23214 67282 23266 67294
rect 13906 67230 13918 67282
rect 13970 67230 13982 67282
rect 9774 67218 9826 67230
rect 23214 67218 23266 67230
rect 2046 67170 2098 67182
rect 2046 67106 2098 67118
rect 8206 67170 8258 67182
rect 8206 67106 8258 67118
rect 8318 67170 8370 67182
rect 8318 67106 8370 67118
rect 8542 67170 8594 67182
rect 8542 67106 8594 67118
rect 8766 67170 8818 67182
rect 8766 67106 8818 67118
rect 8878 67170 8930 67182
rect 8878 67106 8930 67118
rect 10110 67170 10162 67182
rect 16830 67170 16882 67182
rect 11666 67118 11678 67170
rect 11730 67118 11742 67170
rect 10110 67106 10162 67118
rect 16830 67106 16882 67118
rect 17390 67170 17442 67182
rect 17390 67106 17442 67118
rect 20190 67170 20242 67182
rect 20190 67106 20242 67118
rect 25454 67170 25506 67182
rect 25454 67106 25506 67118
rect 25566 67170 25618 67182
rect 25566 67106 25618 67118
rect 26462 67170 26514 67182
rect 26462 67106 26514 67118
rect 27582 67170 27634 67182
rect 27582 67106 27634 67118
rect 1710 67058 1762 67070
rect 1710 66994 1762 67006
rect 9102 67058 9154 67070
rect 9102 66994 9154 67006
rect 9438 67058 9490 67070
rect 9438 66994 9490 67006
rect 9774 67058 9826 67070
rect 17838 67058 17890 67070
rect 10882 67006 10894 67058
rect 10946 67006 10958 67058
rect 9774 66994 9826 67006
rect 17838 66994 17890 67006
rect 18062 67058 18114 67070
rect 25230 67058 25282 67070
rect 26238 67058 26290 67070
rect 20402 67006 20414 67058
rect 20466 67006 20478 67058
rect 21298 67006 21310 67058
rect 21362 67006 21374 67058
rect 22978 67006 22990 67058
rect 23042 67006 23054 67058
rect 25778 67006 25790 67058
rect 25842 67006 25854 67058
rect 18062 66994 18114 67006
rect 25230 66994 25282 67006
rect 26238 66994 26290 67006
rect 26798 67058 26850 67070
rect 27470 67058 27522 67070
rect 27010 67006 27022 67058
rect 27074 67006 27086 67058
rect 26798 66994 26850 67006
rect 27470 66994 27522 67006
rect 2494 66946 2546 66958
rect 18610 66894 18622 66946
rect 18674 66894 18686 66946
rect 21410 66894 21422 66946
rect 21474 66894 21486 66946
rect 2494 66882 2546 66894
rect 16718 66834 16770 66846
rect 16718 66770 16770 66782
rect 17614 66834 17666 66846
rect 26574 66834 26626 66846
rect 21186 66782 21198 66834
rect 21250 66782 21262 66834
rect 17614 66770 17666 66782
rect 26574 66770 26626 66782
rect 27358 66834 27410 66846
rect 27358 66770 27410 66782
rect 1344 66666 38640 66700
rect 1344 66614 4478 66666
rect 4530 66614 4582 66666
rect 4634 66614 4686 66666
rect 4738 66614 35198 66666
rect 35250 66614 35302 66666
rect 35354 66614 35406 66666
rect 35458 66614 38640 66666
rect 1344 66580 38640 66614
rect 26462 66498 26514 66510
rect 26462 66434 26514 66446
rect 26798 66498 26850 66510
rect 26798 66434 26850 66446
rect 9886 66274 9938 66286
rect 9886 66210 9938 66222
rect 10222 66274 10274 66286
rect 10222 66210 10274 66222
rect 12574 66274 12626 66286
rect 12574 66210 12626 66222
rect 12910 66274 12962 66286
rect 26686 66274 26738 66286
rect 26226 66222 26238 66274
rect 26290 66222 26302 66274
rect 12910 66210 12962 66222
rect 26686 66210 26738 66222
rect 9662 66050 9714 66062
rect 9662 65986 9714 65998
rect 9998 66050 10050 66062
rect 9998 65986 10050 65998
rect 12350 66050 12402 66062
rect 12350 65986 12402 65998
rect 12798 66050 12850 66062
rect 12798 65986 12850 65998
rect 27246 66050 27298 66062
rect 27246 65986 27298 65998
rect 1344 65882 38640 65916
rect 1344 65830 19838 65882
rect 19890 65830 19942 65882
rect 19994 65830 20046 65882
rect 20098 65830 38640 65882
rect 1344 65796 38640 65830
rect 24334 65602 24386 65614
rect 24334 65538 24386 65550
rect 24446 65490 24498 65502
rect 23874 65438 23886 65490
rect 23938 65438 23950 65490
rect 24658 65438 24670 65490
rect 24722 65438 24734 65490
rect 24446 65426 24498 65438
rect 2158 65378 2210 65390
rect 2158 65314 2210 65326
rect 25342 65378 25394 65390
rect 25342 65314 25394 65326
rect 25790 65378 25842 65390
rect 25790 65314 25842 65326
rect 1344 65098 38640 65132
rect 1344 65046 4478 65098
rect 4530 65046 4582 65098
rect 4634 65046 4686 65098
rect 4738 65046 35198 65098
rect 35250 65046 35302 65098
rect 35354 65046 35406 65098
rect 35458 65046 38640 65098
rect 1344 65012 38640 65046
rect 14030 64706 14082 64718
rect 1810 64654 1822 64706
rect 1874 64654 1886 64706
rect 9314 64654 9326 64706
rect 9378 64654 9390 64706
rect 14030 64642 14082 64654
rect 14142 64706 14194 64718
rect 14466 64654 14478 64706
rect 14530 64654 14542 64706
rect 14142 64642 14194 64654
rect 2382 64594 2434 64606
rect 2382 64530 2434 64542
rect 2718 64594 2770 64606
rect 2718 64530 2770 64542
rect 8654 64594 8706 64606
rect 8654 64530 8706 64542
rect 8766 64594 8818 64606
rect 13694 64594 13746 64606
rect 9986 64542 9998 64594
rect 10050 64542 10062 64594
rect 8766 64530 8818 64542
rect 13694 64530 13746 64542
rect 2046 64482 2098 64494
rect 2046 64418 2098 64430
rect 3166 64482 3218 64494
rect 3166 64418 3218 64430
rect 8990 64482 9042 64494
rect 25678 64482 25730 64494
rect 12674 64430 12686 64482
rect 12738 64430 12750 64482
rect 14130 64430 14142 64482
rect 14194 64430 14206 64482
rect 8990 64418 9042 64430
rect 25678 64418 25730 64430
rect 38222 64482 38274 64494
rect 38222 64418 38274 64430
rect 1344 64314 38640 64348
rect 1344 64262 19838 64314
rect 19890 64262 19942 64314
rect 19994 64262 20046 64314
rect 20098 64262 38640 64314
rect 1344 64228 38640 64262
rect 10446 64146 10498 64158
rect 9986 64094 9998 64146
rect 10050 64094 10062 64146
rect 10446 64082 10498 64094
rect 11118 64146 11170 64158
rect 11118 64082 11170 64094
rect 11342 64146 11394 64158
rect 11342 64082 11394 64094
rect 13358 64146 13410 64158
rect 13358 64082 13410 64094
rect 14478 64146 14530 64158
rect 14478 64082 14530 64094
rect 2046 64034 2098 64046
rect 2046 63970 2098 63982
rect 10670 64034 10722 64046
rect 10670 63970 10722 63982
rect 13918 64034 13970 64046
rect 13918 63970 13970 63982
rect 14590 64034 14642 64046
rect 20190 64034 20242 64046
rect 17938 63982 17950 64034
rect 18002 63982 18014 64034
rect 14590 63970 14642 63982
rect 20190 63970 20242 63982
rect 26238 64034 26290 64046
rect 26238 63970 26290 63982
rect 1710 63922 1762 63934
rect 1710 63858 1762 63870
rect 2494 63922 2546 63934
rect 10222 63922 10274 63934
rect 9762 63870 9774 63922
rect 9826 63870 9838 63922
rect 2494 63858 2546 63870
rect 10222 63858 10274 63870
rect 10894 63922 10946 63934
rect 10894 63858 10946 63870
rect 11454 63922 11506 63934
rect 25790 63922 25842 63934
rect 18274 63870 18286 63922
rect 18338 63870 18350 63922
rect 18946 63870 18958 63922
rect 19010 63870 19022 63922
rect 24322 63870 24334 63922
rect 24386 63870 24398 63922
rect 26786 63870 26798 63922
rect 26850 63870 26862 63922
rect 11454 63858 11506 63870
rect 25790 63858 25842 63870
rect 13694 63810 13746 63822
rect 13694 63746 13746 63758
rect 13806 63810 13858 63822
rect 13806 63746 13858 63758
rect 19630 63810 19682 63822
rect 25566 63810 25618 63822
rect 29598 63810 29650 63822
rect 21410 63758 21422 63810
rect 21474 63758 21486 63810
rect 23538 63758 23550 63810
rect 23602 63758 23614 63810
rect 27458 63758 27470 63810
rect 27522 63758 27534 63810
rect 19630 63746 19682 63758
rect 25566 63746 25618 63758
rect 29598 63746 29650 63758
rect 14366 63698 14418 63710
rect 14366 63634 14418 63646
rect 19966 63698 20018 63710
rect 19966 63634 20018 63646
rect 20302 63698 20354 63710
rect 20302 63634 20354 63646
rect 25230 63698 25282 63710
rect 25230 63634 25282 63646
rect 1344 63530 38640 63564
rect 1344 63478 4478 63530
rect 4530 63478 4582 63530
rect 4634 63478 4686 63530
rect 4738 63478 35198 63530
rect 35250 63478 35302 63530
rect 35354 63478 35406 63530
rect 35458 63478 38640 63530
rect 1344 63444 38640 63478
rect 18062 63362 18114 63374
rect 18062 63298 18114 63310
rect 27458 63198 27470 63250
rect 27522 63198 27534 63250
rect 9886 63138 9938 63150
rect 17390 63138 17442 63150
rect 13570 63086 13582 63138
rect 13634 63086 13646 63138
rect 9886 63074 9938 63086
rect 17390 63074 17442 63086
rect 17838 63138 17890 63150
rect 22766 63138 22818 63150
rect 19394 63086 19406 63138
rect 19458 63086 19470 63138
rect 20290 63086 20302 63138
rect 20354 63086 20366 63138
rect 17838 63074 17890 63086
rect 22766 63074 22818 63086
rect 23326 63138 23378 63150
rect 24894 63138 24946 63150
rect 24658 63086 24670 63138
rect 24722 63086 24734 63138
rect 23326 63074 23378 63086
rect 24894 63074 24946 63086
rect 25230 63138 25282 63150
rect 25230 63074 25282 63086
rect 26014 63138 26066 63150
rect 28030 63138 28082 63150
rect 26226 63086 26238 63138
rect 26290 63086 26302 63138
rect 27570 63086 27582 63138
rect 27634 63086 27646 63138
rect 26014 63074 26066 63086
rect 28030 63074 28082 63086
rect 1710 63026 1762 63038
rect 1710 62962 1762 62974
rect 2046 63026 2098 63038
rect 2046 62962 2098 62974
rect 8878 63026 8930 63038
rect 8878 62962 8930 62974
rect 8990 63026 9042 63038
rect 17278 63026 17330 63038
rect 23662 63026 23714 63038
rect 14242 62974 14254 63026
rect 14306 62974 14318 63026
rect 18834 62974 18846 63026
rect 18898 62974 18910 63026
rect 8990 62962 9042 62974
rect 17278 62962 17330 62974
rect 23662 62962 23714 62974
rect 23998 63026 24050 63038
rect 23998 62962 24050 62974
rect 24222 63026 24274 63038
rect 24222 62962 24274 62974
rect 25006 63026 25058 63038
rect 25006 62962 25058 62974
rect 26910 63026 26962 63038
rect 26910 62962 26962 62974
rect 27246 63026 27298 63038
rect 27246 62962 27298 62974
rect 2494 62914 2546 62926
rect 2494 62850 2546 62862
rect 9214 62914 9266 62926
rect 18174 62914 18226 62926
rect 10210 62862 10222 62914
rect 10274 62862 10286 62914
rect 16482 62862 16494 62914
rect 16546 62862 16558 62914
rect 20402 62862 20414 62914
rect 20466 62862 20478 62914
rect 9214 62850 9266 62862
rect 18174 62850 18226 62862
rect 1344 62746 38640 62780
rect 1344 62694 19838 62746
rect 19890 62694 19942 62746
rect 19994 62694 20046 62746
rect 20098 62694 38640 62746
rect 1344 62660 38640 62694
rect 13246 62578 13298 62590
rect 8082 62526 8094 62578
rect 8146 62526 8158 62578
rect 13246 62514 13298 62526
rect 14254 62578 14306 62590
rect 16046 62578 16098 62590
rect 14690 62526 14702 62578
rect 14754 62526 14766 62578
rect 14254 62514 14306 62526
rect 16046 62514 16098 62526
rect 16830 62578 16882 62590
rect 16830 62514 16882 62526
rect 17502 62578 17554 62590
rect 17502 62514 17554 62526
rect 24334 62578 24386 62590
rect 24334 62514 24386 62526
rect 15710 62466 15762 62478
rect 14130 62414 14142 62466
rect 14194 62414 14206 62466
rect 15710 62402 15762 62414
rect 19518 62466 19570 62478
rect 24558 62466 24610 62478
rect 20178 62414 20190 62466
rect 20242 62414 20254 62466
rect 21522 62414 21534 62466
rect 21586 62414 21598 62466
rect 19518 62402 19570 62414
rect 24558 62402 24610 62414
rect 24670 62466 24722 62478
rect 24670 62402 24722 62414
rect 8542 62354 8594 62366
rect 7858 62302 7870 62354
rect 7922 62302 7934 62354
rect 8542 62290 8594 62302
rect 8766 62354 8818 62366
rect 8766 62290 8818 62302
rect 9102 62354 9154 62366
rect 14366 62354 14418 62366
rect 15598 62354 15650 62366
rect 17950 62354 18002 62366
rect 9538 62302 9550 62354
rect 9602 62302 9614 62354
rect 13682 62302 13694 62354
rect 13746 62302 13758 62354
rect 14914 62302 14926 62354
rect 14978 62302 14990 62354
rect 17602 62302 17614 62354
rect 17666 62302 17678 62354
rect 9102 62290 9154 62302
rect 14366 62290 14418 62302
rect 15598 62290 15650 62302
rect 17950 62290 18002 62302
rect 18958 62354 19010 62366
rect 24222 62354 24274 62366
rect 19282 62302 19294 62354
rect 19346 62302 19358 62354
rect 29026 62302 29038 62354
rect 29090 62302 29102 62354
rect 18958 62290 19010 62302
rect 24222 62290 24274 62302
rect 8878 62242 8930 62254
rect 19966 62242 20018 62254
rect 10322 62190 10334 62242
rect 10386 62190 10398 62242
rect 12450 62190 12462 62242
rect 12514 62190 12526 62242
rect 22082 62190 22094 62242
rect 22146 62190 22158 62242
rect 28466 62190 28478 62242
rect 28530 62190 28542 62242
rect 8878 62178 8930 62190
rect 19966 62178 20018 62190
rect 13918 62130 13970 62142
rect 13918 62066 13970 62078
rect 19630 62130 19682 62142
rect 19630 62066 19682 62078
rect 1344 61962 38640 61996
rect 1344 61910 4478 61962
rect 4530 61910 4582 61962
rect 4634 61910 4686 61962
rect 4738 61910 35198 61962
rect 35250 61910 35302 61962
rect 35354 61910 35406 61962
rect 35458 61910 38640 61962
rect 1344 61876 38640 61910
rect 19742 61794 19794 61806
rect 19742 61730 19794 61742
rect 23886 61682 23938 61694
rect 27122 61630 27134 61682
rect 27186 61630 27198 61682
rect 23886 61618 23938 61630
rect 8878 61570 8930 61582
rect 8418 61518 8430 61570
rect 8482 61518 8494 61570
rect 8878 61506 8930 61518
rect 9550 61570 9602 61582
rect 9550 61506 9602 61518
rect 10110 61570 10162 61582
rect 19294 61570 19346 61582
rect 13570 61518 13582 61570
rect 13634 61518 13646 61570
rect 10110 61506 10162 61518
rect 19294 61506 19346 61518
rect 19630 61570 19682 61582
rect 19630 61506 19682 61518
rect 20190 61570 20242 61582
rect 20190 61506 20242 61518
rect 20414 61570 20466 61582
rect 20414 61506 20466 61518
rect 23998 61570 24050 61582
rect 23998 61506 24050 61518
rect 24670 61570 24722 61582
rect 24670 61506 24722 61518
rect 24894 61570 24946 61582
rect 25218 61518 25230 61570
rect 25282 61518 25294 61570
rect 26898 61518 26910 61570
rect 26962 61518 26974 61570
rect 24894 61506 24946 61518
rect 10446 61458 10498 61470
rect 18734 61458 18786 61470
rect 13794 61406 13806 61458
rect 13858 61406 13870 61458
rect 10446 61394 10498 61406
rect 18734 61394 18786 61406
rect 18958 61458 19010 61470
rect 20750 61458 20802 61470
rect 18958 61394 19010 61406
rect 19742 61402 19794 61414
rect 9214 61346 9266 61358
rect 9214 61282 9266 61294
rect 10334 61346 10386 61358
rect 10334 61282 10386 61294
rect 19070 61346 19122 61358
rect 20750 61394 20802 61406
rect 23326 61458 23378 61470
rect 25778 61406 25790 61458
rect 25842 61406 25854 61458
rect 27010 61406 27022 61458
rect 27074 61406 27086 61458
rect 23326 61394 23378 61406
rect 19742 61338 19794 61350
rect 20414 61346 20466 61358
rect 19070 61282 19122 61294
rect 20414 61282 20466 61294
rect 23214 61346 23266 61358
rect 23214 61282 23266 61294
rect 24446 61346 24498 61358
rect 24446 61282 24498 61294
rect 24782 61346 24834 61358
rect 24782 61282 24834 61294
rect 1344 61178 38640 61212
rect 1344 61126 19838 61178
rect 19890 61126 19942 61178
rect 19994 61126 20046 61178
rect 20098 61126 38640 61178
rect 1344 61092 38640 61126
rect 22206 61010 22258 61022
rect 22206 60946 22258 60958
rect 18386 60846 18398 60898
rect 18450 60846 18462 60898
rect 20638 60786 20690 60798
rect 16818 60734 16830 60786
rect 16882 60734 16894 60786
rect 18722 60734 18734 60786
rect 18786 60734 18798 60786
rect 19506 60734 19518 60786
rect 19570 60734 19582 60786
rect 20638 60722 20690 60734
rect 20862 60786 20914 60798
rect 20862 60722 20914 60734
rect 21086 60786 21138 60798
rect 28466 60734 28478 60786
rect 28530 60734 28542 60786
rect 21086 60722 21138 60734
rect 17502 60674 17554 60686
rect 11778 60622 11790 60674
rect 11842 60622 11854 60674
rect 17502 60610 17554 60622
rect 20078 60674 20130 60686
rect 22642 60622 22654 60674
rect 22706 60622 22718 60674
rect 25666 60622 25678 60674
rect 25730 60622 25742 60674
rect 27794 60622 27806 60674
rect 27858 60622 27870 60674
rect 20078 60610 20130 60622
rect 21310 60562 21362 60574
rect 21310 60498 21362 60510
rect 21758 60562 21810 60574
rect 21758 60498 21810 60510
rect 1344 60394 38640 60428
rect 1344 60342 4478 60394
rect 4530 60342 4582 60394
rect 4634 60342 4686 60394
rect 4738 60342 35198 60394
rect 35250 60342 35302 60394
rect 35354 60342 35406 60394
rect 35458 60342 38640 60394
rect 1344 60308 38640 60342
rect 19070 60226 19122 60238
rect 19070 60162 19122 60174
rect 19742 60226 19794 60238
rect 19742 60162 19794 60174
rect 19854 60226 19906 60238
rect 19854 60162 19906 60174
rect 18510 60002 18562 60014
rect 6066 59950 6078 60002
rect 6130 59950 6142 60002
rect 14802 59950 14814 60002
rect 14866 59950 14878 60002
rect 18510 59938 18562 59950
rect 19294 60002 19346 60014
rect 19294 59938 19346 59950
rect 19630 60002 19682 60014
rect 19630 59938 19682 59950
rect 24782 60002 24834 60014
rect 25330 59950 25342 60002
rect 25394 59950 25406 60002
rect 24782 59938 24834 59950
rect 1710 59890 1762 59902
rect 1710 59826 1762 59838
rect 2494 59890 2546 59902
rect 13470 59890 13522 59902
rect 6738 59838 6750 59890
rect 6802 59838 6814 59890
rect 2494 59826 2546 59838
rect 13470 59826 13522 59838
rect 14478 59890 14530 59902
rect 14478 59826 14530 59838
rect 15934 59890 15986 59902
rect 15934 59826 15986 59838
rect 17390 59890 17442 59902
rect 25118 59890 25170 59902
rect 24882 59838 24894 59890
rect 24946 59838 24958 59890
rect 17390 59826 17442 59838
rect 25118 59826 25170 59838
rect 25790 59890 25842 59902
rect 25790 59826 25842 59838
rect 26238 59890 26290 59902
rect 26238 59826 26290 59838
rect 26574 59890 26626 59902
rect 26574 59826 26626 59838
rect 2046 59778 2098 59790
rect 13582 59778 13634 59790
rect 8978 59726 8990 59778
rect 9042 59726 9054 59778
rect 2046 59714 2098 59726
rect 13582 59714 13634 59726
rect 13694 59778 13746 59790
rect 13694 59714 13746 59726
rect 14366 59778 14418 59790
rect 24446 59778 24498 59790
rect 15810 59726 15822 59778
rect 15874 59726 15886 59778
rect 14366 59714 14418 59726
rect 24446 59714 24498 59726
rect 1344 59610 38640 59644
rect 1344 59558 19838 59610
rect 19890 59558 19942 59610
rect 19994 59558 20046 59610
rect 20098 59558 38640 59610
rect 1344 59524 38640 59558
rect 7982 59442 8034 59454
rect 7982 59378 8034 59390
rect 11118 59442 11170 59454
rect 11118 59378 11170 59390
rect 16270 59442 16322 59454
rect 18162 59390 18174 59442
rect 18226 59390 18238 59442
rect 18834 59390 18846 59442
rect 18898 59390 18910 59442
rect 16270 59378 16322 59390
rect 9662 59330 9714 59342
rect 17502 59330 17554 59342
rect 11442 59278 11454 59330
rect 11506 59278 11518 59330
rect 9662 59266 9714 59278
rect 17502 59266 17554 59278
rect 17726 59330 17778 59342
rect 17726 59266 17778 59278
rect 7870 59218 7922 59230
rect 7870 59154 7922 59166
rect 8206 59218 8258 59230
rect 8206 59154 8258 59166
rect 8430 59218 8482 59230
rect 8430 59154 8482 59166
rect 9438 59218 9490 59230
rect 9438 59154 9490 59166
rect 9774 59218 9826 59230
rect 16830 59218 16882 59230
rect 12226 59166 12238 59218
rect 12290 59166 12302 59218
rect 9774 59154 9826 59166
rect 16830 59154 16882 59166
rect 17614 59218 17666 59230
rect 17614 59154 17666 59166
rect 18510 59218 18562 59230
rect 18510 59154 18562 59166
rect 25902 59106 25954 59118
rect 12898 59054 12910 59106
rect 12962 59054 12974 59106
rect 15026 59054 15038 59106
rect 15090 59054 15102 59106
rect 25902 59042 25954 59054
rect 1344 58826 38640 58860
rect 1344 58774 4478 58826
rect 4530 58774 4582 58826
rect 4634 58774 4686 58826
rect 4738 58774 35198 58826
rect 35250 58774 35302 58826
rect 35354 58774 35406 58826
rect 35458 58774 38640 58826
rect 1344 58740 38640 58774
rect 25902 58658 25954 58670
rect 13682 58606 13694 58658
rect 13746 58606 13758 58658
rect 25902 58594 25954 58606
rect 25566 58546 25618 58558
rect 18162 58494 18174 58546
rect 18226 58494 18238 58546
rect 25566 58482 25618 58494
rect 26910 58546 26962 58558
rect 27570 58494 27582 58546
rect 27634 58494 27646 58546
rect 26910 58482 26962 58494
rect 14254 58434 14306 58446
rect 25678 58434 25730 58446
rect 10098 58382 10110 58434
rect 10162 58382 10174 58434
rect 13570 58382 13582 58434
rect 13634 58382 13646 58434
rect 14018 58382 14030 58434
rect 14082 58382 14094 58434
rect 16258 58382 16270 58434
rect 16322 58382 16334 58434
rect 17490 58382 17502 58434
rect 17554 58382 17566 58434
rect 17826 58382 17838 58434
rect 17890 58382 17902 58434
rect 14254 58370 14306 58382
rect 25678 58370 25730 58382
rect 1710 58322 1762 58334
rect 1710 58258 1762 58270
rect 10334 58322 10386 58334
rect 10334 58258 10386 58270
rect 16718 58322 16770 58334
rect 27246 58322 27298 58334
rect 18386 58270 18398 58322
rect 18450 58270 18462 58322
rect 24770 58270 24782 58322
rect 24834 58270 24846 58322
rect 16718 58258 16770 58270
rect 27246 58258 27298 58270
rect 27470 58322 27522 58334
rect 27470 58258 27522 58270
rect 2046 58210 2098 58222
rect 2046 58146 2098 58158
rect 2494 58210 2546 58222
rect 2494 58146 2546 58158
rect 9774 58210 9826 58222
rect 9774 58146 9826 58158
rect 13470 58210 13522 58222
rect 13470 58146 13522 58158
rect 18958 58210 19010 58222
rect 18958 58146 19010 58158
rect 25118 58210 25170 58222
rect 25118 58146 25170 58158
rect 25566 58210 25618 58222
rect 25566 58146 25618 58158
rect 1344 58042 38640 58076
rect 1344 57990 19838 58042
rect 19890 57990 19942 58042
rect 19994 57990 20046 58042
rect 20098 57990 38640 58042
rect 1344 57956 38640 57990
rect 8094 57874 8146 57886
rect 8094 57810 8146 57822
rect 2046 57762 2098 57774
rect 2046 57698 2098 57710
rect 7758 57762 7810 57774
rect 7758 57698 7810 57710
rect 7870 57762 7922 57774
rect 13022 57762 13074 57774
rect 16158 57762 16210 57774
rect 9874 57710 9886 57762
rect 9938 57710 9950 57762
rect 15810 57710 15822 57762
rect 15874 57710 15886 57762
rect 17602 57710 17614 57762
rect 17666 57710 17678 57762
rect 23650 57710 23662 57762
rect 23714 57710 23726 57762
rect 7870 57698 7922 57710
rect 13022 57698 13074 57710
rect 16158 57698 16210 57710
rect 1710 57650 1762 57662
rect 1710 57586 1762 57598
rect 10222 57650 10274 57662
rect 13346 57598 13358 57650
rect 13410 57598 13422 57650
rect 17714 57598 17726 57650
rect 17778 57598 17790 57650
rect 24434 57598 24446 57650
rect 24498 57598 24510 57650
rect 26002 57598 26014 57650
rect 26066 57598 26078 57650
rect 10222 57586 10274 57598
rect 2494 57538 2546 57550
rect 25678 57538 25730 57550
rect 15026 57486 15038 57538
rect 15090 57486 15102 57538
rect 18610 57486 18622 57538
rect 18674 57486 18686 57538
rect 21522 57486 21534 57538
rect 21586 57486 21598 57538
rect 26002 57535 26014 57538
rect 2494 57474 2546 57486
rect 25678 57474 25730 57486
rect 25793 57489 26014 57535
rect 13358 57426 13410 57438
rect 13358 57362 13410 57374
rect 16382 57426 16434 57438
rect 16706 57374 16718 57426
rect 16770 57374 16782 57426
rect 25666 57374 25678 57426
rect 25730 57423 25742 57426
rect 25793 57423 25839 57489
rect 26002 57486 26014 57489
rect 26066 57486 26078 57538
rect 28466 57486 28478 57538
rect 28530 57486 28542 57538
rect 25730 57377 25839 57423
rect 25730 57374 25742 57377
rect 16382 57362 16434 57374
rect 1344 57258 38640 57292
rect 1344 57206 4478 57258
rect 4530 57206 4582 57258
rect 4634 57206 4686 57258
rect 4738 57206 35198 57258
rect 35250 57206 35302 57258
rect 35354 57206 35406 57258
rect 35458 57206 38640 57258
rect 1344 57172 38640 57206
rect 25342 57090 25394 57102
rect 28030 57090 28082 57102
rect 13682 57038 13694 57090
rect 13746 57038 13758 57090
rect 27234 57038 27246 57090
rect 27298 57038 27310 57090
rect 25342 57026 25394 57038
rect 28030 57026 28082 57038
rect 17502 56978 17554 56990
rect 17502 56914 17554 56926
rect 18062 56978 18114 56990
rect 21410 56926 21422 56978
rect 21474 56926 21486 56978
rect 18062 56914 18114 56926
rect 22654 56866 22706 56878
rect 13458 56814 13470 56866
rect 13522 56814 13534 56866
rect 14018 56814 14030 56866
rect 14082 56814 14094 56866
rect 16706 56814 16718 56866
rect 16770 56814 16782 56866
rect 17602 56814 17614 56866
rect 17666 56814 17678 56866
rect 21858 56814 21870 56866
rect 21922 56814 21934 56866
rect 22654 56802 22706 56814
rect 23662 56866 23714 56878
rect 23662 56802 23714 56814
rect 24446 56866 24498 56878
rect 25118 56866 25170 56878
rect 27358 56866 27410 56878
rect 24658 56814 24670 56866
rect 24722 56814 24734 56866
rect 26898 56814 26910 56866
rect 26962 56814 26974 56866
rect 24446 56802 24498 56814
rect 25118 56802 25170 56814
rect 27358 56802 27410 56814
rect 28254 56866 28306 56878
rect 28254 56802 28306 56814
rect 28366 56866 28418 56878
rect 28366 56802 28418 56814
rect 1710 56754 1762 56766
rect 1710 56690 1762 56702
rect 7422 56754 7474 56766
rect 7422 56690 7474 56702
rect 7758 56754 7810 56766
rect 7758 56690 7810 56702
rect 7982 56754 8034 56766
rect 7982 56690 8034 56702
rect 8318 56754 8370 56766
rect 8318 56690 8370 56702
rect 8542 56754 8594 56766
rect 14254 56754 14306 56766
rect 12338 56702 12350 56754
rect 12402 56702 12414 56754
rect 8542 56690 8594 56702
rect 14254 56690 14306 56702
rect 15598 56754 15650 56766
rect 15598 56690 15650 56702
rect 16270 56754 16322 56766
rect 16270 56690 16322 56702
rect 22318 56754 22370 56766
rect 22318 56690 22370 56702
rect 24782 56754 24834 56766
rect 24782 56690 24834 56702
rect 27918 56754 27970 56766
rect 27918 56690 27970 56702
rect 2046 56642 2098 56654
rect 2046 56578 2098 56590
rect 2494 56642 2546 56654
rect 2494 56578 2546 56590
rect 7534 56642 7586 56654
rect 7534 56578 7586 56590
rect 8094 56642 8146 56654
rect 8094 56578 8146 56590
rect 12014 56642 12066 56654
rect 12014 56578 12066 56590
rect 13470 56642 13522 56654
rect 13470 56578 13522 56590
rect 15486 56642 15538 56654
rect 15486 56578 15538 56590
rect 17166 56642 17218 56654
rect 17166 56578 17218 56590
rect 17390 56642 17442 56654
rect 17390 56578 17442 56590
rect 22766 56642 22818 56654
rect 22766 56578 22818 56590
rect 23102 56642 23154 56654
rect 25666 56590 25678 56642
rect 25730 56590 25742 56642
rect 23102 56578 23154 56590
rect 1344 56474 38640 56508
rect 1344 56422 19838 56474
rect 19890 56422 19942 56474
rect 19994 56422 20046 56474
rect 20098 56422 38640 56474
rect 1344 56388 38640 56422
rect 2046 56306 2098 56318
rect 2046 56242 2098 56254
rect 17614 56306 17666 56318
rect 17614 56242 17666 56254
rect 10110 56194 10162 56206
rect 10110 56130 10162 56142
rect 24558 56194 24610 56206
rect 27794 56142 27806 56194
rect 27858 56142 27870 56194
rect 24558 56130 24610 56142
rect 1710 56082 1762 56094
rect 9438 56082 9490 56094
rect 5954 56030 5966 56082
rect 6018 56030 6030 56082
rect 1710 56018 1762 56030
rect 9438 56018 9490 56030
rect 9774 56082 9826 56094
rect 17502 56082 17554 56094
rect 16594 56030 16606 56082
rect 16658 56030 16670 56082
rect 9774 56018 9826 56030
rect 17502 56018 17554 56030
rect 17838 56082 17890 56094
rect 18398 56082 18450 56094
rect 24446 56082 24498 56094
rect 18050 56030 18062 56082
rect 18114 56030 18126 56082
rect 21746 56030 21758 56082
rect 21810 56030 21822 56082
rect 17838 56018 17890 56030
rect 18398 56018 18450 56030
rect 24446 56018 24498 56030
rect 24782 56082 24834 56094
rect 25566 56082 25618 56094
rect 25330 56030 25342 56082
rect 25394 56030 25406 56082
rect 24782 56018 24834 56030
rect 25566 56018 25618 56030
rect 25902 56082 25954 56094
rect 27122 56030 27134 56082
rect 27186 56030 27198 56082
rect 25902 56018 25954 56030
rect 2494 55970 2546 55982
rect 8766 55970 8818 55982
rect 6626 55918 6638 55970
rect 6690 55918 6702 55970
rect 2494 55906 2546 55918
rect 8766 55906 8818 55918
rect 9662 55970 9714 55982
rect 17726 55970 17778 55982
rect 12002 55918 12014 55970
rect 12066 55918 12078 55970
rect 9662 55906 9714 55918
rect 17726 55906 17778 55918
rect 18958 55970 19010 55982
rect 18958 55906 19010 55918
rect 21086 55970 21138 55982
rect 21410 55918 21422 55970
rect 21474 55918 21486 55970
rect 29922 55918 29934 55970
rect 29986 55918 29998 55970
rect 21086 55906 21138 55918
rect 25790 55858 25842 55870
rect 25790 55794 25842 55806
rect 1344 55690 38640 55724
rect 1344 55638 4478 55690
rect 4530 55638 4582 55690
rect 4634 55638 4686 55690
rect 4738 55638 35198 55690
rect 35250 55638 35302 55690
rect 35354 55638 35406 55690
rect 35458 55638 38640 55690
rect 1344 55604 38640 55638
rect 22194 55470 22206 55522
rect 22258 55470 22270 55522
rect 11566 55410 11618 55422
rect 29262 55410 29314 55422
rect 9090 55358 9102 55410
rect 9154 55358 9166 55410
rect 17266 55358 17278 55410
rect 17330 55358 17342 55410
rect 21970 55358 21982 55410
rect 22034 55358 22046 55410
rect 27682 55358 27694 55410
rect 27746 55358 27758 55410
rect 11566 55346 11618 55358
rect 29262 55346 29314 55358
rect 9326 55298 9378 55310
rect 6290 55246 6302 55298
rect 6354 55246 6366 55298
rect 9326 55234 9378 55246
rect 9662 55298 9714 55310
rect 26910 55298 26962 55310
rect 10546 55246 10558 55298
rect 10610 55246 10622 55298
rect 15026 55246 15038 55298
rect 15090 55246 15102 55298
rect 15586 55246 15598 55298
rect 15650 55246 15662 55298
rect 18386 55246 18398 55298
rect 18450 55246 18462 55298
rect 22082 55246 22094 55298
rect 22146 55246 22158 55298
rect 26338 55246 26350 55298
rect 26402 55246 26414 55298
rect 9662 55234 9714 55246
rect 26910 55234 26962 55246
rect 29038 55298 29090 55310
rect 29038 55234 29090 55246
rect 29374 55298 29426 55310
rect 29374 55234 29426 55246
rect 29598 55298 29650 55310
rect 29598 55234 29650 55246
rect 1710 55186 1762 55198
rect 2494 55186 2546 55198
rect 10334 55186 10386 55198
rect 2034 55134 2046 55186
rect 2098 55134 2110 55186
rect 6962 55134 6974 55186
rect 7026 55134 7038 55186
rect 1710 55122 1762 55134
rect 2494 55122 2546 55134
rect 10334 55122 10386 55134
rect 11902 55186 11954 55198
rect 19182 55186 19234 55198
rect 12898 55134 12910 55186
rect 12962 55134 12974 55186
rect 17154 55134 17166 55186
rect 17218 55134 17230 55186
rect 18162 55134 18174 55186
rect 18226 55134 18238 55186
rect 11902 55122 11954 55134
rect 19182 55122 19234 55134
rect 25342 55186 25394 55198
rect 25342 55122 25394 55134
rect 27358 55186 27410 55198
rect 27358 55122 27410 55134
rect 9550 55074 9602 55086
rect 9550 55010 9602 55022
rect 11006 55074 11058 55086
rect 11006 55010 11058 55022
rect 12238 55074 12290 55086
rect 12238 55010 12290 55022
rect 12574 55074 12626 55086
rect 12574 55010 12626 55022
rect 15262 55074 15314 55086
rect 15262 55010 15314 55022
rect 19294 55074 19346 55086
rect 19294 55010 19346 55022
rect 1344 54906 38640 54940
rect 1344 54854 19838 54906
rect 19890 54854 19942 54906
rect 19994 54854 20046 54906
rect 20098 54854 38640 54906
rect 1344 54820 38640 54854
rect 8094 54738 8146 54750
rect 8094 54674 8146 54686
rect 9102 54738 9154 54750
rect 10110 54738 10162 54750
rect 9762 54686 9774 54738
rect 9826 54686 9838 54738
rect 14914 54686 14926 54738
rect 14978 54686 14990 54738
rect 9102 54674 9154 54686
rect 10110 54674 10162 54686
rect 7758 54626 7810 54638
rect 7758 54562 7810 54574
rect 7870 54626 7922 54638
rect 7870 54562 7922 54574
rect 8878 54626 8930 54638
rect 25454 54626 25506 54638
rect 12674 54574 12686 54626
rect 12738 54574 12750 54626
rect 16594 54574 16606 54626
rect 16658 54574 16670 54626
rect 18834 54574 18846 54626
rect 18898 54574 18910 54626
rect 27794 54574 27806 54626
rect 27858 54574 27870 54626
rect 8878 54562 8930 54574
rect 25454 54562 25506 54574
rect 8766 54514 8818 54526
rect 12002 54462 12014 54514
rect 12066 54462 12078 54514
rect 17602 54462 17614 54514
rect 17666 54462 17678 54514
rect 20066 54462 20078 54514
rect 20130 54462 20142 54514
rect 27122 54462 27134 54514
rect 27186 54462 27198 54514
rect 35970 54462 35982 54514
rect 36034 54462 36046 54514
rect 8766 54450 8818 54462
rect 18174 54402 18226 54414
rect 17714 54350 17726 54402
rect 17778 54350 17790 54402
rect 18174 54338 18226 54350
rect 18734 54402 18786 54414
rect 18734 54338 18786 54350
rect 20750 54402 20802 54414
rect 20750 54338 20802 54350
rect 25342 54402 25394 54414
rect 29922 54350 29934 54402
rect 29986 54350 29998 54402
rect 25342 54338 25394 54350
rect 16046 54290 16098 54302
rect 16046 54226 16098 54238
rect 25230 54290 25282 54302
rect 25230 54226 25282 54238
rect 37998 54290 38050 54302
rect 37998 54226 38050 54238
rect 1344 54122 38640 54156
rect 1344 54070 4478 54122
rect 4530 54070 4582 54122
rect 4634 54070 4686 54122
rect 4738 54070 35198 54122
rect 35250 54070 35302 54122
rect 35354 54070 35406 54122
rect 35458 54070 38640 54122
rect 1344 54036 38640 54070
rect 27582 53954 27634 53966
rect 27582 53890 27634 53902
rect 19406 53842 19458 53854
rect 27234 53790 27246 53842
rect 27298 53790 27310 53842
rect 19406 53778 19458 53790
rect 19182 53730 19234 53742
rect 16930 53678 16942 53730
rect 16994 53678 17006 53730
rect 17378 53678 17390 53730
rect 17442 53678 17454 53730
rect 19182 53666 19234 53678
rect 21310 53730 21362 53742
rect 21310 53666 21362 53678
rect 21982 53730 22034 53742
rect 22418 53678 22430 53730
rect 22482 53678 22494 53730
rect 24434 53678 24446 53730
rect 24498 53678 24510 53730
rect 26898 53678 26910 53730
rect 26962 53678 26974 53730
rect 21982 53666 22034 53678
rect 16382 53618 16434 53630
rect 16382 53554 16434 53566
rect 17838 53618 17890 53630
rect 17838 53554 17890 53566
rect 21534 53618 21586 53630
rect 25006 53618 25058 53630
rect 22530 53566 22542 53618
rect 22594 53566 22606 53618
rect 21534 53554 21586 53566
rect 25006 53554 25058 53566
rect 1710 53506 1762 53518
rect 2494 53506 2546 53518
rect 2034 53454 2046 53506
rect 2098 53454 2110 53506
rect 1710 53442 1762 53454
rect 2494 53442 2546 53454
rect 15934 53506 15986 53518
rect 15934 53442 15986 53454
rect 19518 53506 19570 53518
rect 19518 53442 19570 53454
rect 19742 53506 19794 53518
rect 19742 53442 19794 53454
rect 21758 53506 21810 53518
rect 26798 53506 26850 53518
rect 23986 53454 23998 53506
rect 24050 53454 24062 53506
rect 21758 53442 21810 53454
rect 26798 53442 26850 53454
rect 27358 53506 27410 53518
rect 27358 53442 27410 53454
rect 1344 53338 38640 53372
rect 1344 53286 19838 53338
rect 19890 53286 19942 53338
rect 19994 53286 20046 53338
rect 20098 53286 38640 53338
rect 1344 53252 38640 53286
rect 10334 53170 10386 53182
rect 17490 53118 17502 53170
rect 17554 53118 17566 53170
rect 17714 53118 17726 53170
rect 17778 53118 17790 53170
rect 10334 53106 10386 53118
rect 15262 53058 15314 53070
rect 24670 53058 24722 53070
rect 18722 53006 18734 53058
rect 18786 53006 18798 53058
rect 21298 53006 21310 53058
rect 21362 53006 21374 53058
rect 22978 53006 22990 53058
rect 23042 53006 23054 53058
rect 15262 52994 15314 53006
rect 24670 52994 24722 53006
rect 14802 52894 14814 52946
rect 14866 52894 14878 52946
rect 15026 52894 15038 52946
rect 15090 52894 15102 52946
rect 16594 52894 16606 52946
rect 16658 52894 16670 52946
rect 17378 52894 17390 52946
rect 17442 52894 17454 52946
rect 18498 52894 18510 52946
rect 18562 52894 18574 52946
rect 19394 52894 19406 52946
rect 19458 52894 19470 52946
rect 19730 52894 19742 52946
rect 19794 52894 19806 52946
rect 21858 52894 21870 52946
rect 21922 52894 21934 52946
rect 22306 52894 22318 52946
rect 22370 52894 22382 52946
rect 24098 52894 24110 52946
rect 24162 52894 24174 52946
rect 25890 52894 25902 52946
rect 25954 52894 25966 52946
rect 33058 52894 33070 52946
rect 33122 52894 33134 52946
rect 10222 52834 10274 52846
rect 10222 52770 10274 52782
rect 16270 52834 16322 52846
rect 20962 52782 20974 52834
rect 21026 52782 21038 52834
rect 22194 52782 22206 52834
rect 22258 52782 22270 52834
rect 24210 52782 24222 52834
rect 24274 52782 24286 52834
rect 26562 52782 26574 52834
rect 26626 52782 26638 52834
rect 28690 52782 28702 52834
rect 28754 52782 28766 52834
rect 33842 52782 33854 52834
rect 33906 52782 33918 52834
rect 35970 52782 35982 52834
rect 36034 52782 36046 52834
rect 16270 52770 16322 52782
rect 15374 52722 15426 52734
rect 15374 52658 15426 52670
rect 1344 52554 38640 52588
rect 1344 52502 4478 52554
rect 4530 52502 4582 52554
rect 4634 52502 4686 52554
rect 4738 52502 35198 52554
rect 35250 52502 35302 52554
rect 35354 52502 35406 52554
rect 35458 52502 38640 52554
rect 1344 52468 38640 52502
rect 12462 52386 12514 52398
rect 12462 52322 12514 52334
rect 26574 52386 26626 52398
rect 26574 52322 26626 52334
rect 26686 52386 26738 52398
rect 26686 52322 26738 52334
rect 26910 52386 26962 52398
rect 27346 52334 27358 52386
rect 27410 52383 27422 52386
rect 27570 52383 27582 52386
rect 27410 52337 27582 52383
rect 27410 52334 27422 52337
rect 27570 52334 27582 52337
rect 27634 52334 27646 52386
rect 26910 52322 26962 52334
rect 27582 52274 27634 52286
rect 11778 52222 11790 52274
rect 11842 52222 11854 52274
rect 15698 52222 15710 52274
rect 15762 52222 15774 52274
rect 16706 52222 16718 52274
rect 16770 52222 16782 52274
rect 18386 52222 18398 52274
rect 18450 52222 18462 52274
rect 27582 52210 27634 52222
rect 1710 52162 1762 52174
rect 1710 52098 1762 52110
rect 2494 52162 2546 52174
rect 2494 52098 2546 52110
rect 11454 52162 11506 52174
rect 20190 52162 20242 52174
rect 33742 52162 33794 52174
rect 12114 52110 12126 52162
rect 12178 52110 12190 52162
rect 15474 52110 15486 52162
rect 15538 52110 15550 52162
rect 18162 52110 18174 52162
rect 18226 52110 18238 52162
rect 21858 52110 21870 52162
rect 21922 52110 21934 52162
rect 23874 52110 23886 52162
rect 23938 52110 23950 52162
rect 27122 52110 27134 52162
rect 27186 52110 27198 52162
rect 11454 52098 11506 52110
rect 20190 52098 20242 52110
rect 33742 52098 33794 52110
rect 2046 52050 2098 52062
rect 12910 52050 12962 52062
rect 24446 52050 24498 52062
rect 12674 51998 12686 52050
rect 12738 51998 12750 52050
rect 17938 51998 17950 52050
rect 18002 51998 18014 52050
rect 18610 51998 18622 52050
rect 18674 51998 18686 52050
rect 21970 51998 21982 52050
rect 22034 51998 22046 52050
rect 2046 51986 2098 51998
rect 12910 51986 12962 51998
rect 24446 51986 24498 51998
rect 34078 52050 34130 52062
rect 34078 51986 34130 51998
rect 11678 51938 11730 51950
rect 12450 51886 12462 51938
rect 12514 51886 12526 51938
rect 23426 51886 23438 51938
rect 23490 51886 23502 51938
rect 11678 51874 11730 51886
rect 1344 51770 38640 51804
rect 1344 51718 19838 51770
rect 19890 51718 19942 51770
rect 19994 51718 20046 51770
rect 20098 51718 38640 51770
rect 1344 51684 38640 51718
rect 10222 51602 10274 51614
rect 10222 51538 10274 51550
rect 15598 51602 15650 51614
rect 15598 51538 15650 51550
rect 16046 51602 16098 51614
rect 23314 51550 23326 51602
rect 23378 51550 23390 51602
rect 26562 51550 26574 51602
rect 26626 51550 26638 51602
rect 16046 51538 16098 51550
rect 2046 51490 2098 51502
rect 16606 51490 16658 51502
rect 25678 51490 25730 51502
rect 9538 51438 9550 51490
rect 9602 51438 9614 51490
rect 10546 51438 10558 51490
rect 10610 51438 10622 51490
rect 12450 51438 12462 51490
rect 12514 51438 12526 51490
rect 17938 51438 17950 51490
rect 18002 51438 18014 51490
rect 19170 51438 19182 51490
rect 19234 51438 19246 51490
rect 23090 51438 23102 51490
rect 23154 51438 23166 51490
rect 24098 51438 24110 51490
rect 24162 51438 24174 51490
rect 2046 51426 2098 51438
rect 16606 51426 16658 51438
rect 25678 51426 25730 51438
rect 26910 51490 26962 51502
rect 26910 51426 26962 51438
rect 1710 51378 1762 51390
rect 15710 51378 15762 51390
rect 24670 51378 24722 51390
rect 6178 51326 6190 51378
rect 6242 51326 6254 51378
rect 9762 51326 9774 51378
rect 9826 51326 9838 51378
rect 11778 51326 11790 51378
rect 11842 51326 11854 51378
rect 18050 51326 18062 51378
rect 18114 51326 18126 51378
rect 19058 51326 19070 51378
rect 19122 51326 19134 51378
rect 22418 51326 22430 51378
rect 22482 51326 22494 51378
rect 22978 51326 22990 51378
rect 23042 51326 23054 51378
rect 23762 51326 23774 51378
rect 23826 51326 23838 51378
rect 1710 51314 1762 51326
rect 15710 51314 15762 51326
rect 24670 51314 24722 51326
rect 26238 51378 26290 51390
rect 37762 51326 37774 51378
rect 37826 51326 37838 51378
rect 26238 51314 26290 51326
rect 2494 51266 2546 51278
rect 27358 51266 27410 51278
rect 6850 51214 6862 51266
rect 6914 51214 6926 51266
rect 8978 51214 8990 51266
rect 9042 51214 9054 51266
rect 14578 51214 14590 51266
rect 14642 51214 14654 51266
rect 18610 51214 18622 51266
rect 18674 51214 18686 51266
rect 2494 51202 2546 51214
rect 27358 51202 27410 51214
rect 27806 51266 27858 51278
rect 27806 51202 27858 51214
rect 27346 51102 27358 51154
rect 27410 51151 27422 51154
rect 27794 51151 27806 51154
rect 27410 51105 27806 51151
rect 27410 51102 27422 51105
rect 27794 51102 27806 51105
rect 27858 51102 27870 51154
rect 36754 51102 36766 51154
rect 36818 51102 36830 51154
rect 1344 50986 38640 51020
rect 1344 50934 4478 50986
rect 4530 50934 4582 50986
rect 4634 50934 4686 50986
rect 4738 50934 35198 50986
rect 35250 50934 35302 50986
rect 35354 50934 35406 50986
rect 35458 50934 38640 50986
rect 1344 50900 38640 50934
rect 11454 50818 11506 50830
rect 12338 50766 12350 50818
rect 12402 50766 12414 50818
rect 32946 50766 32958 50818
rect 33010 50766 33022 50818
rect 11454 50754 11506 50766
rect 17614 50706 17666 50718
rect 11666 50654 11678 50706
rect 11730 50654 11742 50706
rect 17614 50642 17666 50654
rect 17726 50706 17778 50718
rect 33518 50706 33570 50718
rect 19730 50654 19742 50706
rect 19794 50654 19806 50706
rect 17726 50642 17778 50654
rect 33518 50642 33570 50654
rect 7422 50594 7474 50606
rect 9438 50594 9490 50606
rect 33294 50594 33346 50606
rect 8530 50542 8542 50594
rect 8594 50542 8606 50594
rect 10546 50542 10558 50594
rect 10610 50542 10622 50594
rect 12114 50542 12126 50594
rect 12178 50542 12190 50594
rect 12674 50542 12686 50594
rect 12738 50542 12750 50594
rect 15810 50542 15822 50594
rect 15874 50542 15886 50594
rect 20738 50542 20750 50594
rect 20802 50542 20814 50594
rect 26562 50542 26574 50594
rect 26626 50542 26638 50594
rect 7422 50530 7474 50542
rect 9438 50530 9490 50542
rect 33294 50530 33346 50542
rect 1710 50482 1762 50494
rect 1710 50418 1762 50430
rect 2382 50482 2434 50494
rect 2382 50418 2434 50430
rect 2718 50482 2770 50494
rect 2718 50418 2770 50430
rect 3166 50482 3218 50494
rect 3166 50418 3218 50430
rect 7758 50482 7810 50494
rect 9550 50482 9602 50494
rect 8306 50430 8318 50482
rect 8370 50430 8382 50482
rect 7758 50418 7810 50430
rect 9550 50418 9602 50430
rect 9774 50482 9826 50494
rect 9774 50418 9826 50430
rect 9998 50482 10050 50494
rect 9998 50418 10050 50430
rect 12910 50482 12962 50494
rect 12910 50418 12962 50430
rect 15150 50482 15202 50494
rect 15150 50418 15202 50430
rect 15262 50482 15314 50494
rect 15262 50418 15314 50430
rect 16382 50482 16434 50494
rect 27022 50482 27074 50494
rect 20626 50430 20638 50482
rect 20690 50430 20702 50482
rect 22978 50430 22990 50482
rect 23042 50430 23054 50482
rect 16382 50418 16434 50430
rect 27022 50418 27074 50430
rect 2046 50370 2098 50382
rect 2046 50306 2098 50318
rect 7646 50370 7698 50382
rect 11678 50370 11730 50382
rect 10322 50318 10334 50370
rect 10386 50318 10398 50370
rect 7646 50306 7698 50318
rect 11678 50306 11730 50318
rect 12798 50370 12850 50382
rect 12798 50306 12850 50318
rect 1344 50202 38640 50236
rect 1344 50150 19838 50202
rect 19890 50150 19942 50202
rect 19994 50150 20046 50202
rect 20098 50150 38640 50202
rect 1344 50116 38640 50150
rect 2494 50034 2546 50046
rect 2494 49970 2546 49982
rect 10446 50034 10498 50046
rect 15586 49982 15598 50034
rect 15650 49982 15662 50034
rect 23874 49982 23886 50034
rect 23938 49982 23950 50034
rect 10446 49970 10498 49982
rect 2046 49922 2098 49934
rect 2046 49858 2098 49870
rect 9550 49922 9602 49934
rect 9550 49858 9602 49870
rect 9662 49922 9714 49934
rect 9662 49858 9714 49870
rect 11230 49922 11282 49934
rect 12674 49870 12686 49922
rect 12738 49870 12750 49922
rect 15362 49870 15374 49922
rect 15426 49870 15438 49922
rect 15922 49870 15934 49922
rect 15986 49870 15998 49922
rect 19058 49870 19070 49922
rect 19122 49870 19134 49922
rect 21074 49870 21086 49922
rect 21138 49870 21150 49922
rect 22642 49870 22654 49922
rect 22706 49870 22718 49922
rect 23314 49870 23326 49922
rect 23378 49870 23390 49922
rect 23538 49870 23550 49922
rect 23602 49870 23614 49922
rect 11230 49858 11282 49870
rect 1710 49810 1762 49822
rect 9886 49810 9938 49822
rect 5282 49758 5294 49810
rect 5346 49758 5358 49810
rect 1710 49746 1762 49758
rect 9886 49746 9938 49758
rect 10222 49810 10274 49822
rect 22094 49810 22146 49822
rect 11554 49758 11566 49810
rect 11618 49758 11630 49810
rect 11890 49758 11902 49810
rect 11954 49758 11966 49810
rect 16258 49758 16270 49810
rect 16322 49758 16334 49810
rect 17602 49758 17614 49810
rect 17666 49758 17678 49810
rect 18386 49758 18398 49810
rect 18450 49758 18462 49810
rect 21634 49758 21646 49810
rect 21698 49758 21710 49810
rect 10222 49746 10274 49758
rect 22094 49746 22146 49758
rect 23998 49810 24050 49822
rect 31154 49758 31166 49810
rect 31218 49758 31230 49810
rect 34850 49758 34862 49810
rect 34914 49758 34926 49810
rect 23998 49746 24050 49758
rect 2942 49698 2994 49710
rect 11342 49698 11394 49710
rect 5954 49646 5966 49698
rect 6018 49646 6030 49698
rect 8194 49646 8206 49698
rect 8258 49646 8270 49698
rect 14802 49646 14814 49698
rect 14866 49646 14878 49698
rect 18498 49646 18510 49698
rect 18562 49646 18574 49698
rect 22194 49646 22206 49698
rect 22258 49646 22270 49698
rect 28354 49646 28366 49698
rect 28418 49646 28430 49698
rect 30482 49646 30494 49698
rect 30546 49646 30558 49698
rect 35634 49646 35646 49698
rect 35698 49646 35710 49698
rect 37762 49646 37774 49698
rect 37826 49646 37838 49698
rect 2942 49634 2994 49646
rect 11342 49634 11394 49646
rect 10558 49586 10610 49598
rect 10558 49522 10610 49534
rect 1344 49418 38640 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 38640 49418
rect 1344 49332 38640 49366
rect 9886 49138 9938 49150
rect 32398 49138 32450 49150
rect 18050 49086 18062 49138
rect 18114 49086 18126 49138
rect 22754 49086 22766 49138
rect 22818 49086 22830 49138
rect 24210 49086 24222 49138
rect 24274 49086 24286 49138
rect 29138 49086 29150 49138
rect 29202 49086 29214 49138
rect 9886 49074 9938 49086
rect 32398 49074 32450 49086
rect 33406 49138 33458 49150
rect 35634 49086 35646 49138
rect 35698 49086 35710 49138
rect 33406 49074 33458 49086
rect 7198 49026 7250 49038
rect 7198 48962 7250 48974
rect 7534 49026 7586 49038
rect 7534 48962 7586 48974
rect 8206 49026 8258 49038
rect 8206 48962 8258 48974
rect 8654 49026 8706 49038
rect 8654 48962 8706 48974
rect 15486 49026 15538 49038
rect 15486 48962 15538 48974
rect 15710 49026 15762 49038
rect 15710 48962 15762 48974
rect 15934 49026 15986 49038
rect 20414 49026 20466 49038
rect 17826 48974 17838 49026
rect 17890 48974 17902 49026
rect 19170 48974 19182 49026
rect 19234 48974 19246 49026
rect 15934 48962 15986 48974
rect 20414 48962 20466 48974
rect 22318 49026 22370 49038
rect 33294 49026 33346 49038
rect 35982 49026 36034 49038
rect 23090 48974 23102 49026
rect 23154 48974 23166 49026
rect 23650 48974 23662 49026
rect 23714 48974 23726 49026
rect 27010 48974 27022 49026
rect 27074 48974 27086 49026
rect 31938 48974 31950 49026
rect 32002 48974 32014 49026
rect 35074 48974 35086 49026
rect 35138 48974 35150 49026
rect 35410 48974 35422 49026
rect 35474 48974 35486 49026
rect 22318 48962 22370 48974
rect 33294 48962 33346 48974
rect 35982 48962 36034 48974
rect 1710 48914 1762 48926
rect 1710 48850 1762 48862
rect 2046 48914 2098 48926
rect 2046 48850 2098 48862
rect 6638 48914 6690 48926
rect 6638 48850 6690 48862
rect 8878 48914 8930 48926
rect 8878 48850 8930 48862
rect 19966 48914 20018 48926
rect 34414 48914 34466 48926
rect 22754 48862 22766 48914
rect 22818 48862 22830 48914
rect 26338 48862 26350 48914
rect 26402 48862 26414 48914
rect 31266 48862 31278 48914
rect 31330 48862 31342 48914
rect 19966 48850 20018 48862
rect 34414 48850 34466 48862
rect 2494 48802 2546 48814
rect 2494 48738 2546 48750
rect 6750 48802 6802 48814
rect 6750 48738 6802 48750
rect 6974 48802 7026 48814
rect 6974 48738 7026 48750
rect 7310 48802 7362 48814
rect 7310 48738 7362 48750
rect 8430 48802 8482 48814
rect 21758 48802 21810 48814
rect 16258 48750 16270 48802
rect 16322 48750 16334 48802
rect 8430 48738 8482 48750
rect 21758 48738 21810 48750
rect 32958 48802 33010 48814
rect 32958 48738 33010 48750
rect 33518 48802 33570 48814
rect 33518 48738 33570 48750
rect 33742 48802 33794 48814
rect 33742 48738 33794 48750
rect 34638 48802 34690 48814
rect 34638 48738 34690 48750
rect 34750 48802 34802 48814
rect 34750 48738 34802 48750
rect 34862 48802 34914 48814
rect 34862 48738 34914 48750
rect 35646 48802 35698 48814
rect 35646 48738 35698 48750
rect 35870 48802 35922 48814
rect 35870 48738 35922 48750
rect 1344 48634 38640 48668
rect 1344 48582 19838 48634
rect 19890 48582 19942 48634
rect 19994 48582 20046 48634
rect 20098 48582 38640 48634
rect 1344 48548 38640 48582
rect 6638 48466 6690 48478
rect 6638 48402 6690 48414
rect 6862 48466 6914 48478
rect 6862 48402 6914 48414
rect 7646 48466 7698 48478
rect 7646 48402 7698 48414
rect 11118 48466 11170 48478
rect 11118 48402 11170 48414
rect 18398 48466 18450 48478
rect 18398 48402 18450 48414
rect 18622 48466 18674 48478
rect 21422 48466 21474 48478
rect 20850 48414 20862 48466
rect 20914 48414 20926 48466
rect 18622 48402 18674 48414
rect 21422 48402 21474 48414
rect 26126 48466 26178 48478
rect 26126 48402 26178 48414
rect 31278 48466 31330 48478
rect 31278 48402 31330 48414
rect 32510 48466 32562 48478
rect 32510 48402 32562 48414
rect 2046 48354 2098 48366
rect 2046 48290 2098 48302
rect 6974 48354 7026 48366
rect 18174 48354 18226 48366
rect 7298 48302 7310 48354
rect 7362 48302 7374 48354
rect 6974 48290 7026 48302
rect 18174 48290 18226 48302
rect 21198 48354 21250 48366
rect 21198 48290 21250 48302
rect 22206 48354 22258 48366
rect 22206 48290 22258 48302
rect 23998 48354 24050 48366
rect 23998 48290 24050 48302
rect 24110 48354 24162 48366
rect 24110 48290 24162 48302
rect 25566 48354 25618 48366
rect 25566 48290 25618 48302
rect 26798 48354 26850 48366
rect 27470 48354 27522 48366
rect 27122 48302 27134 48354
rect 27186 48302 27198 48354
rect 26798 48290 26850 48302
rect 27470 48290 27522 48302
rect 32174 48354 32226 48366
rect 32174 48290 32226 48302
rect 32286 48354 32338 48366
rect 32286 48290 32338 48302
rect 33630 48354 33682 48366
rect 33630 48290 33682 48302
rect 1710 48242 1762 48254
rect 11566 48242 11618 48254
rect 11330 48190 11342 48242
rect 11394 48190 11406 48242
rect 1710 48178 1762 48190
rect 11566 48178 11618 48190
rect 11902 48242 11954 48254
rect 11902 48178 11954 48190
rect 18734 48242 18786 48254
rect 18734 48178 18786 48190
rect 20302 48242 20354 48254
rect 20302 48178 20354 48190
rect 21534 48242 21586 48254
rect 21534 48178 21586 48190
rect 21646 48242 21698 48254
rect 22318 48242 22370 48254
rect 21858 48190 21870 48242
rect 21922 48190 21934 48242
rect 21646 48178 21698 48190
rect 22318 48178 22370 48190
rect 22542 48242 22594 48254
rect 22542 48178 22594 48190
rect 22766 48242 22818 48254
rect 22766 48178 22818 48190
rect 24222 48242 24274 48254
rect 26462 48242 26514 48254
rect 24658 48190 24670 48242
rect 24722 48190 24734 48242
rect 25330 48190 25342 48242
rect 25394 48190 25406 48242
rect 31826 48190 31838 48242
rect 31890 48190 31902 48242
rect 33282 48190 33294 48242
rect 33346 48190 33358 48242
rect 38210 48190 38222 48242
rect 38274 48190 38286 48242
rect 24222 48178 24274 48190
rect 26462 48178 26514 48190
rect 2494 48130 2546 48142
rect 2494 48066 2546 48078
rect 18510 48130 18562 48142
rect 18510 48066 18562 48078
rect 28030 48130 28082 48142
rect 33170 48078 33182 48130
rect 33234 48078 33246 48130
rect 34850 48078 34862 48130
rect 34914 48078 34926 48130
rect 36866 48078 36878 48130
rect 36930 48078 36942 48130
rect 28030 48066 28082 48078
rect 20526 48018 20578 48030
rect 11330 47966 11342 48018
rect 11394 47966 11406 48018
rect 23202 47966 23214 48018
rect 23266 47966 23278 48018
rect 20526 47954 20578 47966
rect 1344 47850 38640 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 38640 47850
rect 1344 47764 38640 47798
rect 20750 47682 20802 47694
rect 33730 47630 33742 47682
rect 33794 47630 33806 47682
rect 20750 47618 20802 47630
rect 25006 47570 25058 47582
rect 25006 47506 25058 47518
rect 25342 47570 25394 47582
rect 25342 47506 25394 47518
rect 26574 47570 26626 47582
rect 26574 47506 26626 47518
rect 27246 47570 27298 47582
rect 27246 47506 27298 47518
rect 29934 47570 29986 47582
rect 29934 47506 29986 47518
rect 31838 47570 31890 47582
rect 31838 47506 31890 47518
rect 7982 47458 8034 47470
rect 7982 47394 8034 47406
rect 18286 47458 18338 47470
rect 18286 47394 18338 47406
rect 30158 47458 30210 47470
rect 34078 47458 34130 47470
rect 32610 47406 32622 47458
rect 32674 47406 32686 47458
rect 34290 47406 34302 47458
rect 34354 47406 34366 47458
rect 30158 47394 30210 47406
rect 34078 47394 34130 47406
rect 8094 47346 8146 47358
rect 20414 47346 20466 47358
rect 17602 47294 17614 47346
rect 17666 47294 17678 47346
rect 17938 47294 17950 47346
rect 18002 47294 18014 47346
rect 30482 47294 30494 47346
rect 30546 47294 30558 47346
rect 30818 47294 30830 47346
rect 30882 47294 30894 47346
rect 32946 47294 32958 47346
rect 33010 47294 33022 47346
rect 8094 47282 8146 47294
rect 20414 47282 20466 47294
rect 8318 47234 8370 47246
rect 8318 47170 8370 47182
rect 9214 47234 9266 47246
rect 20638 47234 20690 47246
rect 18162 47182 18174 47234
rect 18226 47182 18238 47234
rect 9214 47170 9266 47182
rect 20638 47170 20690 47182
rect 1344 47066 38640 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 38640 47066
rect 1344 46980 38640 47014
rect 10446 46898 10498 46910
rect 10446 46834 10498 46846
rect 11342 46898 11394 46910
rect 11342 46834 11394 46846
rect 15486 46898 15538 46910
rect 15486 46834 15538 46846
rect 21870 46898 21922 46910
rect 21870 46834 21922 46846
rect 32062 46898 32114 46910
rect 32062 46834 32114 46846
rect 8430 46786 8482 46798
rect 8430 46722 8482 46734
rect 8766 46786 8818 46798
rect 8766 46722 8818 46734
rect 9438 46786 9490 46798
rect 9438 46722 9490 46734
rect 9662 46786 9714 46798
rect 9662 46722 9714 46734
rect 10782 46786 10834 46798
rect 31726 46786 31778 46798
rect 30818 46734 30830 46786
rect 30882 46734 30894 46786
rect 31378 46734 31390 46786
rect 31442 46734 31454 46786
rect 10782 46722 10834 46734
rect 31726 46722 31778 46734
rect 31950 46786 32002 46798
rect 31950 46722 32002 46734
rect 32286 46786 32338 46798
rect 33058 46734 33070 46786
rect 33122 46734 33134 46786
rect 36082 46734 36094 46786
rect 36146 46734 36158 46786
rect 32286 46722 32338 46734
rect 8990 46674 9042 46686
rect 8990 46610 9042 46622
rect 9774 46674 9826 46686
rect 9774 46610 9826 46622
rect 10110 46674 10162 46686
rect 10110 46610 10162 46622
rect 10558 46674 10610 46686
rect 17950 46674 18002 46686
rect 21758 46674 21810 46686
rect 17490 46622 17502 46674
rect 17554 46622 17566 46674
rect 19170 46622 19182 46674
rect 19234 46622 19246 46674
rect 10558 46610 10610 46622
rect 17950 46610 18002 46622
rect 21758 46610 21810 46622
rect 21982 46674 22034 46686
rect 31614 46674 31666 46686
rect 22082 46622 22094 46674
rect 22146 46622 22158 46674
rect 28018 46622 28030 46674
rect 28082 46622 28094 46674
rect 21982 46610 22034 46622
rect 31614 46610 31666 46622
rect 32510 46674 32562 46686
rect 33282 46622 33294 46674
rect 33346 46622 33358 46674
rect 33730 46622 33742 46674
rect 33794 46622 33806 46674
rect 35298 46622 35310 46674
rect 35362 46622 35374 46674
rect 32510 46610 32562 46622
rect 8542 46562 8594 46574
rect 8542 46498 8594 46510
rect 15374 46562 15426 46574
rect 15374 46498 15426 46510
rect 15822 46562 15874 46574
rect 19282 46510 19294 46562
rect 19346 46510 19358 46562
rect 25218 46510 25230 46562
rect 25282 46510 25294 46562
rect 27346 46510 27358 46562
rect 27410 46510 27422 46562
rect 34626 46510 34638 46562
rect 34690 46510 34702 46562
rect 38210 46510 38222 46562
rect 38274 46510 38286 46562
rect 15822 46498 15874 46510
rect 15934 46450 15986 46462
rect 22430 46450 22482 46462
rect 19506 46398 19518 46450
rect 19570 46398 19582 46450
rect 15934 46386 15986 46398
rect 22430 46386 22482 46398
rect 1344 46282 38640 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 38640 46282
rect 1344 46196 38640 46230
rect 21646 46114 21698 46126
rect 21646 46050 21698 46062
rect 23998 46114 24050 46126
rect 23998 46050 24050 46062
rect 16942 46002 16994 46014
rect 30382 46002 30434 46014
rect 7298 45950 7310 46002
rect 7362 45950 7374 46002
rect 9426 45950 9438 46002
rect 9490 45950 9502 46002
rect 10770 45950 10782 46002
rect 10834 45950 10846 46002
rect 12898 45950 12910 46002
rect 12962 45950 12974 46002
rect 14914 45950 14926 46002
rect 14978 45950 14990 46002
rect 15810 45950 15822 46002
rect 15874 45950 15886 46002
rect 25666 45950 25678 46002
rect 25730 45950 25742 46002
rect 34738 45950 34750 46002
rect 34802 45950 34814 46002
rect 16942 45938 16994 45950
rect 30382 45938 30434 45950
rect 25230 45890 25282 45902
rect 30046 45890 30098 45902
rect 6514 45838 6526 45890
rect 6578 45838 6590 45890
rect 10098 45838 10110 45890
rect 10162 45838 10174 45890
rect 15362 45838 15374 45890
rect 15426 45838 15438 45890
rect 15922 45838 15934 45890
rect 15986 45838 15998 45890
rect 22082 45838 22094 45890
rect 22146 45838 22158 45890
rect 22418 45838 22430 45890
rect 22482 45838 22494 45890
rect 29586 45838 29598 45890
rect 29650 45838 29662 45890
rect 31378 45838 31390 45890
rect 31442 45838 31454 45890
rect 36418 45838 36430 45890
rect 36482 45838 36494 45890
rect 25230 45826 25282 45838
rect 30046 45826 30098 45838
rect 14590 45778 14642 45790
rect 21534 45778 21586 45790
rect 24110 45778 24162 45790
rect 14242 45726 14254 45778
rect 14306 45726 14318 45778
rect 16594 45726 16606 45778
rect 16658 45726 16670 45778
rect 23538 45726 23550 45778
rect 23602 45726 23614 45778
rect 14590 45714 14642 45726
rect 21534 45714 21586 45726
rect 24110 45714 24162 45726
rect 24558 45778 24610 45790
rect 24558 45714 24610 45726
rect 24894 45778 24946 45790
rect 33182 45778 33234 45790
rect 29250 45726 29262 45778
rect 29314 45726 29326 45778
rect 32274 45726 32286 45778
rect 32338 45726 32350 45778
rect 24894 45714 24946 45726
rect 33182 45714 33234 45726
rect 13918 45666 13970 45678
rect 13918 45602 13970 45614
rect 14814 45666 14866 45678
rect 14814 45602 14866 45614
rect 17054 45666 17106 45678
rect 33294 45666 33346 45678
rect 32386 45614 32398 45666
rect 32450 45614 32462 45666
rect 17054 45602 17106 45614
rect 33294 45602 33346 45614
rect 33406 45666 33458 45678
rect 33406 45602 33458 45614
rect 1344 45498 38640 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 38640 45498
rect 1344 45412 38640 45446
rect 8990 45330 9042 45342
rect 8990 45266 9042 45278
rect 9886 45330 9938 45342
rect 9886 45266 9938 45278
rect 10558 45330 10610 45342
rect 10558 45266 10610 45278
rect 10782 45330 10834 45342
rect 10782 45266 10834 45278
rect 14814 45330 14866 45342
rect 14814 45266 14866 45278
rect 17838 45330 17890 45342
rect 17838 45266 17890 45278
rect 18622 45330 18674 45342
rect 18622 45266 18674 45278
rect 25566 45330 25618 45342
rect 25566 45266 25618 45278
rect 26014 45330 26066 45342
rect 26014 45266 26066 45278
rect 26126 45330 26178 45342
rect 33058 45278 33070 45330
rect 33122 45278 33134 45330
rect 26126 45266 26178 45278
rect 2046 45218 2098 45230
rect 2046 45154 2098 45166
rect 6862 45218 6914 45230
rect 15038 45218 15090 45230
rect 10210 45166 10222 45218
rect 10274 45166 10286 45218
rect 6862 45154 6914 45166
rect 15038 45154 15090 45166
rect 18062 45218 18114 45230
rect 18062 45154 18114 45166
rect 18398 45218 18450 45230
rect 18398 45154 18450 45166
rect 18846 45218 18898 45230
rect 34638 45218 34690 45230
rect 23202 45166 23214 45218
rect 23266 45166 23278 45218
rect 30818 45166 30830 45218
rect 30882 45166 30894 45218
rect 32162 45166 32174 45218
rect 32226 45166 32238 45218
rect 18846 45154 18898 45166
rect 34638 45154 34690 45166
rect 1710 45106 1762 45118
rect 1710 45042 1762 45054
rect 6974 45106 7026 45118
rect 6974 45042 7026 45054
rect 10894 45106 10946 45118
rect 14478 45106 14530 45118
rect 16606 45106 16658 45118
rect 14018 45054 14030 45106
rect 14082 45054 14094 45106
rect 16034 45054 16046 45106
rect 16098 45054 16110 45106
rect 10894 45042 10946 45054
rect 14478 45042 14530 45054
rect 16606 45042 16658 45054
rect 17502 45106 17554 45118
rect 17502 45042 17554 45054
rect 19854 45106 19906 45118
rect 19854 45042 19906 45054
rect 19966 45106 20018 45118
rect 19966 45042 20018 45054
rect 22878 45106 22930 45118
rect 34078 45106 34130 45118
rect 29586 45054 29598 45106
rect 29650 45054 29662 45106
rect 30146 45054 30158 45106
rect 30210 45054 30222 45106
rect 32386 45054 32398 45106
rect 32450 45054 32462 45106
rect 33282 45054 33294 45106
rect 33346 45054 33358 45106
rect 22878 45042 22930 45054
rect 34078 45042 34130 45054
rect 34302 45106 34354 45118
rect 35298 45054 35310 45106
rect 35362 45054 35374 45106
rect 34302 45042 34354 45054
rect 2494 44994 2546 45006
rect 14242 44942 14254 44994
rect 14306 44942 14318 44994
rect 18722 44942 18734 44994
rect 18786 44942 18798 44994
rect 31938 44942 31950 44994
rect 32002 44942 32014 44994
rect 36082 44942 36094 44994
rect 36146 44942 36158 44994
rect 38210 44942 38222 44994
rect 38274 44942 38286 44994
rect 2494 44930 2546 44942
rect 6862 44882 6914 44894
rect 16718 44882 16770 44894
rect 15586 44830 15598 44882
rect 15650 44830 15662 44882
rect 6862 44818 6914 44830
rect 16718 44818 16770 44830
rect 18174 44882 18226 44894
rect 18174 44818 18226 44830
rect 20190 44882 20242 44894
rect 20190 44818 20242 44830
rect 20302 44882 20354 44894
rect 20302 44818 20354 44830
rect 26238 44882 26290 44894
rect 26238 44818 26290 44830
rect 34750 44882 34802 44894
rect 34750 44818 34802 44830
rect 34862 44882 34914 44894
rect 34862 44818 34914 44830
rect 1344 44714 38640 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 38640 44714
rect 1344 44628 38640 44662
rect 6750 44546 6802 44558
rect 20750 44546 20802 44558
rect 19954 44494 19966 44546
rect 20018 44494 20030 44546
rect 6750 44482 6802 44494
rect 20750 44482 20802 44494
rect 8318 44434 8370 44446
rect 10770 44382 10782 44434
rect 10834 44382 10846 44434
rect 12898 44382 12910 44434
rect 12962 44382 12974 44434
rect 21858 44382 21870 44434
rect 21922 44382 21934 44434
rect 24882 44382 24894 44434
rect 24946 44382 24958 44434
rect 35074 44382 35086 44434
rect 35138 44382 35150 44434
rect 8318 44370 8370 44382
rect 6638 44322 6690 44334
rect 6638 44258 6690 44270
rect 8542 44322 8594 44334
rect 8542 44258 8594 44270
rect 8766 44322 8818 44334
rect 15710 44322 15762 44334
rect 30606 44322 30658 44334
rect 10098 44270 10110 44322
rect 10162 44270 10174 44322
rect 13570 44270 13582 44322
rect 13634 44270 13646 44322
rect 17714 44270 17726 44322
rect 17778 44270 17790 44322
rect 21634 44270 21646 44322
rect 21698 44270 21710 44322
rect 23650 44270 23662 44322
rect 23714 44270 23726 44322
rect 26450 44270 26462 44322
rect 26514 44270 26526 44322
rect 30930 44270 30942 44322
rect 30994 44270 31006 44322
rect 8766 44258 8818 44270
rect 15710 44258 15762 44270
rect 30606 44258 30658 44270
rect 1710 44210 1762 44222
rect 1710 44146 1762 44158
rect 6750 44210 6802 44222
rect 6750 44146 6802 44158
rect 7534 44210 7586 44222
rect 7534 44146 7586 44158
rect 8206 44210 8258 44222
rect 16158 44210 16210 44222
rect 18958 44210 19010 44222
rect 13682 44158 13694 44210
rect 13746 44158 13758 44210
rect 17938 44158 17950 44210
rect 18002 44158 18014 44210
rect 18274 44158 18286 44210
rect 18338 44158 18350 44210
rect 8206 44146 8258 44158
rect 16158 44146 16210 44158
rect 18958 44146 19010 44158
rect 19182 44210 19234 44222
rect 19182 44146 19234 44158
rect 19406 44210 19458 44222
rect 19406 44146 19458 44158
rect 19630 44210 19682 44222
rect 19630 44146 19682 44158
rect 20414 44210 20466 44222
rect 20414 44146 20466 44158
rect 22318 44210 22370 44222
rect 23762 44158 23774 44210
rect 23826 44158 23838 44210
rect 24770 44158 24782 44210
rect 24834 44158 24846 44210
rect 22318 44146 22370 44158
rect 2046 44098 2098 44110
rect 2046 44034 2098 44046
rect 2494 44098 2546 44110
rect 2494 44034 2546 44046
rect 7646 44098 7698 44110
rect 7646 44034 7698 44046
rect 7870 44098 7922 44110
rect 20638 44098 20690 44110
rect 17266 44046 17278 44098
rect 17330 44046 17342 44098
rect 7870 44034 7922 44046
rect 20638 44034 20690 44046
rect 1344 43930 38640 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 38640 43930
rect 1344 43844 38640 43878
rect 9886 43762 9938 43774
rect 8194 43710 8206 43762
rect 8258 43710 8270 43762
rect 9886 43698 9938 43710
rect 12910 43762 12962 43774
rect 26450 43710 26462 43762
rect 26514 43710 26526 43762
rect 32162 43710 32174 43762
rect 32226 43710 32238 43762
rect 34402 43710 34414 43762
rect 34466 43710 34478 43762
rect 12910 43698 12962 43710
rect 10110 43650 10162 43662
rect 5954 43598 5966 43650
rect 6018 43598 6030 43650
rect 10110 43586 10162 43598
rect 10446 43650 10498 43662
rect 21422 43650 21474 43662
rect 27470 43650 27522 43662
rect 28590 43650 28642 43662
rect 12562 43598 12574 43650
rect 12626 43598 12638 43650
rect 24322 43598 24334 43650
rect 24386 43598 24398 43650
rect 27122 43598 27134 43650
rect 27186 43598 27198 43650
rect 27794 43598 27806 43650
rect 27858 43598 27870 43650
rect 10446 43586 10498 43598
rect 21422 43586 21474 43598
rect 27470 43586 27522 43598
rect 28590 43586 28642 43598
rect 30718 43650 30770 43662
rect 30818 43598 30830 43650
rect 30882 43647 30894 43650
rect 31154 43647 31166 43650
rect 30882 43601 31166 43647
rect 30882 43598 30894 43601
rect 31154 43598 31166 43601
rect 31218 43598 31230 43650
rect 31714 43598 31726 43650
rect 31778 43598 31790 43650
rect 32274 43598 32286 43650
rect 32338 43598 32350 43650
rect 33506 43598 33518 43650
rect 33570 43598 33582 43650
rect 30718 43586 30770 43598
rect 16382 43538 16434 43550
rect 5282 43486 5294 43538
rect 5346 43486 5358 43538
rect 13906 43486 13918 43538
rect 13970 43486 13982 43538
rect 16146 43486 16158 43538
rect 16210 43486 16222 43538
rect 16382 43474 16434 43486
rect 18286 43538 18338 43550
rect 18286 43474 18338 43486
rect 19854 43538 19906 43550
rect 19854 43474 19906 43486
rect 21198 43538 21250 43550
rect 21198 43474 21250 43486
rect 21534 43538 21586 43550
rect 23214 43538 23266 43550
rect 21858 43486 21870 43538
rect 21922 43486 21934 43538
rect 22194 43486 22206 43538
rect 22258 43486 22270 43538
rect 21534 43474 21586 43486
rect 23214 43474 23266 43486
rect 23550 43538 23602 43550
rect 23550 43474 23602 43486
rect 23662 43538 23714 43550
rect 23662 43474 23714 43486
rect 23886 43538 23938 43550
rect 23886 43474 23938 43486
rect 25566 43538 25618 43550
rect 25566 43474 25618 43486
rect 26126 43538 26178 43550
rect 26126 43474 26178 43486
rect 26798 43538 26850 43550
rect 28366 43538 28418 43550
rect 28018 43486 28030 43538
rect 28082 43486 28094 43538
rect 26798 43474 26850 43486
rect 28366 43474 28418 43486
rect 28702 43538 28754 43550
rect 28702 43474 28754 43486
rect 29598 43538 29650 43550
rect 29598 43474 29650 43486
rect 29822 43538 29874 43550
rect 29822 43474 29874 43486
rect 30046 43538 30098 43550
rect 30046 43474 30098 43486
rect 30270 43538 30322 43550
rect 30270 43474 30322 43486
rect 32398 43538 32450 43550
rect 33394 43486 33406 43538
rect 33458 43486 33470 43538
rect 33954 43486 33966 43538
rect 34018 43486 34030 43538
rect 35298 43486 35310 43538
rect 35362 43486 35374 43538
rect 32398 43474 32450 43486
rect 15934 43426 15986 43438
rect 19742 43426 19794 43438
rect 14018 43374 14030 43426
rect 14082 43374 14094 43426
rect 18610 43374 18622 43426
rect 18674 43374 18686 43426
rect 33730 43374 33742 43426
rect 33794 43374 33806 43426
rect 36082 43374 36094 43426
rect 36146 43374 36158 43426
rect 38210 43374 38222 43426
rect 38274 43374 38286 43426
rect 15934 43362 15986 43374
rect 19742 43362 19794 43374
rect 30158 43314 30210 43326
rect 18498 43262 18510 43314
rect 18562 43262 18574 43314
rect 30158 43250 30210 43262
rect 30606 43314 30658 43326
rect 30606 43250 30658 43262
rect 1344 43146 38640 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 38640 43146
rect 1344 43060 38640 43094
rect 14142 42978 14194 42990
rect 14142 42914 14194 42926
rect 20190 42978 20242 42990
rect 20190 42914 20242 42926
rect 20414 42978 20466 42990
rect 26226 42926 26238 42978
rect 26290 42926 26302 42978
rect 20414 42914 20466 42926
rect 31726 42866 31778 42878
rect 9874 42814 9886 42866
rect 9938 42814 9950 42866
rect 18386 42814 18398 42866
rect 18450 42814 18462 42866
rect 26002 42814 26014 42866
rect 26066 42814 26078 42866
rect 31726 42802 31778 42814
rect 32622 42866 32674 42878
rect 32622 42802 32674 42814
rect 10334 42754 10386 42766
rect 7074 42702 7086 42754
rect 7138 42702 7150 42754
rect 10334 42690 10386 42702
rect 10558 42754 10610 42766
rect 10558 42690 10610 42702
rect 10894 42754 10946 42766
rect 20638 42754 20690 42766
rect 28366 42754 28418 42766
rect 15138 42702 15150 42754
rect 15202 42702 15214 42754
rect 16034 42702 16046 42754
rect 16098 42702 16110 42754
rect 17714 42702 17726 42754
rect 17778 42702 17790 42754
rect 19954 42702 19966 42754
rect 20018 42702 20030 42754
rect 25666 42702 25678 42754
rect 25730 42702 25742 42754
rect 10894 42690 10946 42702
rect 20638 42690 20690 42702
rect 28366 42690 28418 42702
rect 28702 42754 28754 42766
rect 33070 42754 33122 42766
rect 29474 42702 29486 42754
rect 29538 42702 29550 42754
rect 29698 42702 29710 42754
rect 29762 42702 29774 42754
rect 30594 42702 30606 42754
rect 30658 42702 30670 42754
rect 28702 42690 28754 42702
rect 33070 42690 33122 42702
rect 33294 42754 33346 42766
rect 33294 42690 33346 42702
rect 33406 42754 33458 42766
rect 36418 42702 36430 42754
rect 36482 42702 36494 42754
rect 33406 42690 33458 42702
rect 15374 42642 15426 42654
rect 20750 42642 20802 42654
rect 7746 42590 7758 42642
rect 7810 42590 7822 42642
rect 14690 42590 14702 42642
rect 14754 42590 14766 42642
rect 16594 42590 16606 42642
rect 16658 42590 16670 42642
rect 17602 42590 17614 42642
rect 17666 42590 17678 42642
rect 15374 42578 15426 42590
rect 20750 42578 20802 42590
rect 21310 42642 21362 42654
rect 31166 42642 31218 42654
rect 30034 42590 30046 42642
rect 30098 42590 30110 42642
rect 21310 42578 21362 42590
rect 31166 42578 31218 42590
rect 31278 42642 31330 42654
rect 31278 42578 31330 42590
rect 31614 42642 31666 42654
rect 31614 42578 31666 42590
rect 32062 42642 32114 42654
rect 32062 42578 32114 42590
rect 32846 42642 32898 42654
rect 32846 42578 32898 42590
rect 10558 42530 10610 42542
rect 10558 42466 10610 42478
rect 11230 42530 11282 42542
rect 11230 42466 11282 42478
rect 21422 42530 21474 42542
rect 21422 42466 21474 42478
rect 21646 42530 21698 42542
rect 21646 42466 21698 42478
rect 26798 42530 26850 42542
rect 26798 42466 26850 42478
rect 28478 42530 28530 42542
rect 28478 42466 28530 42478
rect 30942 42530 30994 42542
rect 30942 42466 30994 42478
rect 32286 42530 32338 42542
rect 32286 42466 32338 42478
rect 32510 42530 32562 42542
rect 32510 42466 32562 42478
rect 33182 42530 33234 42542
rect 33182 42466 33234 42478
rect 35422 42530 35474 42542
rect 35422 42466 35474 42478
rect 1344 42362 38640 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 38640 42362
rect 1344 42276 38640 42310
rect 7982 42194 8034 42206
rect 7982 42130 8034 42142
rect 8206 42194 8258 42206
rect 8206 42130 8258 42142
rect 16046 42194 16098 42206
rect 28142 42194 28194 42206
rect 20402 42142 20414 42194
rect 20466 42142 20478 42194
rect 16046 42130 16098 42142
rect 28142 42130 28194 42142
rect 33294 42194 33346 42206
rect 33294 42130 33346 42142
rect 34414 42194 34466 42206
rect 34414 42130 34466 42142
rect 8318 42082 8370 42094
rect 8318 42018 8370 42030
rect 22766 42082 22818 42094
rect 22766 42018 22818 42030
rect 22878 42082 22930 42094
rect 31278 42082 31330 42094
rect 30258 42030 30270 42082
rect 30322 42030 30334 42082
rect 30594 42030 30606 42082
rect 30658 42030 30670 42082
rect 22878 42018 22930 42030
rect 31278 42018 31330 42030
rect 14814 41970 14866 41982
rect 18286 41970 18338 41982
rect 16594 41918 16606 41970
rect 16658 41918 16670 41970
rect 14814 41906 14866 41918
rect 18286 41906 18338 41918
rect 18622 41970 18674 41982
rect 18622 41906 18674 41918
rect 18734 41970 18786 41982
rect 18734 41906 18786 41918
rect 18958 41970 19010 41982
rect 19854 41970 19906 41982
rect 19618 41918 19630 41970
rect 19682 41918 19694 41970
rect 18958 41906 19010 41918
rect 19854 41906 19906 41918
rect 19966 41970 20018 41982
rect 19966 41906 20018 41918
rect 22542 41970 22594 41982
rect 22542 41906 22594 41918
rect 25230 41970 25282 41982
rect 28254 41970 28306 41982
rect 27794 41918 27806 41970
rect 27858 41918 27870 41970
rect 25230 41906 25282 41918
rect 28254 41906 28306 41918
rect 28366 41970 28418 41982
rect 31054 41970 31106 41982
rect 29250 41918 29262 41970
rect 29314 41918 29326 41970
rect 29474 41918 29486 41970
rect 29538 41918 29550 41970
rect 28366 41906 28418 41918
rect 31054 41906 31106 41918
rect 31502 41970 31554 41982
rect 31502 41906 31554 41918
rect 31726 41970 31778 41982
rect 31726 41906 31778 41918
rect 31950 41970 32002 41982
rect 32958 41970 33010 41982
rect 32274 41918 32286 41970
rect 32338 41918 32350 41970
rect 31950 41906 32002 41918
rect 32958 41906 33010 41918
rect 33294 41970 33346 41982
rect 33294 41906 33346 41918
rect 33630 41970 33682 41982
rect 34526 41970 34578 41982
rect 34178 41918 34190 41970
rect 34242 41918 34254 41970
rect 33630 41906 33682 41918
rect 34526 41906 34578 41918
rect 34638 41970 34690 41982
rect 34638 41906 34690 41918
rect 34750 41970 34802 41982
rect 35410 41918 35422 41970
rect 35474 41918 35486 41970
rect 34750 41906 34802 41918
rect 17502 41858 17554 41870
rect 17502 41794 17554 41806
rect 25678 41858 25730 41870
rect 25678 41794 25730 41806
rect 29710 41858 29762 41870
rect 36082 41806 36094 41858
rect 36146 41806 36158 41858
rect 38210 41806 38222 41858
rect 38274 41806 38286 41858
rect 29710 41794 29762 41806
rect 14926 41746 14978 41758
rect 14926 41682 14978 41694
rect 25454 41746 25506 41758
rect 25454 41682 25506 41694
rect 25902 41746 25954 41758
rect 25902 41682 25954 41694
rect 26350 41746 26402 41758
rect 26350 41682 26402 41694
rect 1344 41578 38640 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 38640 41578
rect 1344 41492 38640 41526
rect 22542 41410 22594 41422
rect 29362 41358 29374 41410
rect 29426 41358 29438 41410
rect 34962 41358 34974 41410
rect 35026 41358 35038 41410
rect 22542 41346 22594 41358
rect 20078 41298 20130 41310
rect 20078 41234 20130 41246
rect 20638 41298 20690 41310
rect 30606 41298 30658 41310
rect 29586 41246 29598 41298
rect 29650 41246 29662 41298
rect 20638 41234 20690 41246
rect 30606 41234 30658 41246
rect 31390 41298 31442 41310
rect 31390 41234 31442 41246
rect 10894 41186 10946 41198
rect 1810 41134 1822 41186
rect 1874 41134 1886 41186
rect 10894 41122 10946 41134
rect 11230 41186 11282 41198
rect 11230 41122 11282 41134
rect 11566 41186 11618 41198
rect 11566 41122 11618 41134
rect 11902 41186 11954 41198
rect 19854 41186 19906 41198
rect 19170 41134 19182 41186
rect 19234 41134 19246 41186
rect 11902 41122 11954 41134
rect 19854 41122 19906 41134
rect 21646 41186 21698 41198
rect 22990 41186 23042 41198
rect 26238 41186 26290 41198
rect 22082 41134 22094 41186
rect 22146 41134 22158 41186
rect 24098 41134 24110 41186
rect 24162 41134 24174 41186
rect 21646 41122 21698 41134
rect 22990 41122 23042 41134
rect 26238 41122 26290 41134
rect 28702 41186 28754 41198
rect 28702 41122 28754 41134
rect 31054 41186 31106 41198
rect 31054 41122 31106 41134
rect 31278 41186 31330 41198
rect 32622 41186 32674 41198
rect 31714 41134 31726 41186
rect 31778 41134 31790 41186
rect 31278 41122 31330 41134
rect 32622 41122 32674 41134
rect 33182 41186 33234 41198
rect 36306 41134 36318 41186
rect 36370 41134 36382 41186
rect 33182 41122 33234 41134
rect 2494 41074 2546 41086
rect 19630 41074 19682 41086
rect 14130 41022 14142 41074
rect 14194 41022 14206 41074
rect 2494 41010 2546 41022
rect 19630 41010 19682 41022
rect 20190 41074 20242 41086
rect 20190 41010 20242 41022
rect 21758 41074 21810 41086
rect 21758 41010 21810 41022
rect 21870 41074 21922 41086
rect 21870 41010 21922 41022
rect 24782 41074 24834 41086
rect 24782 41010 24834 41022
rect 26798 41074 26850 41086
rect 26798 41010 26850 41022
rect 28366 41074 28418 41086
rect 32734 41074 32786 41086
rect 29250 41022 29262 41074
rect 29314 41022 29326 41074
rect 31826 41022 31838 41074
rect 31890 41022 31902 41074
rect 28366 41010 28418 41022
rect 32734 41010 32786 41022
rect 33518 41074 33570 41086
rect 33518 41010 33570 41022
rect 2046 40962 2098 40974
rect 2046 40898 2098 40910
rect 11342 40962 11394 40974
rect 11342 40898 11394 40910
rect 23102 40962 23154 40974
rect 23102 40898 23154 40910
rect 23214 40962 23266 40974
rect 23214 40898 23266 40910
rect 23438 40962 23490 40974
rect 28478 40962 28530 40974
rect 27794 40910 27806 40962
rect 27858 40910 27870 40962
rect 23438 40898 23490 40910
rect 28478 40898 28530 40910
rect 31502 40962 31554 40974
rect 31502 40898 31554 40910
rect 32958 40962 33010 40974
rect 32958 40898 33010 40910
rect 1344 40794 38640 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 38640 40794
rect 1344 40708 38640 40742
rect 9774 40626 9826 40638
rect 9774 40562 9826 40574
rect 10334 40626 10386 40638
rect 10334 40562 10386 40574
rect 14254 40626 14306 40638
rect 14254 40562 14306 40574
rect 18846 40626 18898 40638
rect 18846 40562 18898 40574
rect 19854 40626 19906 40638
rect 19854 40562 19906 40574
rect 20190 40626 20242 40638
rect 20190 40562 20242 40574
rect 22430 40626 22482 40638
rect 22430 40562 22482 40574
rect 30158 40626 30210 40638
rect 30158 40562 30210 40574
rect 30382 40626 30434 40638
rect 30382 40562 30434 40574
rect 30718 40626 30770 40638
rect 30718 40562 30770 40574
rect 31950 40626 32002 40638
rect 31950 40562 32002 40574
rect 32398 40626 32450 40638
rect 32398 40562 32450 40574
rect 2046 40514 2098 40526
rect 2046 40450 2098 40462
rect 9662 40514 9714 40526
rect 9662 40450 9714 40462
rect 20078 40514 20130 40526
rect 20078 40450 20130 40462
rect 20414 40514 20466 40526
rect 20414 40450 20466 40462
rect 23326 40514 23378 40526
rect 23326 40450 23378 40462
rect 32510 40514 32562 40526
rect 33842 40462 33854 40514
rect 33906 40462 33918 40514
rect 32510 40450 32562 40462
rect 1710 40402 1762 40414
rect 1710 40338 1762 40350
rect 2494 40402 2546 40414
rect 19518 40402 19570 40414
rect 13234 40350 13246 40402
rect 13298 40350 13310 40402
rect 13458 40350 13470 40402
rect 13522 40350 13534 40402
rect 2494 40338 2546 40350
rect 19518 40338 19570 40350
rect 21310 40402 21362 40414
rect 30046 40402 30098 40414
rect 24322 40350 24334 40402
rect 24386 40350 24398 40402
rect 21310 40338 21362 40350
rect 30046 40338 30098 40350
rect 30606 40402 30658 40414
rect 30606 40338 30658 40350
rect 30942 40402 30994 40414
rect 32062 40402 32114 40414
rect 31378 40350 31390 40402
rect 31442 40350 31454 40402
rect 33170 40350 33182 40402
rect 33234 40350 33246 40402
rect 30942 40338 30994 40350
rect 32062 40338 32114 40350
rect 20974 40290 21026 40302
rect 13682 40238 13694 40290
rect 13746 40238 13758 40290
rect 20974 40226 21026 40238
rect 21534 40290 21586 40302
rect 21534 40226 21586 40238
rect 21758 40290 21810 40302
rect 21758 40226 21810 40238
rect 23662 40290 23714 40302
rect 23986 40238 23998 40290
rect 24050 40238 24062 40290
rect 35970 40238 35982 40290
rect 36034 40238 36046 40290
rect 23662 40226 23714 40238
rect 9774 40178 9826 40190
rect 9774 40114 9826 40126
rect 20638 40178 20690 40190
rect 20638 40114 20690 40126
rect 21982 40178 22034 40190
rect 21982 40114 22034 40126
rect 1344 40010 38640 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 38640 40010
rect 1344 39924 38640 39958
rect 18834 39790 18846 39842
rect 18898 39839 18910 39842
rect 18898 39793 19119 39839
rect 18898 39790 18910 39793
rect 19073 39730 19119 39793
rect 19630 39730 19682 39742
rect 12898 39678 12910 39730
rect 12962 39678 12974 39730
rect 19058 39678 19070 39730
rect 19122 39678 19134 39730
rect 19630 39666 19682 39678
rect 20190 39730 20242 39742
rect 29598 39730 29650 39742
rect 25554 39678 25566 39730
rect 25618 39678 25630 39730
rect 33170 39678 33182 39730
rect 33234 39678 33246 39730
rect 20190 39666 20242 39678
rect 29598 39666 29650 39678
rect 8542 39618 8594 39630
rect 8542 39554 8594 39566
rect 8766 39618 8818 39630
rect 8766 39554 8818 39566
rect 9214 39618 9266 39630
rect 9214 39554 9266 39566
rect 9774 39618 9826 39630
rect 18510 39618 18562 39630
rect 10098 39566 10110 39618
rect 10162 39566 10174 39618
rect 16370 39566 16382 39618
rect 16434 39566 16446 39618
rect 9774 39554 9826 39566
rect 18510 39554 18562 39566
rect 19518 39618 19570 39630
rect 19518 39554 19570 39566
rect 19966 39618 20018 39630
rect 19966 39554 20018 39566
rect 20302 39618 20354 39630
rect 22754 39566 22766 39618
rect 22818 39566 22830 39618
rect 22978 39566 22990 39618
rect 23042 39566 23054 39618
rect 24770 39566 24782 39618
rect 24834 39566 24846 39618
rect 30818 39566 30830 39618
rect 30882 39566 30894 39618
rect 20302 39554 20354 39566
rect 1710 39506 1762 39518
rect 1710 39442 1762 39454
rect 8206 39506 8258 39518
rect 8206 39442 8258 39454
rect 9326 39506 9378 39518
rect 17390 39506 17442 39518
rect 10770 39454 10782 39506
rect 10834 39454 10846 39506
rect 14914 39454 14926 39506
rect 14978 39454 14990 39506
rect 9326 39442 9378 39454
rect 17390 39442 17442 39454
rect 19294 39506 19346 39518
rect 19294 39442 19346 39454
rect 20638 39506 20690 39518
rect 25778 39454 25790 39506
rect 25842 39454 25854 39506
rect 20638 39442 20690 39454
rect 2046 39394 2098 39406
rect 2046 39330 2098 39342
rect 2494 39394 2546 39406
rect 2494 39330 2546 39342
rect 8430 39394 8482 39406
rect 8430 39330 8482 39342
rect 9438 39394 9490 39406
rect 19742 39394 19794 39406
rect 15026 39342 15038 39394
rect 15090 39342 15102 39394
rect 9438 39330 9490 39342
rect 19742 39330 19794 39342
rect 1344 39226 38640 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 38640 39226
rect 1344 39140 38640 39174
rect 8206 39058 8258 39070
rect 8206 38994 8258 39006
rect 9662 39058 9714 39070
rect 9662 38994 9714 39006
rect 10334 39058 10386 39070
rect 10334 38994 10386 39006
rect 10670 39058 10722 39070
rect 10670 38994 10722 39006
rect 11118 39058 11170 39070
rect 26238 39058 26290 39070
rect 18386 39006 18398 39058
rect 18450 39006 18462 39058
rect 11118 38994 11170 39006
rect 26238 38994 26290 39006
rect 26910 39058 26962 39070
rect 26910 38994 26962 39006
rect 7534 38946 7586 38958
rect 7534 38882 7586 38894
rect 7646 38946 7698 38958
rect 7646 38882 7698 38894
rect 8094 38946 8146 38958
rect 8094 38882 8146 38894
rect 8766 38946 8818 38958
rect 8766 38882 8818 38894
rect 9550 38946 9602 38958
rect 9550 38882 9602 38894
rect 9886 38946 9938 38958
rect 9886 38882 9938 38894
rect 11342 38946 11394 38958
rect 11342 38882 11394 38894
rect 11454 38946 11506 38958
rect 11454 38882 11506 38894
rect 12574 38946 12626 38958
rect 12574 38882 12626 38894
rect 12686 38946 12738 38958
rect 12686 38882 12738 38894
rect 13022 38946 13074 38958
rect 15710 38946 15762 38958
rect 19070 38946 19122 38958
rect 14018 38894 14030 38946
rect 14082 38894 14094 38946
rect 17826 38894 17838 38946
rect 17890 38894 17902 38946
rect 13022 38882 13074 38894
rect 15710 38882 15762 38894
rect 19070 38882 19122 38894
rect 19182 38946 19234 38958
rect 25342 38946 25394 38958
rect 23314 38894 23326 38946
rect 23378 38894 23390 38946
rect 19182 38882 19234 38894
rect 25342 38882 25394 38894
rect 26126 38946 26178 38958
rect 34178 38894 34190 38946
rect 34242 38894 34254 38946
rect 26126 38882 26178 38894
rect 7870 38834 7922 38846
rect 7870 38770 7922 38782
rect 8430 38834 8482 38846
rect 8430 38770 8482 38782
rect 8654 38834 8706 38846
rect 8654 38770 8706 38782
rect 8990 38834 9042 38846
rect 25230 38834 25282 38846
rect 15138 38782 15150 38834
rect 15202 38782 15214 38834
rect 17378 38782 17390 38834
rect 17442 38782 17454 38834
rect 18274 38782 18286 38834
rect 18338 38782 18350 38834
rect 18834 38782 18846 38834
rect 18898 38782 18910 38834
rect 19618 38782 19630 38834
rect 19682 38782 19694 38834
rect 20402 38782 20414 38834
rect 20466 38782 20478 38834
rect 20626 38782 20638 38834
rect 20690 38782 20702 38834
rect 21634 38782 21646 38834
rect 21698 38782 21710 38834
rect 23650 38782 23662 38834
rect 23714 38782 23726 38834
rect 24322 38782 24334 38834
rect 24386 38782 24398 38834
rect 8990 38770 9042 38782
rect 25230 38770 25282 38782
rect 26462 38834 26514 38846
rect 33394 38782 33406 38834
rect 33458 38782 33470 38834
rect 26462 38770 26514 38782
rect 13694 38722 13746 38734
rect 22766 38722 22818 38734
rect 21522 38670 21534 38722
rect 21586 38670 21598 38722
rect 22082 38670 22094 38722
rect 22146 38670 22158 38722
rect 13694 38658 13746 38670
rect 22766 38658 22818 38670
rect 23550 38722 23602 38734
rect 36306 38670 36318 38722
rect 36370 38670 36382 38722
rect 23550 38658 23602 38670
rect 13134 38610 13186 38622
rect 13134 38546 13186 38558
rect 22542 38610 22594 38622
rect 22542 38546 22594 38558
rect 22878 38610 22930 38622
rect 22878 38546 22930 38558
rect 1344 38442 38640 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 38640 38442
rect 1344 38356 38640 38390
rect 23774 38274 23826 38286
rect 23774 38210 23826 38222
rect 24446 38274 24498 38286
rect 26014 38274 26066 38286
rect 24770 38222 24782 38274
rect 24834 38222 24846 38274
rect 25666 38222 25678 38274
rect 25730 38222 25742 38274
rect 24446 38210 24498 38222
rect 26014 38210 26066 38222
rect 26910 38274 26962 38286
rect 26910 38210 26962 38222
rect 27582 38274 27634 38286
rect 34962 38222 34974 38274
rect 35026 38222 35038 38274
rect 27582 38210 27634 38222
rect 6974 38162 7026 38174
rect 22094 38162 22146 38174
rect 9090 38110 9102 38162
rect 9154 38110 9166 38162
rect 14914 38110 14926 38162
rect 14978 38110 14990 38162
rect 6974 38098 7026 38110
rect 22094 38098 22146 38110
rect 24222 38162 24274 38174
rect 24222 38098 24274 38110
rect 25454 38162 25506 38174
rect 28030 38162 28082 38174
rect 26562 38110 26574 38162
rect 26626 38110 26638 38162
rect 29474 38110 29486 38162
rect 29538 38110 29550 38162
rect 31602 38110 31614 38162
rect 31666 38110 31678 38162
rect 25454 38098 25506 38110
rect 28030 38098 28082 38110
rect 21646 38050 21698 38062
rect 26238 38050 26290 38062
rect 9874 37998 9886 38050
rect 9938 37998 9950 38050
rect 14018 37998 14030 38050
rect 14082 37998 14094 38050
rect 15026 37998 15038 38050
rect 15090 37998 15102 38050
rect 20066 37998 20078 38050
rect 20130 37998 20142 38050
rect 22642 37998 22654 38050
rect 22706 37998 22718 38050
rect 22866 37998 22878 38050
rect 22930 37998 22942 38050
rect 23538 37998 23550 38050
rect 23602 37998 23614 38050
rect 27234 37998 27246 38050
rect 27298 37998 27310 38050
rect 32386 37998 32398 38050
rect 32450 37998 32462 38050
rect 36306 37998 36318 38050
rect 36370 37998 36382 38050
rect 21646 37986 21698 37998
rect 26238 37986 26290 37998
rect 21310 37938 21362 37950
rect 14690 37886 14702 37938
rect 14754 37886 14766 37938
rect 16930 37886 16942 37938
rect 16994 37886 17006 37938
rect 21310 37874 21362 37886
rect 26686 37938 26738 37950
rect 26686 37874 26738 37886
rect 10334 37826 10386 37838
rect 10334 37762 10386 37774
rect 21422 37826 21474 37838
rect 21422 37762 21474 37774
rect 27470 37826 27522 37838
rect 27470 37762 27522 37774
rect 1344 37658 38640 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 38640 37658
rect 1344 37572 38640 37606
rect 16270 37490 16322 37502
rect 16270 37426 16322 37438
rect 28478 37490 28530 37502
rect 28478 37426 28530 37438
rect 19742 37378 19794 37390
rect 19742 37314 19794 37326
rect 19854 37378 19906 37390
rect 19854 37314 19906 37326
rect 25342 37378 25394 37390
rect 25342 37314 25394 37326
rect 26462 37378 26514 37390
rect 26462 37314 26514 37326
rect 28030 37378 28082 37390
rect 28030 37314 28082 37326
rect 27134 37266 27186 37278
rect 25442 37214 25454 37266
rect 25506 37214 25518 37266
rect 25890 37214 25902 37266
rect 25954 37214 25966 37266
rect 26674 37214 26686 37266
rect 26738 37214 26750 37266
rect 27346 37214 27358 37266
rect 27410 37214 27422 37266
rect 27134 37202 27186 37214
rect 16158 37154 16210 37166
rect 16158 37090 16210 37102
rect 28926 37154 28978 37166
rect 28926 37090 28978 37102
rect 19854 37042 19906 37054
rect 19854 36978 19906 36990
rect 1344 36874 38640 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 38640 36874
rect 1344 36788 38640 36822
rect 17950 36594 18002 36606
rect 8754 36542 8766 36594
rect 8818 36542 8830 36594
rect 10882 36542 10894 36594
rect 10946 36542 10958 36594
rect 24658 36542 24670 36594
rect 24722 36542 24734 36594
rect 17950 36530 18002 36542
rect 18622 36482 18674 36494
rect 8082 36430 8094 36482
rect 8146 36430 8158 36482
rect 16370 36430 16382 36482
rect 16434 36430 16446 36482
rect 27570 36430 27582 36482
rect 27634 36430 27646 36482
rect 18622 36418 18674 36430
rect 18286 36370 18338 36382
rect 38222 36370 38274 36382
rect 16034 36318 16046 36370
rect 16098 36318 16110 36370
rect 17714 36318 17726 36370
rect 17778 36318 17790 36370
rect 26786 36318 26798 36370
rect 26850 36318 26862 36370
rect 18286 36306 18338 36318
rect 38222 36306 38274 36318
rect 11342 36258 11394 36270
rect 11342 36194 11394 36206
rect 14590 36258 14642 36270
rect 14590 36194 14642 36206
rect 28030 36258 28082 36270
rect 28030 36194 28082 36206
rect 1344 36090 38640 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 38640 36090
rect 1344 36004 38640 36038
rect 22542 35922 22594 35934
rect 22542 35858 22594 35870
rect 25790 35922 25842 35934
rect 25790 35858 25842 35870
rect 14926 35810 14978 35822
rect 14926 35746 14978 35758
rect 15262 35810 15314 35822
rect 15262 35746 15314 35758
rect 22654 35810 22706 35822
rect 27682 35758 27694 35810
rect 27746 35758 27758 35810
rect 22654 35746 22706 35758
rect 25678 35698 25730 35710
rect 11554 35646 11566 35698
rect 11618 35646 11630 35698
rect 17714 35646 17726 35698
rect 17778 35646 17790 35698
rect 21858 35646 21870 35698
rect 21922 35646 21934 35698
rect 26898 35646 26910 35698
rect 26962 35646 26974 35698
rect 25678 35634 25730 35646
rect 15822 35586 15874 35598
rect 22094 35586 22146 35598
rect 12226 35534 12238 35586
rect 12290 35534 12302 35586
rect 14354 35534 14366 35586
rect 14418 35534 14430 35586
rect 17602 35534 17614 35586
rect 17666 35534 17678 35586
rect 29810 35534 29822 35586
rect 29874 35534 29886 35586
rect 15822 35522 15874 35534
rect 22094 35522 22146 35534
rect 17390 35474 17442 35486
rect 17390 35410 17442 35422
rect 22206 35474 22258 35486
rect 22206 35410 22258 35422
rect 25454 35474 25506 35486
rect 25454 35410 25506 35422
rect 25790 35474 25842 35486
rect 25790 35410 25842 35422
rect 1344 35306 38640 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 38640 35306
rect 1344 35220 38640 35254
rect 13470 35138 13522 35150
rect 13470 35074 13522 35086
rect 15150 35026 15202 35038
rect 22654 35026 22706 35038
rect 19170 34974 19182 35026
rect 19234 34974 19246 35026
rect 15150 34962 15202 34974
rect 22654 34962 22706 34974
rect 23102 35026 23154 35038
rect 23102 34962 23154 34974
rect 14366 34914 14418 34926
rect 14366 34850 14418 34862
rect 14814 34914 14866 34926
rect 14814 34850 14866 34862
rect 15262 34914 15314 34926
rect 15262 34850 15314 34862
rect 15598 34914 15650 34926
rect 21758 34914 21810 34926
rect 16370 34862 16382 34914
rect 16434 34862 16446 34914
rect 22194 34862 22206 34914
rect 22258 34862 22270 34914
rect 15598 34850 15650 34862
rect 21758 34850 21810 34862
rect 13582 34802 13634 34814
rect 13582 34738 13634 34750
rect 14254 34802 14306 34814
rect 14254 34738 14306 34750
rect 15038 34802 15090 34814
rect 17042 34750 17054 34802
rect 17106 34750 17118 34802
rect 15038 34738 15090 34750
rect 14142 34690 14194 34702
rect 14142 34626 14194 34638
rect 19630 34690 19682 34702
rect 19630 34626 19682 34638
rect 1344 34522 38640 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 38640 34522
rect 1344 34436 38640 34470
rect 15150 34354 15202 34366
rect 15150 34290 15202 34302
rect 17502 34354 17554 34366
rect 22766 34354 22818 34366
rect 21074 34302 21086 34354
rect 21138 34302 21150 34354
rect 24658 34302 24670 34354
rect 24722 34302 24734 34354
rect 17502 34290 17554 34302
rect 22766 34290 22818 34302
rect 16270 34242 16322 34254
rect 16270 34178 16322 34190
rect 16382 34242 16434 34254
rect 22318 34242 22370 34254
rect 20290 34190 20302 34242
rect 20354 34190 20366 34242
rect 16382 34178 16434 34190
rect 22318 34178 22370 34190
rect 17614 34130 17666 34142
rect 20526 34130 20578 34142
rect 11778 34078 11790 34130
rect 11842 34078 11854 34130
rect 16034 34078 16046 34130
rect 16098 34078 16110 34130
rect 17378 34078 17390 34130
rect 17442 34078 17454 34130
rect 20066 34078 20078 34130
rect 20130 34078 20142 34130
rect 17614 34066 17666 34078
rect 20526 34066 20578 34078
rect 20638 34130 20690 34142
rect 20638 34066 20690 34078
rect 21646 34130 21698 34142
rect 25342 34130 25394 34142
rect 21970 34078 21982 34130
rect 22034 34078 22046 34130
rect 24434 34078 24446 34130
rect 24498 34078 24510 34130
rect 25554 34078 25566 34130
rect 25618 34078 25630 34130
rect 21646 34066 21698 34078
rect 25342 34066 25394 34078
rect 16606 34018 16658 34030
rect 12562 33966 12574 34018
rect 12626 33966 12638 34018
rect 14690 33966 14702 34018
rect 14754 33966 14766 34018
rect 16606 33954 16658 33966
rect 21422 34018 21474 34030
rect 21422 33954 21474 33966
rect 26238 34018 26290 34030
rect 26238 33954 26290 33966
rect 15598 33906 15650 33918
rect 15598 33842 15650 33854
rect 17838 33906 17890 33918
rect 17838 33842 17890 33854
rect 19742 33906 19794 33918
rect 19742 33842 19794 33854
rect 21982 33906 22034 33918
rect 21982 33842 22034 33854
rect 1344 33738 38640 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 38640 33738
rect 1344 33652 38640 33686
rect 13918 33570 13970 33582
rect 13918 33506 13970 33518
rect 14366 33570 14418 33582
rect 14366 33506 14418 33518
rect 17166 33570 17218 33582
rect 17166 33506 17218 33518
rect 18734 33570 18786 33582
rect 18734 33506 18786 33518
rect 19070 33570 19122 33582
rect 19070 33506 19122 33518
rect 21422 33570 21474 33582
rect 21422 33506 21474 33518
rect 21646 33570 21698 33582
rect 21646 33506 21698 33518
rect 26014 33570 26066 33582
rect 26014 33506 26066 33518
rect 13694 33458 13746 33470
rect 13694 33394 13746 33406
rect 14030 33458 14082 33470
rect 14030 33394 14082 33406
rect 17390 33458 17442 33470
rect 17390 33394 17442 33406
rect 22318 33458 22370 33470
rect 22318 33394 22370 33406
rect 23998 33458 24050 33470
rect 23998 33394 24050 33406
rect 24894 33458 24946 33470
rect 24894 33394 24946 33406
rect 26798 33458 26850 33470
rect 26798 33394 26850 33406
rect 14254 33346 14306 33358
rect 14254 33282 14306 33294
rect 14814 33346 14866 33358
rect 14814 33282 14866 33294
rect 15150 33346 15202 33358
rect 15150 33282 15202 33294
rect 15374 33346 15426 33358
rect 18958 33346 19010 33358
rect 16818 33294 16830 33346
rect 16882 33294 16894 33346
rect 15374 33282 15426 33294
rect 18958 33282 19010 33294
rect 19966 33346 20018 33358
rect 19966 33282 20018 33294
rect 20190 33346 20242 33358
rect 20190 33282 20242 33294
rect 20302 33346 20354 33358
rect 20302 33282 20354 33294
rect 20526 33346 20578 33358
rect 20526 33282 20578 33294
rect 21758 33346 21810 33358
rect 26338 33294 26350 33346
rect 26402 33294 26414 33346
rect 21758 33282 21810 33294
rect 14926 33234 14978 33246
rect 14926 33170 14978 33182
rect 18622 33234 18674 33246
rect 18622 33170 18674 33182
rect 21310 33234 21362 33246
rect 21310 33170 21362 33182
rect 1710 33122 1762 33134
rect 1710 33058 1762 33070
rect 26126 33122 26178 33134
rect 26126 33058 26178 33070
rect 1344 32954 38640 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 38640 32954
rect 1344 32868 38640 32902
rect 24222 32786 24274 32798
rect 24222 32722 24274 32734
rect 23550 32674 23602 32686
rect 21074 32622 21086 32674
rect 21138 32622 21150 32674
rect 23550 32610 23602 32622
rect 23774 32674 23826 32686
rect 27458 32622 27470 32674
rect 27522 32622 27534 32674
rect 23774 32610 23826 32622
rect 14702 32562 14754 32574
rect 14018 32510 14030 32562
rect 14082 32510 14094 32562
rect 14702 32498 14754 32510
rect 14926 32562 14978 32574
rect 23214 32562 23266 32574
rect 21858 32510 21870 32562
rect 21922 32510 21934 32562
rect 14926 32498 14978 32510
rect 23214 32498 23266 32510
rect 24334 32562 24386 32574
rect 28130 32510 28142 32562
rect 28194 32510 28206 32562
rect 24334 32498 24386 32510
rect 14366 32450 14418 32462
rect 14366 32386 14418 32398
rect 18622 32450 18674 32462
rect 23326 32450 23378 32462
rect 18946 32398 18958 32450
rect 19010 32398 19022 32450
rect 25330 32398 25342 32450
rect 25394 32398 25406 32450
rect 18622 32386 18674 32398
rect 23326 32386 23378 32398
rect 14030 32338 14082 32350
rect 24222 32338 24274 32350
rect 15250 32286 15262 32338
rect 15314 32286 15326 32338
rect 14030 32274 14082 32286
rect 24222 32274 24274 32286
rect 1344 32170 38640 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 38640 32170
rect 1344 32084 38640 32118
rect 14702 32002 14754 32014
rect 14702 31938 14754 31950
rect 23426 31838 23438 31890
rect 23490 31838 23502 31890
rect 14478 31778 14530 31790
rect 15486 31778 15538 31790
rect 14914 31726 14926 31778
rect 14978 31726 14990 31778
rect 14478 31714 14530 31726
rect 15486 31714 15538 31726
rect 22542 31778 22594 31790
rect 22542 31714 22594 31726
rect 22766 31778 22818 31790
rect 22766 31714 22818 31726
rect 23214 31778 23266 31790
rect 26338 31726 26350 31778
rect 26402 31726 26414 31778
rect 23214 31714 23266 31726
rect 14366 31666 14418 31678
rect 25554 31614 25566 31666
rect 25618 31614 25630 31666
rect 14366 31602 14418 31614
rect 22654 31554 22706 31566
rect 22654 31490 22706 31502
rect 1344 31386 38640 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 38640 31386
rect 1344 31300 38640 31334
rect 20750 31218 20802 31230
rect 25454 31218 25506 31230
rect 22866 31166 22878 31218
rect 22930 31166 22942 31218
rect 20750 31154 20802 31166
rect 25454 31154 25506 31166
rect 26126 31218 26178 31230
rect 26126 31154 26178 31166
rect 21870 31106 21922 31118
rect 12114 31054 12126 31106
rect 12178 31054 12190 31106
rect 18162 31054 18174 31106
rect 18226 31054 18238 31106
rect 21870 31042 21922 31054
rect 38222 31106 38274 31118
rect 38222 31042 38274 31054
rect 14702 30994 14754 31006
rect 23214 30994 23266 31006
rect 24670 30994 24722 31006
rect 11442 30942 11454 30994
rect 11506 30942 11518 30994
rect 17490 30942 17502 30994
rect 17554 30942 17566 30994
rect 23986 30942 23998 30994
rect 24050 30942 24062 30994
rect 14702 30930 14754 30942
rect 23214 30930 23266 30942
rect 24670 30930 24722 30942
rect 25230 30994 25282 31006
rect 25230 30930 25282 30942
rect 14242 30830 14254 30882
rect 14306 30830 14318 30882
rect 20290 30830 20302 30882
rect 20354 30830 20366 30882
rect 24210 30830 24222 30882
rect 24274 30830 24286 30882
rect 25554 30830 25566 30882
rect 25618 30830 25630 30882
rect 21982 30770 22034 30782
rect 21982 30706 22034 30718
rect 1344 30602 38640 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 38640 30602
rect 1344 30516 38640 30550
rect 20862 30322 20914 30334
rect 22082 30270 22094 30322
rect 22146 30270 22158 30322
rect 24210 30270 24222 30322
rect 24274 30270 24286 30322
rect 20862 30258 20914 30270
rect 21298 30158 21310 30210
rect 21362 30158 21374 30210
rect 1344 29818 38640 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 38640 29818
rect 1344 29732 38640 29766
rect 1344 29034 38640 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 38640 29034
rect 1344 28948 38640 28982
rect 1344 28250 38640 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 38640 28250
rect 1344 28164 38640 28198
rect 1344 27466 38640 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 38640 27466
rect 1344 27380 38640 27414
rect 1344 26682 38640 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 38640 26682
rect 1344 26596 38640 26630
rect 1344 25898 38640 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 38640 25898
rect 1344 25812 38640 25846
rect 1344 25114 38640 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 38640 25114
rect 1344 25028 38640 25062
rect 1344 24330 38640 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 38640 24330
rect 1344 24244 38640 24278
rect 1344 23546 38640 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 38640 23546
rect 1344 23460 38640 23494
rect 38222 23266 38274 23278
rect 38222 23202 38274 23214
rect 1344 22762 38640 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 38640 22762
rect 1344 22676 38640 22710
rect 1344 21978 38640 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 38640 21978
rect 1344 21892 38640 21926
rect 1344 21194 38640 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 38640 21194
rect 1344 21108 38640 21142
rect 1344 20410 38640 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 38640 20410
rect 1344 20324 38640 20358
rect 1344 19626 38640 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 38640 19626
rect 1344 19540 38640 19574
rect 1344 18842 38640 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 38640 18842
rect 1344 18756 38640 18790
rect 1344 18058 38640 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 38640 18058
rect 1344 17972 38640 18006
rect 1344 17274 38640 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 38640 17274
rect 1344 17188 38640 17222
rect 1344 16490 38640 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 38640 16490
rect 1344 16404 38640 16438
rect 1344 15706 38640 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 38640 15706
rect 1344 15620 38640 15654
rect 1344 14922 38640 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 38640 14922
rect 1344 14836 38640 14870
rect 1344 14138 38640 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 38640 14138
rect 1344 14052 38640 14086
rect 1344 13354 38640 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 38640 13354
rect 1344 13268 38640 13302
rect 1344 12570 38640 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 38640 12570
rect 1344 12484 38640 12518
rect 1344 11786 38640 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 38640 11786
rect 1344 11700 38640 11734
rect 1344 11002 38640 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 38640 11002
rect 1344 10916 38640 10950
rect 1344 10218 38640 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 38640 10218
rect 1344 10132 38640 10166
rect 1344 9434 38640 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 38640 9434
rect 1344 9348 38640 9382
rect 1344 8650 38640 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 38640 8650
rect 1344 8564 38640 8598
rect 1344 7866 38640 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 38640 7866
rect 1344 7780 38640 7814
rect 1344 7082 38640 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 38640 7082
rect 1344 6996 38640 7030
rect 1344 6298 38640 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 38640 6298
rect 1344 6212 38640 6246
rect 1344 5514 38640 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 38640 5514
rect 1344 5428 38640 5462
rect 1344 4730 38640 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 38640 4730
rect 1344 4644 38640 4678
rect 1344 3946 38640 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 38640 3946
rect 1344 3860 38640 3894
rect 2942 3330 2994 3342
rect 2942 3266 2994 3278
rect 1344 3162 38640 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 38640 3162
rect 1344 3076 38640 3110
<< via1 >>
rect 4478 96406 4530 96458
rect 4582 96406 4634 96458
rect 4686 96406 4738 96458
rect 35198 96406 35250 96458
rect 35302 96406 35354 96458
rect 35406 96406 35458 96458
rect 3614 95902 3666 95954
rect 19838 95622 19890 95674
rect 19942 95622 19994 95674
rect 20046 95622 20098 95674
rect 4478 94838 4530 94890
rect 4582 94838 4634 94890
rect 4686 94838 4738 94890
rect 35198 94838 35250 94890
rect 35302 94838 35354 94890
rect 35406 94838 35458 94890
rect 19838 94054 19890 94106
rect 19942 94054 19994 94106
rect 20046 94054 20098 94106
rect 4478 93270 4530 93322
rect 4582 93270 4634 93322
rect 4686 93270 4738 93322
rect 35198 93270 35250 93322
rect 35302 93270 35354 93322
rect 35406 93270 35458 93322
rect 19838 92486 19890 92538
rect 19942 92486 19994 92538
rect 20046 92486 20098 92538
rect 4478 91702 4530 91754
rect 4582 91702 4634 91754
rect 4686 91702 4738 91754
rect 35198 91702 35250 91754
rect 35302 91702 35354 91754
rect 35406 91702 35458 91754
rect 19838 90918 19890 90970
rect 19942 90918 19994 90970
rect 20046 90918 20098 90970
rect 4478 90134 4530 90186
rect 4582 90134 4634 90186
rect 4686 90134 4738 90186
rect 35198 90134 35250 90186
rect 35302 90134 35354 90186
rect 35406 90134 35458 90186
rect 19838 89350 19890 89402
rect 19942 89350 19994 89402
rect 20046 89350 20098 89402
rect 4478 88566 4530 88618
rect 4582 88566 4634 88618
rect 4686 88566 4738 88618
rect 35198 88566 35250 88618
rect 35302 88566 35354 88618
rect 35406 88566 35458 88618
rect 19838 87782 19890 87834
rect 19942 87782 19994 87834
rect 20046 87782 20098 87834
rect 4478 86998 4530 87050
rect 4582 86998 4634 87050
rect 4686 86998 4738 87050
rect 35198 86998 35250 87050
rect 35302 86998 35354 87050
rect 35406 86998 35458 87050
rect 19838 86214 19890 86266
rect 19942 86214 19994 86266
rect 20046 86214 20098 86266
rect 4478 85430 4530 85482
rect 4582 85430 4634 85482
rect 4686 85430 4738 85482
rect 35198 85430 35250 85482
rect 35302 85430 35354 85482
rect 35406 85430 35458 85482
rect 19838 84646 19890 84698
rect 19942 84646 19994 84698
rect 20046 84646 20098 84698
rect 4478 83862 4530 83914
rect 4582 83862 4634 83914
rect 4686 83862 4738 83914
rect 35198 83862 35250 83914
rect 35302 83862 35354 83914
rect 35406 83862 35458 83914
rect 19838 83078 19890 83130
rect 19942 83078 19994 83130
rect 20046 83078 20098 83130
rect 4478 82294 4530 82346
rect 4582 82294 4634 82346
rect 4686 82294 4738 82346
rect 35198 82294 35250 82346
rect 35302 82294 35354 82346
rect 35406 82294 35458 82346
rect 19838 81510 19890 81562
rect 19942 81510 19994 81562
rect 20046 81510 20098 81562
rect 4478 80726 4530 80778
rect 4582 80726 4634 80778
rect 4686 80726 4738 80778
rect 35198 80726 35250 80778
rect 35302 80726 35354 80778
rect 35406 80726 35458 80778
rect 19838 79942 19890 79994
rect 19942 79942 19994 79994
rect 20046 79942 20098 79994
rect 4478 79158 4530 79210
rect 4582 79158 4634 79210
rect 4686 79158 4738 79210
rect 35198 79158 35250 79210
rect 35302 79158 35354 79210
rect 35406 79158 35458 79210
rect 19838 78374 19890 78426
rect 19942 78374 19994 78426
rect 20046 78374 20098 78426
rect 4478 77590 4530 77642
rect 4582 77590 4634 77642
rect 4686 77590 4738 77642
rect 35198 77590 35250 77642
rect 35302 77590 35354 77642
rect 35406 77590 35458 77642
rect 19838 76806 19890 76858
rect 19942 76806 19994 76858
rect 20046 76806 20098 76858
rect 4478 76022 4530 76074
rect 4582 76022 4634 76074
rect 4686 76022 4738 76074
rect 35198 76022 35250 76074
rect 35302 76022 35354 76074
rect 35406 76022 35458 76074
rect 19838 75238 19890 75290
rect 19942 75238 19994 75290
rect 20046 75238 20098 75290
rect 4478 74454 4530 74506
rect 4582 74454 4634 74506
rect 4686 74454 4738 74506
rect 35198 74454 35250 74506
rect 35302 74454 35354 74506
rect 35406 74454 35458 74506
rect 19838 73670 19890 73722
rect 19942 73670 19994 73722
rect 20046 73670 20098 73722
rect 4478 72886 4530 72938
rect 4582 72886 4634 72938
rect 4686 72886 4738 72938
rect 35198 72886 35250 72938
rect 35302 72886 35354 72938
rect 35406 72886 35458 72938
rect 19838 72102 19890 72154
rect 19942 72102 19994 72154
rect 20046 72102 20098 72154
rect 4478 71318 4530 71370
rect 4582 71318 4634 71370
rect 4686 71318 4738 71370
rect 35198 71318 35250 71370
rect 35302 71318 35354 71370
rect 35406 71318 35458 71370
rect 19838 70534 19890 70586
rect 19942 70534 19994 70586
rect 20046 70534 20098 70586
rect 25342 70254 25394 70306
rect 17950 70142 18002 70194
rect 19854 70142 19906 70194
rect 20078 70142 20130 70194
rect 20190 70142 20242 70194
rect 25566 70030 25618 70082
rect 26126 70030 26178 70082
rect 18174 69918 18226 69970
rect 18398 69918 18450 69970
rect 18510 69918 18562 69970
rect 20638 69918 20690 69970
rect 25230 69918 25282 69970
rect 4478 69750 4530 69802
rect 4582 69750 4634 69802
rect 4686 69750 4738 69802
rect 35198 69750 35250 69802
rect 35302 69750 35354 69802
rect 35406 69750 35458 69802
rect 20638 69582 20690 69634
rect 20414 69470 20466 69522
rect 22318 69470 22370 69522
rect 24446 69470 24498 69522
rect 15262 69358 15314 69410
rect 16606 69358 16658 69410
rect 17838 69358 17890 69410
rect 18398 69358 18450 69410
rect 19070 69358 19122 69410
rect 20190 69358 20242 69410
rect 25230 69358 25282 69410
rect 25566 69358 25618 69410
rect 19630 69246 19682 69298
rect 20750 69246 20802 69298
rect 25790 69246 25842 69298
rect 25902 69246 25954 69298
rect 15822 69134 15874 69186
rect 16830 69134 16882 69186
rect 26350 69134 26402 69186
rect 19838 68966 19890 69018
rect 19942 68966 19994 69018
rect 20046 68966 20098 69018
rect 17614 68798 17666 68850
rect 2046 68686 2098 68738
rect 9662 68686 9714 68738
rect 9774 68686 9826 68738
rect 17390 68686 17442 68738
rect 24670 68686 24722 68738
rect 25230 68686 25282 68738
rect 25790 68686 25842 68738
rect 1710 68574 1762 68626
rect 10334 68574 10386 68626
rect 13694 68574 13746 68626
rect 18510 68574 18562 68626
rect 18958 68574 19010 68626
rect 19630 68574 19682 68626
rect 23998 68574 24050 68626
rect 24334 68574 24386 68626
rect 25454 68574 25506 68626
rect 28926 68574 28978 68626
rect 2494 68462 2546 68514
rect 11006 68462 11058 68514
rect 13246 68462 13298 68514
rect 14478 68462 14530 68514
rect 16606 68462 16658 68514
rect 17726 68462 17778 68514
rect 21086 68462 21138 68514
rect 23214 68462 23266 68514
rect 25678 68462 25730 68514
rect 26126 68462 26178 68514
rect 28254 68462 28306 68514
rect 9774 68350 9826 68402
rect 20190 68350 20242 68402
rect 4478 68182 4530 68234
rect 4582 68182 4634 68234
rect 4686 68182 4738 68234
rect 35198 68182 35250 68234
rect 35302 68182 35354 68234
rect 35406 68182 35458 68234
rect 7646 67902 7698 67954
rect 11006 67902 11058 67954
rect 19630 67902 19682 67954
rect 20526 67902 20578 67954
rect 24558 67902 24610 67954
rect 28590 67902 28642 67954
rect 10558 67790 10610 67842
rect 10782 67790 10834 67842
rect 11790 67790 11842 67842
rect 12126 67790 12178 67842
rect 12574 67790 12626 67842
rect 14142 67790 14194 67842
rect 15486 67790 15538 67842
rect 17726 67790 17778 67842
rect 20078 67790 20130 67842
rect 23550 67790 23602 67842
rect 24670 67790 24722 67842
rect 25790 67790 25842 67842
rect 1710 67678 1762 67730
rect 9774 67678 9826 67730
rect 11230 67678 11282 67730
rect 11454 67678 11506 67730
rect 12350 67678 12402 67730
rect 12910 67678 12962 67730
rect 16718 67678 16770 67730
rect 18174 67678 18226 67730
rect 23886 67678 23938 67730
rect 24222 67678 24274 67730
rect 26462 67678 26514 67730
rect 2046 67566 2098 67618
rect 2494 67566 2546 67618
rect 11902 67566 11954 67618
rect 12798 67566 12850 67618
rect 13582 67566 13634 67618
rect 14478 67566 14530 67618
rect 16270 67566 16322 67618
rect 19838 67398 19890 67450
rect 19942 67398 19994 67450
rect 20046 67398 20098 67450
rect 9774 67230 9826 67282
rect 13918 67230 13970 67282
rect 23214 67230 23266 67282
rect 2046 67118 2098 67170
rect 8206 67118 8258 67170
rect 8318 67118 8370 67170
rect 8542 67118 8594 67170
rect 8766 67118 8818 67170
rect 8878 67118 8930 67170
rect 10110 67118 10162 67170
rect 11678 67118 11730 67170
rect 16830 67118 16882 67170
rect 17390 67118 17442 67170
rect 20190 67118 20242 67170
rect 25454 67118 25506 67170
rect 25566 67118 25618 67170
rect 26462 67118 26514 67170
rect 27582 67118 27634 67170
rect 1710 67006 1762 67058
rect 9102 67006 9154 67058
rect 9438 67006 9490 67058
rect 9774 67006 9826 67058
rect 10894 67006 10946 67058
rect 17838 67006 17890 67058
rect 18062 67006 18114 67058
rect 20414 67006 20466 67058
rect 21310 67006 21362 67058
rect 22990 67006 23042 67058
rect 25230 67006 25282 67058
rect 25790 67006 25842 67058
rect 26238 67006 26290 67058
rect 26798 67006 26850 67058
rect 27022 67006 27074 67058
rect 27470 67006 27522 67058
rect 2494 66894 2546 66946
rect 18622 66894 18674 66946
rect 21422 66894 21474 66946
rect 16718 66782 16770 66834
rect 17614 66782 17666 66834
rect 21198 66782 21250 66834
rect 26574 66782 26626 66834
rect 27358 66782 27410 66834
rect 4478 66614 4530 66666
rect 4582 66614 4634 66666
rect 4686 66614 4738 66666
rect 35198 66614 35250 66666
rect 35302 66614 35354 66666
rect 35406 66614 35458 66666
rect 26462 66446 26514 66498
rect 26798 66446 26850 66498
rect 9886 66222 9938 66274
rect 10222 66222 10274 66274
rect 12574 66222 12626 66274
rect 12910 66222 12962 66274
rect 26238 66222 26290 66274
rect 26686 66222 26738 66274
rect 9662 65998 9714 66050
rect 9998 65998 10050 66050
rect 12350 65998 12402 66050
rect 12798 65998 12850 66050
rect 27246 65998 27298 66050
rect 19838 65830 19890 65882
rect 19942 65830 19994 65882
rect 20046 65830 20098 65882
rect 24334 65550 24386 65602
rect 23886 65438 23938 65490
rect 24446 65438 24498 65490
rect 24670 65438 24722 65490
rect 2158 65326 2210 65378
rect 25342 65326 25394 65378
rect 25790 65326 25842 65378
rect 4478 65046 4530 65098
rect 4582 65046 4634 65098
rect 4686 65046 4738 65098
rect 35198 65046 35250 65098
rect 35302 65046 35354 65098
rect 35406 65046 35458 65098
rect 1822 64654 1874 64706
rect 9326 64654 9378 64706
rect 14030 64654 14082 64706
rect 14142 64654 14194 64706
rect 14478 64654 14530 64706
rect 2382 64542 2434 64594
rect 2718 64542 2770 64594
rect 8654 64542 8706 64594
rect 8766 64542 8818 64594
rect 9998 64542 10050 64594
rect 13694 64542 13746 64594
rect 2046 64430 2098 64482
rect 3166 64430 3218 64482
rect 8990 64430 9042 64482
rect 12686 64430 12738 64482
rect 14142 64430 14194 64482
rect 25678 64430 25730 64482
rect 38222 64430 38274 64482
rect 19838 64262 19890 64314
rect 19942 64262 19994 64314
rect 20046 64262 20098 64314
rect 9998 64094 10050 64146
rect 10446 64094 10498 64146
rect 11118 64094 11170 64146
rect 11342 64094 11394 64146
rect 13358 64094 13410 64146
rect 14478 64094 14530 64146
rect 2046 63982 2098 64034
rect 10670 63982 10722 64034
rect 13918 63982 13970 64034
rect 14590 63982 14642 64034
rect 17950 63982 18002 64034
rect 20190 63982 20242 64034
rect 26238 63982 26290 64034
rect 1710 63870 1762 63922
rect 2494 63870 2546 63922
rect 9774 63870 9826 63922
rect 10222 63870 10274 63922
rect 10894 63870 10946 63922
rect 11454 63870 11506 63922
rect 18286 63870 18338 63922
rect 18958 63870 19010 63922
rect 24334 63870 24386 63922
rect 25790 63870 25842 63922
rect 26798 63870 26850 63922
rect 13694 63758 13746 63810
rect 13806 63758 13858 63810
rect 19630 63758 19682 63810
rect 21422 63758 21474 63810
rect 23550 63758 23602 63810
rect 25566 63758 25618 63810
rect 27470 63758 27522 63810
rect 29598 63758 29650 63810
rect 14366 63646 14418 63698
rect 19966 63646 20018 63698
rect 20302 63646 20354 63698
rect 25230 63646 25282 63698
rect 4478 63478 4530 63530
rect 4582 63478 4634 63530
rect 4686 63478 4738 63530
rect 35198 63478 35250 63530
rect 35302 63478 35354 63530
rect 35406 63478 35458 63530
rect 18062 63310 18114 63362
rect 27470 63198 27522 63250
rect 9886 63086 9938 63138
rect 13582 63086 13634 63138
rect 17390 63086 17442 63138
rect 17838 63086 17890 63138
rect 19406 63086 19458 63138
rect 20302 63086 20354 63138
rect 22766 63086 22818 63138
rect 23326 63086 23378 63138
rect 24670 63086 24722 63138
rect 24894 63086 24946 63138
rect 25230 63086 25282 63138
rect 26014 63086 26066 63138
rect 26238 63086 26290 63138
rect 27582 63086 27634 63138
rect 28030 63086 28082 63138
rect 1710 62974 1762 63026
rect 2046 62974 2098 63026
rect 8878 62974 8930 63026
rect 8990 62974 9042 63026
rect 14254 62974 14306 63026
rect 17278 62974 17330 63026
rect 18846 62974 18898 63026
rect 23662 62974 23714 63026
rect 23998 62974 24050 63026
rect 24222 62974 24274 63026
rect 25006 62974 25058 63026
rect 26910 62974 26962 63026
rect 27246 62974 27298 63026
rect 2494 62862 2546 62914
rect 9214 62862 9266 62914
rect 10222 62862 10274 62914
rect 16494 62862 16546 62914
rect 18174 62862 18226 62914
rect 20414 62862 20466 62914
rect 19838 62694 19890 62746
rect 19942 62694 19994 62746
rect 20046 62694 20098 62746
rect 8094 62526 8146 62578
rect 13246 62526 13298 62578
rect 14254 62526 14306 62578
rect 14702 62526 14754 62578
rect 16046 62526 16098 62578
rect 16830 62526 16882 62578
rect 17502 62526 17554 62578
rect 24334 62526 24386 62578
rect 14142 62414 14194 62466
rect 15710 62414 15762 62466
rect 19518 62414 19570 62466
rect 20190 62414 20242 62466
rect 21534 62414 21586 62466
rect 24558 62414 24610 62466
rect 24670 62414 24722 62466
rect 7870 62302 7922 62354
rect 8542 62302 8594 62354
rect 8766 62302 8818 62354
rect 9102 62302 9154 62354
rect 9550 62302 9602 62354
rect 13694 62302 13746 62354
rect 14366 62302 14418 62354
rect 14926 62302 14978 62354
rect 15598 62302 15650 62354
rect 17614 62302 17666 62354
rect 17950 62302 18002 62354
rect 18958 62302 19010 62354
rect 19294 62302 19346 62354
rect 24222 62302 24274 62354
rect 29038 62302 29090 62354
rect 8878 62190 8930 62242
rect 10334 62190 10386 62242
rect 12462 62190 12514 62242
rect 19966 62190 20018 62242
rect 22094 62190 22146 62242
rect 28478 62190 28530 62242
rect 13918 62078 13970 62130
rect 19630 62078 19682 62130
rect 4478 61910 4530 61962
rect 4582 61910 4634 61962
rect 4686 61910 4738 61962
rect 35198 61910 35250 61962
rect 35302 61910 35354 61962
rect 35406 61910 35458 61962
rect 19742 61742 19794 61794
rect 23886 61630 23938 61682
rect 27134 61630 27186 61682
rect 8430 61518 8482 61570
rect 8878 61518 8930 61570
rect 9550 61518 9602 61570
rect 10110 61518 10162 61570
rect 13582 61518 13634 61570
rect 19294 61518 19346 61570
rect 19630 61518 19682 61570
rect 20190 61518 20242 61570
rect 20414 61518 20466 61570
rect 23998 61518 24050 61570
rect 24670 61518 24722 61570
rect 24894 61518 24946 61570
rect 25230 61518 25282 61570
rect 26910 61518 26962 61570
rect 10446 61406 10498 61458
rect 13806 61406 13858 61458
rect 18734 61406 18786 61458
rect 18958 61406 19010 61458
rect 9214 61294 9266 61346
rect 10334 61294 10386 61346
rect 19070 61294 19122 61346
rect 19742 61350 19794 61402
rect 20750 61406 20802 61458
rect 23326 61406 23378 61458
rect 25790 61406 25842 61458
rect 27022 61406 27074 61458
rect 20414 61294 20466 61346
rect 23214 61294 23266 61346
rect 24446 61294 24498 61346
rect 24782 61294 24834 61346
rect 19838 61126 19890 61178
rect 19942 61126 19994 61178
rect 20046 61126 20098 61178
rect 22206 60958 22258 61010
rect 18398 60846 18450 60898
rect 16830 60734 16882 60786
rect 18734 60734 18786 60786
rect 19518 60734 19570 60786
rect 20638 60734 20690 60786
rect 20862 60734 20914 60786
rect 21086 60734 21138 60786
rect 28478 60734 28530 60786
rect 11790 60622 11842 60674
rect 17502 60622 17554 60674
rect 20078 60622 20130 60674
rect 22654 60622 22706 60674
rect 25678 60622 25730 60674
rect 27806 60622 27858 60674
rect 21310 60510 21362 60562
rect 21758 60510 21810 60562
rect 4478 60342 4530 60394
rect 4582 60342 4634 60394
rect 4686 60342 4738 60394
rect 35198 60342 35250 60394
rect 35302 60342 35354 60394
rect 35406 60342 35458 60394
rect 19070 60174 19122 60226
rect 19742 60174 19794 60226
rect 19854 60174 19906 60226
rect 6078 59950 6130 60002
rect 14814 59950 14866 60002
rect 18510 59950 18562 60002
rect 19294 59950 19346 60002
rect 19630 59950 19682 60002
rect 24782 59950 24834 60002
rect 25342 59950 25394 60002
rect 1710 59838 1762 59890
rect 2494 59838 2546 59890
rect 6750 59838 6802 59890
rect 13470 59838 13522 59890
rect 14478 59838 14530 59890
rect 15934 59838 15986 59890
rect 17390 59838 17442 59890
rect 24894 59838 24946 59890
rect 25118 59838 25170 59890
rect 25790 59838 25842 59890
rect 26238 59838 26290 59890
rect 26574 59838 26626 59890
rect 2046 59726 2098 59778
rect 8990 59726 9042 59778
rect 13582 59726 13634 59778
rect 13694 59726 13746 59778
rect 14366 59726 14418 59778
rect 15822 59726 15874 59778
rect 24446 59726 24498 59778
rect 19838 59558 19890 59610
rect 19942 59558 19994 59610
rect 20046 59558 20098 59610
rect 7982 59390 8034 59442
rect 11118 59390 11170 59442
rect 16270 59390 16322 59442
rect 18174 59390 18226 59442
rect 18846 59390 18898 59442
rect 9662 59278 9714 59330
rect 11454 59278 11506 59330
rect 17502 59278 17554 59330
rect 17726 59278 17778 59330
rect 7870 59166 7922 59218
rect 8206 59166 8258 59218
rect 8430 59166 8482 59218
rect 9438 59166 9490 59218
rect 9774 59166 9826 59218
rect 12238 59166 12290 59218
rect 16830 59166 16882 59218
rect 17614 59166 17666 59218
rect 18510 59166 18562 59218
rect 12910 59054 12962 59106
rect 15038 59054 15090 59106
rect 25902 59054 25954 59106
rect 4478 58774 4530 58826
rect 4582 58774 4634 58826
rect 4686 58774 4738 58826
rect 35198 58774 35250 58826
rect 35302 58774 35354 58826
rect 35406 58774 35458 58826
rect 13694 58606 13746 58658
rect 25902 58606 25954 58658
rect 18174 58494 18226 58546
rect 25566 58494 25618 58546
rect 26910 58494 26962 58546
rect 27582 58494 27634 58546
rect 10110 58382 10162 58434
rect 13582 58382 13634 58434
rect 14030 58382 14082 58434
rect 14254 58382 14306 58434
rect 16270 58382 16322 58434
rect 17502 58382 17554 58434
rect 17838 58382 17890 58434
rect 25678 58382 25730 58434
rect 1710 58270 1762 58322
rect 10334 58270 10386 58322
rect 16718 58270 16770 58322
rect 18398 58270 18450 58322
rect 24782 58270 24834 58322
rect 27246 58270 27298 58322
rect 27470 58270 27522 58322
rect 2046 58158 2098 58210
rect 2494 58158 2546 58210
rect 9774 58158 9826 58210
rect 13470 58158 13522 58210
rect 18958 58158 19010 58210
rect 25118 58158 25170 58210
rect 25566 58158 25618 58210
rect 19838 57990 19890 58042
rect 19942 57990 19994 58042
rect 20046 57990 20098 58042
rect 8094 57822 8146 57874
rect 2046 57710 2098 57762
rect 7758 57710 7810 57762
rect 7870 57710 7922 57762
rect 9886 57710 9938 57762
rect 13022 57710 13074 57762
rect 15822 57710 15874 57762
rect 16158 57710 16210 57762
rect 17614 57710 17666 57762
rect 23662 57710 23714 57762
rect 1710 57598 1762 57650
rect 10222 57598 10274 57650
rect 13358 57598 13410 57650
rect 17726 57598 17778 57650
rect 24446 57598 24498 57650
rect 26014 57598 26066 57650
rect 2494 57486 2546 57538
rect 15038 57486 15090 57538
rect 18622 57486 18674 57538
rect 21534 57486 21586 57538
rect 25678 57486 25730 57538
rect 13358 57374 13410 57426
rect 16382 57374 16434 57426
rect 16718 57374 16770 57426
rect 25678 57374 25730 57426
rect 26014 57486 26066 57538
rect 28478 57486 28530 57538
rect 4478 57206 4530 57258
rect 4582 57206 4634 57258
rect 4686 57206 4738 57258
rect 35198 57206 35250 57258
rect 35302 57206 35354 57258
rect 35406 57206 35458 57258
rect 13694 57038 13746 57090
rect 25342 57038 25394 57090
rect 27246 57038 27298 57090
rect 28030 57038 28082 57090
rect 17502 56926 17554 56978
rect 18062 56926 18114 56978
rect 21422 56926 21474 56978
rect 13470 56814 13522 56866
rect 14030 56814 14082 56866
rect 16718 56814 16770 56866
rect 17614 56814 17666 56866
rect 21870 56814 21922 56866
rect 22654 56814 22706 56866
rect 23662 56814 23714 56866
rect 24446 56814 24498 56866
rect 24670 56814 24722 56866
rect 25118 56814 25170 56866
rect 26910 56814 26962 56866
rect 27358 56814 27410 56866
rect 28254 56814 28306 56866
rect 28366 56814 28418 56866
rect 1710 56702 1762 56754
rect 7422 56702 7474 56754
rect 7758 56702 7810 56754
rect 7982 56702 8034 56754
rect 8318 56702 8370 56754
rect 8542 56702 8594 56754
rect 12350 56702 12402 56754
rect 14254 56702 14306 56754
rect 15598 56702 15650 56754
rect 16270 56702 16322 56754
rect 22318 56702 22370 56754
rect 24782 56702 24834 56754
rect 27918 56702 27970 56754
rect 2046 56590 2098 56642
rect 2494 56590 2546 56642
rect 7534 56590 7586 56642
rect 8094 56590 8146 56642
rect 12014 56590 12066 56642
rect 13470 56590 13522 56642
rect 15486 56590 15538 56642
rect 17166 56590 17218 56642
rect 17390 56590 17442 56642
rect 22766 56590 22818 56642
rect 23102 56590 23154 56642
rect 25678 56590 25730 56642
rect 19838 56422 19890 56474
rect 19942 56422 19994 56474
rect 20046 56422 20098 56474
rect 2046 56254 2098 56306
rect 17614 56254 17666 56306
rect 10110 56142 10162 56194
rect 24558 56142 24610 56194
rect 27806 56142 27858 56194
rect 1710 56030 1762 56082
rect 5966 56030 6018 56082
rect 9438 56030 9490 56082
rect 9774 56030 9826 56082
rect 16606 56030 16658 56082
rect 17502 56030 17554 56082
rect 17838 56030 17890 56082
rect 18062 56030 18114 56082
rect 18398 56030 18450 56082
rect 21758 56030 21810 56082
rect 24446 56030 24498 56082
rect 24782 56030 24834 56082
rect 25342 56030 25394 56082
rect 25566 56030 25618 56082
rect 25902 56030 25954 56082
rect 27134 56030 27186 56082
rect 2494 55918 2546 55970
rect 6638 55918 6690 55970
rect 8766 55918 8818 55970
rect 9662 55918 9714 55970
rect 12014 55918 12066 55970
rect 17726 55918 17778 55970
rect 18958 55918 19010 55970
rect 21086 55918 21138 55970
rect 21422 55918 21474 55970
rect 29934 55918 29986 55970
rect 25790 55806 25842 55858
rect 4478 55638 4530 55690
rect 4582 55638 4634 55690
rect 4686 55638 4738 55690
rect 35198 55638 35250 55690
rect 35302 55638 35354 55690
rect 35406 55638 35458 55690
rect 22206 55470 22258 55522
rect 9102 55358 9154 55410
rect 11566 55358 11618 55410
rect 17278 55358 17330 55410
rect 21982 55358 22034 55410
rect 27694 55358 27746 55410
rect 29262 55358 29314 55410
rect 6302 55246 6354 55298
rect 9326 55246 9378 55298
rect 9662 55246 9714 55298
rect 10558 55246 10610 55298
rect 15038 55246 15090 55298
rect 15598 55246 15650 55298
rect 18398 55246 18450 55298
rect 22094 55246 22146 55298
rect 26350 55246 26402 55298
rect 26910 55246 26962 55298
rect 29038 55246 29090 55298
rect 29374 55246 29426 55298
rect 29598 55246 29650 55298
rect 1710 55134 1762 55186
rect 2046 55134 2098 55186
rect 2494 55134 2546 55186
rect 6974 55134 7026 55186
rect 10334 55134 10386 55186
rect 11902 55134 11954 55186
rect 12910 55134 12962 55186
rect 17166 55134 17218 55186
rect 18174 55134 18226 55186
rect 19182 55134 19234 55186
rect 25342 55134 25394 55186
rect 27358 55134 27410 55186
rect 9550 55022 9602 55074
rect 11006 55022 11058 55074
rect 12238 55022 12290 55074
rect 12574 55022 12626 55074
rect 15262 55022 15314 55074
rect 19294 55022 19346 55074
rect 19838 54854 19890 54906
rect 19942 54854 19994 54906
rect 20046 54854 20098 54906
rect 8094 54686 8146 54738
rect 9102 54686 9154 54738
rect 9774 54686 9826 54738
rect 10110 54686 10162 54738
rect 14926 54686 14978 54738
rect 7758 54574 7810 54626
rect 7870 54574 7922 54626
rect 8878 54574 8930 54626
rect 12686 54574 12738 54626
rect 16606 54574 16658 54626
rect 18846 54574 18898 54626
rect 25454 54574 25506 54626
rect 27806 54574 27858 54626
rect 8766 54462 8818 54514
rect 12014 54462 12066 54514
rect 17614 54462 17666 54514
rect 20078 54462 20130 54514
rect 27134 54462 27186 54514
rect 35982 54462 36034 54514
rect 17726 54350 17778 54402
rect 18174 54350 18226 54402
rect 18734 54350 18786 54402
rect 20750 54350 20802 54402
rect 25342 54350 25394 54402
rect 29934 54350 29986 54402
rect 16046 54238 16098 54290
rect 25230 54238 25282 54290
rect 37998 54238 38050 54290
rect 4478 54070 4530 54122
rect 4582 54070 4634 54122
rect 4686 54070 4738 54122
rect 35198 54070 35250 54122
rect 35302 54070 35354 54122
rect 35406 54070 35458 54122
rect 27582 53902 27634 53954
rect 19406 53790 19458 53842
rect 27246 53790 27298 53842
rect 16942 53678 16994 53730
rect 17390 53678 17442 53730
rect 19182 53678 19234 53730
rect 21310 53678 21362 53730
rect 21982 53678 22034 53730
rect 22430 53678 22482 53730
rect 24446 53678 24498 53730
rect 26910 53678 26962 53730
rect 16382 53566 16434 53618
rect 17838 53566 17890 53618
rect 21534 53566 21586 53618
rect 22542 53566 22594 53618
rect 25006 53566 25058 53618
rect 1710 53454 1762 53506
rect 2046 53454 2098 53506
rect 2494 53454 2546 53506
rect 15934 53454 15986 53506
rect 19518 53454 19570 53506
rect 19742 53454 19794 53506
rect 21758 53454 21810 53506
rect 23998 53454 24050 53506
rect 26798 53454 26850 53506
rect 27358 53454 27410 53506
rect 19838 53286 19890 53338
rect 19942 53286 19994 53338
rect 20046 53286 20098 53338
rect 10334 53118 10386 53170
rect 17502 53118 17554 53170
rect 17726 53118 17778 53170
rect 15262 53006 15314 53058
rect 18734 53006 18786 53058
rect 21310 53006 21362 53058
rect 22990 53006 23042 53058
rect 24670 53006 24722 53058
rect 14814 52894 14866 52946
rect 15038 52894 15090 52946
rect 16606 52894 16658 52946
rect 17390 52894 17442 52946
rect 18510 52894 18562 52946
rect 19406 52894 19458 52946
rect 19742 52894 19794 52946
rect 21870 52894 21922 52946
rect 22318 52894 22370 52946
rect 24110 52894 24162 52946
rect 25902 52894 25954 52946
rect 33070 52894 33122 52946
rect 10222 52782 10274 52834
rect 16270 52782 16322 52834
rect 20974 52782 21026 52834
rect 22206 52782 22258 52834
rect 24222 52782 24274 52834
rect 26574 52782 26626 52834
rect 28702 52782 28754 52834
rect 33854 52782 33906 52834
rect 35982 52782 36034 52834
rect 15374 52670 15426 52722
rect 4478 52502 4530 52554
rect 4582 52502 4634 52554
rect 4686 52502 4738 52554
rect 35198 52502 35250 52554
rect 35302 52502 35354 52554
rect 35406 52502 35458 52554
rect 12462 52334 12514 52386
rect 26574 52334 26626 52386
rect 26686 52334 26738 52386
rect 26910 52334 26962 52386
rect 27358 52334 27410 52386
rect 27582 52334 27634 52386
rect 11790 52222 11842 52274
rect 15710 52222 15762 52274
rect 16718 52222 16770 52274
rect 18398 52222 18450 52274
rect 27582 52222 27634 52274
rect 1710 52110 1762 52162
rect 2494 52110 2546 52162
rect 11454 52110 11506 52162
rect 12126 52110 12178 52162
rect 15486 52110 15538 52162
rect 18174 52110 18226 52162
rect 20190 52110 20242 52162
rect 21870 52110 21922 52162
rect 23886 52110 23938 52162
rect 27134 52110 27186 52162
rect 33742 52110 33794 52162
rect 2046 51998 2098 52050
rect 12686 51998 12738 52050
rect 12910 51998 12962 52050
rect 17950 51998 18002 52050
rect 18622 51998 18674 52050
rect 21982 51998 22034 52050
rect 24446 51998 24498 52050
rect 34078 51998 34130 52050
rect 11678 51886 11730 51938
rect 12462 51886 12514 51938
rect 23438 51886 23490 51938
rect 19838 51718 19890 51770
rect 19942 51718 19994 51770
rect 20046 51718 20098 51770
rect 10222 51550 10274 51602
rect 15598 51550 15650 51602
rect 16046 51550 16098 51602
rect 23326 51550 23378 51602
rect 26574 51550 26626 51602
rect 2046 51438 2098 51490
rect 9550 51438 9602 51490
rect 10558 51438 10610 51490
rect 12462 51438 12514 51490
rect 16606 51438 16658 51490
rect 17950 51438 18002 51490
rect 19182 51438 19234 51490
rect 23102 51438 23154 51490
rect 24110 51438 24162 51490
rect 25678 51438 25730 51490
rect 26910 51438 26962 51490
rect 1710 51326 1762 51378
rect 6190 51326 6242 51378
rect 9774 51326 9826 51378
rect 11790 51326 11842 51378
rect 15710 51326 15762 51378
rect 18062 51326 18114 51378
rect 19070 51326 19122 51378
rect 22430 51326 22482 51378
rect 22990 51326 23042 51378
rect 23774 51326 23826 51378
rect 24670 51326 24722 51378
rect 26238 51326 26290 51378
rect 37774 51326 37826 51378
rect 2494 51214 2546 51266
rect 6862 51214 6914 51266
rect 8990 51214 9042 51266
rect 14590 51214 14642 51266
rect 18622 51214 18674 51266
rect 27358 51214 27410 51266
rect 27806 51214 27858 51266
rect 27358 51102 27410 51154
rect 27806 51102 27858 51154
rect 36766 51102 36818 51154
rect 4478 50934 4530 50986
rect 4582 50934 4634 50986
rect 4686 50934 4738 50986
rect 35198 50934 35250 50986
rect 35302 50934 35354 50986
rect 35406 50934 35458 50986
rect 11454 50766 11506 50818
rect 12350 50766 12402 50818
rect 32958 50766 33010 50818
rect 11678 50654 11730 50706
rect 17614 50654 17666 50706
rect 17726 50654 17778 50706
rect 19742 50654 19794 50706
rect 33518 50654 33570 50706
rect 7422 50542 7474 50594
rect 8542 50542 8594 50594
rect 9438 50542 9490 50594
rect 10558 50542 10610 50594
rect 12126 50542 12178 50594
rect 12686 50542 12738 50594
rect 15822 50542 15874 50594
rect 20750 50542 20802 50594
rect 26574 50542 26626 50594
rect 33294 50542 33346 50594
rect 1710 50430 1762 50482
rect 2382 50430 2434 50482
rect 2718 50430 2770 50482
rect 3166 50430 3218 50482
rect 7758 50430 7810 50482
rect 8318 50430 8370 50482
rect 9550 50430 9602 50482
rect 9774 50430 9826 50482
rect 9998 50430 10050 50482
rect 12910 50430 12962 50482
rect 15150 50430 15202 50482
rect 15262 50430 15314 50482
rect 16382 50430 16434 50482
rect 20638 50430 20690 50482
rect 22990 50430 23042 50482
rect 27022 50430 27074 50482
rect 2046 50318 2098 50370
rect 7646 50318 7698 50370
rect 10334 50318 10386 50370
rect 11678 50318 11730 50370
rect 12798 50318 12850 50370
rect 19838 50150 19890 50202
rect 19942 50150 19994 50202
rect 20046 50150 20098 50202
rect 2494 49982 2546 50034
rect 10446 49982 10498 50034
rect 15598 49982 15650 50034
rect 23886 49982 23938 50034
rect 2046 49870 2098 49922
rect 9550 49870 9602 49922
rect 9662 49870 9714 49922
rect 11230 49870 11282 49922
rect 12686 49870 12738 49922
rect 15374 49870 15426 49922
rect 15934 49870 15986 49922
rect 19070 49870 19122 49922
rect 21086 49870 21138 49922
rect 22654 49870 22706 49922
rect 23326 49870 23378 49922
rect 23550 49870 23602 49922
rect 1710 49758 1762 49810
rect 5294 49758 5346 49810
rect 9886 49758 9938 49810
rect 10222 49758 10274 49810
rect 11566 49758 11618 49810
rect 11902 49758 11954 49810
rect 16270 49758 16322 49810
rect 17614 49758 17666 49810
rect 18398 49758 18450 49810
rect 21646 49758 21698 49810
rect 22094 49758 22146 49810
rect 23998 49758 24050 49810
rect 31166 49758 31218 49810
rect 34862 49758 34914 49810
rect 2942 49646 2994 49698
rect 5966 49646 6018 49698
rect 8206 49646 8258 49698
rect 11342 49646 11394 49698
rect 14814 49646 14866 49698
rect 18510 49646 18562 49698
rect 22206 49646 22258 49698
rect 28366 49646 28418 49698
rect 30494 49646 30546 49698
rect 35646 49646 35698 49698
rect 37774 49646 37826 49698
rect 10558 49534 10610 49586
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 9886 49086 9938 49138
rect 18062 49086 18114 49138
rect 22766 49086 22818 49138
rect 24222 49086 24274 49138
rect 29150 49086 29202 49138
rect 32398 49086 32450 49138
rect 33406 49086 33458 49138
rect 35646 49086 35698 49138
rect 7198 48974 7250 49026
rect 7534 48974 7586 49026
rect 8206 48974 8258 49026
rect 8654 48974 8706 49026
rect 15486 48974 15538 49026
rect 15710 48974 15762 49026
rect 15934 48974 15986 49026
rect 17838 48974 17890 49026
rect 19182 48974 19234 49026
rect 20414 48974 20466 49026
rect 22318 48974 22370 49026
rect 23102 48974 23154 49026
rect 23662 48974 23714 49026
rect 27022 48974 27074 49026
rect 31950 48974 32002 49026
rect 33294 48974 33346 49026
rect 35086 48974 35138 49026
rect 35422 48974 35474 49026
rect 35982 48974 36034 49026
rect 1710 48862 1762 48914
rect 2046 48862 2098 48914
rect 6638 48862 6690 48914
rect 8878 48862 8930 48914
rect 19966 48862 20018 48914
rect 22766 48862 22818 48914
rect 26350 48862 26402 48914
rect 31278 48862 31330 48914
rect 34414 48862 34466 48914
rect 2494 48750 2546 48802
rect 6750 48750 6802 48802
rect 6974 48750 7026 48802
rect 7310 48750 7362 48802
rect 8430 48750 8482 48802
rect 16270 48750 16322 48802
rect 21758 48750 21810 48802
rect 32958 48750 33010 48802
rect 33518 48750 33570 48802
rect 33742 48750 33794 48802
rect 34638 48750 34690 48802
rect 34750 48750 34802 48802
rect 34862 48750 34914 48802
rect 35646 48750 35698 48802
rect 35870 48750 35922 48802
rect 19838 48582 19890 48634
rect 19942 48582 19994 48634
rect 20046 48582 20098 48634
rect 6638 48414 6690 48466
rect 6862 48414 6914 48466
rect 7646 48414 7698 48466
rect 11118 48414 11170 48466
rect 18398 48414 18450 48466
rect 18622 48414 18674 48466
rect 20862 48414 20914 48466
rect 21422 48414 21474 48466
rect 26126 48414 26178 48466
rect 31278 48414 31330 48466
rect 32510 48414 32562 48466
rect 2046 48302 2098 48354
rect 6974 48302 7026 48354
rect 7310 48302 7362 48354
rect 18174 48302 18226 48354
rect 21198 48302 21250 48354
rect 22206 48302 22258 48354
rect 23998 48302 24050 48354
rect 24110 48302 24162 48354
rect 25566 48302 25618 48354
rect 26798 48302 26850 48354
rect 27134 48302 27186 48354
rect 27470 48302 27522 48354
rect 32174 48302 32226 48354
rect 32286 48302 32338 48354
rect 33630 48302 33682 48354
rect 1710 48190 1762 48242
rect 11342 48190 11394 48242
rect 11566 48190 11618 48242
rect 11902 48190 11954 48242
rect 18734 48190 18786 48242
rect 20302 48190 20354 48242
rect 21534 48190 21586 48242
rect 21646 48190 21698 48242
rect 21870 48190 21922 48242
rect 22318 48190 22370 48242
rect 22542 48190 22594 48242
rect 22766 48190 22818 48242
rect 24222 48190 24274 48242
rect 24670 48190 24722 48242
rect 25342 48190 25394 48242
rect 26462 48190 26514 48242
rect 31838 48190 31890 48242
rect 33294 48190 33346 48242
rect 38222 48190 38274 48242
rect 2494 48078 2546 48130
rect 18510 48078 18562 48130
rect 28030 48078 28082 48130
rect 33182 48078 33234 48130
rect 34862 48078 34914 48130
rect 36878 48078 36930 48130
rect 11342 47966 11394 48018
rect 20526 47966 20578 48018
rect 23214 47966 23266 48018
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 20750 47630 20802 47682
rect 33742 47630 33794 47682
rect 25006 47518 25058 47570
rect 25342 47518 25394 47570
rect 26574 47518 26626 47570
rect 27246 47518 27298 47570
rect 29934 47518 29986 47570
rect 31838 47518 31890 47570
rect 7982 47406 8034 47458
rect 18286 47406 18338 47458
rect 30158 47406 30210 47458
rect 32622 47406 32674 47458
rect 34078 47406 34130 47458
rect 34302 47406 34354 47458
rect 8094 47294 8146 47346
rect 17614 47294 17666 47346
rect 17950 47294 18002 47346
rect 20414 47294 20466 47346
rect 30494 47294 30546 47346
rect 30830 47294 30882 47346
rect 32958 47294 33010 47346
rect 8318 47182 8370 47234
rect 9214 47182 9266 47234
rect 18174 47182 18226 47234
rect 20638 47182 20690 47234
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 10446 46846 10498 46898
rect 11342 46846 11394 46898
rect 15486 46846 15538 46898
rect 21870 46846 21922 46898
rect 32062 46846 32114 46898
rect 8430 46734 8482 46786
rect 8766 46734 8818 46786
rect 9438 46734 9490 46786
rect 9662 46734 9714 46786
rect 10782 46734 10834 46786
rect 30830 46734 30882 46786
rect 31390 46734 31442 46786
rect 31726 46734 31778 46786
rect 31950 46734 32002 46786
rect 32286 46734 32338 46786
rect 33070 46734 33122 46786
rect 36094 46734 36146 46786
rect 8990 46622 9042 46674
rect 9774 46622 9826 46674
rect 10110 46622 10162 46674
rect 10558 46622 10610 46674
rect 17502 46622 17554 46674
rect 17950 46622 18002 46674
rect 19182 46622 19234 46674
rect 21758 46622 21810 46674
rect 21982 46622 22034 46674
rect 22094 46622 22146 46674
rect 28030 46622 28082 46674
rect 31614 46622 31666 46674
rect 32510 46622 32562 46674
rect 33294 46622 33346 46674
rect 33742 46622 33794 46674
rect 35310 46622 35362 46674
rect 8542 46510 8594 46562
rect 15374 46510 15426 46562
rect 15822 46510 15874 46562
rect 19294 46510 19346 46562
rect 25230 46510 25282 46562
rect 27358 46510 27410 46562
rect 34638 46510 34690 46562
rect 38222 46510 38274 46562
rect 15934 46398 15986 46450
rect 19518 46398 19570 46450
rect 22430 46398 22482 46450
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 21646 46062 21698 46114
rect 23998 46062 24050 46114
rect 7310 45950 7362 46002
rect 9438 45950 9490 46002
rect 10782 45950 10834 46002
rect 12910 45950 12962 46002
rect 14926 45950 14978 46002
rect 15822 45950 15874 46002
rect 16942 45950 16994 46002
rect 25678 45950 25730 46002
rect 30382 45950 30434 46002
rect 34750 45950 34802 46002
rect 6526 45838 6578 45890
rect 10110 45838 10162 45890
rect 15374 45838 15426 45890
rect 15934 45838 15986 45890
rect 22094 45838 22146 45890
rect 22430 45838 22482 45890
rect 25230 45838 25282 45890
rect 29598 45838 29650 45890
rect 30046 45838 30098 45890
rect 31390 45838 31442 45890
rect 36430 45838 36482 45890
rect 14254 45726 14306 45778
rect 14590 45726 14642 45778
rect 16606 45726 16658 45778
rect 21534 45726 21586 45778
rect 23550 45726 23602 45778
rect 24110 45726 24162 45778
rect 24558 45726 24610 45778
rect 24894 45726 24946 45778
rect 29262 45726 29314 45778
rect 32286 45726 32338 45778
rect 33182 45726 33234 45778
rect 13918 45614 13970 45666
rect 14814 45614 14866 45666
rect 17054 45614 17106 45666
rect 32398 45614 32450 45666
rect 33294 45614 33346 45666
rect 33406 45614 33458 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 8990 45278 9042 45330
rect 9886 45278 9938 45330
rect 10558 45278 10610 45330
rect 10782 45278 10834 45330
rect 14814 45278 14866 45330
rect 17838 45278 17890 45330
rect 18622 45278 18674 45330
rect 25566 45278 25618 45330
rect 26014 45278 26066 45330
rect 26126 45278 26178 45330
rect 33070 45278 33122 45330
rect 2046 45166 2098 45218
rect 6862 45166 6914 45218
rect 10222 45166 10274 45218
rect 15038 45166 15090 45218
rect 18062 45166 18114 45218
rect 18398 45166 18450 45218
rect 18846 45166 18898 45218
rect 23214 45166 23266 45218
rect 30830 45166 30882 45218
rect 32174 45166 32226 45218
rect 34638 45166 34690 45218
rect 1710 45054 1762 45106
rect 6974 45054 7026 45106
rect 10894 45054 10946 45106
rect 14030 45054 14082 45106
rect 14478 45054 14530 45106
rect 16046 45054 16098 45106
rect 16606 45054 16658 45106
rect 17502 45054 17554 45106
rect 19854 45054 19906 45106
rect 19966 45054 20018 45106
rect 22878 45054 22930 45106
rect 29598 45054 29650 45106
rect 30158 45054 30210 45106
rect 32398 45054 32450 45106
rect 33294 45054 33346 45106
rect 34078 45054 34130 45106
rect 34302 45054 34354 45106
rect 35310 45054 35362 45106
rect 2494 44942 2546 44994
rect 14254 44942 14306 44994
rect 18734 44942 18786 44994
rect 31950 44942 32002 44994
rect 36094 44942 36146 44994
rect 38222 44942 38274 44994
rect 6862 44830 6914 44882
rect 15598 44830 15650 44882
rect 16718 44830 16770 44882
rect 18174 44830 18226 44882
rect 20190 44830 20242 44882
rect 20302 44830 20354 44882
rect 26238 44830 26290 44882
rect 34750 44830 34802 44882
rect 34862 44830 34914 44882
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 6750 44494 6802 44546
rect 19966 44494 20018 44546
rect 20750 44494 20802 44546
rect 8318 44382 8370 44434
rect 10782 44382 10834 44434
rect 12910 44382 12962 44434
rect 21870 44382 21922 44434
rect 24894 44382 24946 44434
rect 35086 44382 35138 44434
rect 6638 44270 6690 44322
rect 8542 44270 8594 44322
rect 8766 44270 8818 44322
rect 10110 44270 10162 44322
rect 13582 44270 13634 44322
rect 15710 44270 15762 44322
rect 17726 44270 17778 44322
rect 21646 44270 21698 44322
rect 23662 44270 23714 44322
rect 26462 44270 26514 44322
rect 30606 44270 30658 44322
rect 30942 44270 30994 44322
rect 1710 44158 1762 44210
rect 6750 44158 6802 44210
rect 7534 44158 7586 44210
rect 8206 44158 8258 44210
rect 13694 44158 13746 44210
rect 16158 44158 16210 44210
rect 17950 44158 18002 44210
rect 18286 44158 18338 44210
rect 18958 44158 19010 44210
rect 19182 44158 19234 44210
rect 19406 44158 19458 44210
rect 19630 44158 19682 44210
rect 20414 44158 20466 44210
rect 22318 44158 22370 44210
rect 23774 44158 23826 44210
rect 24782 44158 24834 44210
rect 2046 44046 2098 44098
rect 2494 44046 2546 44098
rect 7646 44046 7698 44098
rect 7870 44046 7922 44098
rect 17278 44046 17330 44098
rect 20638 44046 20690 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 8206 43710 8258 43762
rect 9886 43710 9938 43762
rect 12910 43710 12962 43762
rect 26462 43710 26514 43762
rect 32174 43710 32226 43762
rect 34414 43710 34466 43762
rect 5966 43598 6018 43650
rect 10110 43598 10162 43650
rect 10446 43598 10498 43650
rect 12574 43598 12626 43650
rect 21422 43598 21474 43650
rect 24334 43598 24386 43650
rect 27134 43598 27186 43650
rect 27470 43598 27522 43650
rect 27806 43598 27858 43650
rect 28590 43598 28642 43650
rect 30718 43598 30770 43650
rect 30830 43598 30882 43650
rect 31166 43598 31218 43650
rect 31726 43598 31778 43650
rect 32286 43598 32338 43650
rect 33518 43598 33570 43650
rect 5294 43486 5346 43538
rect 13918 43486 13970 43538
rect 16158 43486 16210 43538
rect 16382 43486 16434 43538
rect 18286 43486 18338 43538
rect 19854 43486 19906 43538
rect 21198 43486 21250 43538
rect 21534 43486 21586 43538
rect 21870 43486 21922 43538
rect 22206 43486 22258 43538
rect 23214 43486 23266 43538
rect 23550 43486 23602 43538
rect 23662 43486 23714 43538
rect 23886 43486 23938 43538
rect 25566 43486 25618 43538
rect 26126 43486 26178 43538
rect 26798 43486 26850 43538
rect 28030 43486 28082 43538
rect 28366 43486 28418 43538
rect 28702 43486 28754 43538
rect 29598 43486 29650 43538
rect 29822 43486 29874 43538
rect 30046 43486 30098 43538
rect 30270 43486 30322 43538
rect 32398 43486 32450 43538
rect 33406 43486 33458 43538
rect 33966 43486 34018 43538
rect 35310 43486 35362 43538
rect 14030 43374 14082 43426
rect 15934 43374 15986 43426
rect 18622 43374 18674 43426
rect 19742 43374 19794 43426
rect 33742 43374 33794 43426
rect 36094 43374 36146 43426
rect 38222 43374 38274 43426
rect 18510 43262 18562 43314
rect 30158 43262 30210 43314
rect 30606 43262 30658 43314
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 14142 42926 14194 42978
rect 20190 42926 20242 42978
rect 20414 42926 20466 42978
rect 26238 42926 26290 42978
rect 9886 42814 9938 42866
rect 18398 42814 18450 42866
rect 26014 42814 26066 42866
rect 31726 42814 31778 42866
rect 32622 42814 32674 42866
rect 7086 42702 7138 42754
rect 10334 42702 10386 42754
rect 10558 42702 10610 42754
rect 10894 42702 10946 42754
rect 15150 42702 15202 42754
rect 16046 42702 16098 42754
rect 17726 42702 17778 42754
rect 19966 42702 20018 42754
rect 20638 42702 20690 42754
rect 25678 42702 25730 42754
rect 28366 42702 28418 42754
rect 28702 42702 28754 42754
rect 29486 42702 29538 42754
rect 29710 42702 29762 42754
rect 30606 42702 30658 42754
rect 33070 42702 33122 42754
rect 33294 42702 33346 42754
rect 33406 42702 33458 42754
rect 36430 42702 36482 42754
rect 7758 42590 7810 42642
rect 14702 42590 14754 42642
rect 15374 42590 15426 42642
rect 16606 42590 16658 42642
rect 17614 42590 17666 42642
rect 20750 42590 20802 42642
rect 21310 42590 21362 42642
rect 30046 42590 30098 42642
rect 31166 42590 31218 42642
rect 31278 42590 31330 42642
rect 31614 42590 31666 42642
rect 32062 42590 32114 42642
rect 32846 42590 32898 42642
rect 10558 42478 10610 42530
rect 11230 42478 11282 42530
rect 21422 42478 21474 42530
rect 21646 42478 21698 42530
rect 26798 42478 26850 42530
rect 28478 42478 28530 42530
rect 30942 42478 30994 42530
rect 32286 42478 32338 42530
rect 32510 42478 32562 42530
rect 33182 42478 33234 42530
rect 35422 42478 35474 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 7982 42142 8034 42194
rect 8206 42142 8258 42194
rect 16046 42142 16098 42194
rect 20414 42142 20466 42194
rect 28142 42142 28194 42194
rect 33294 42142 33346 42194
rect 34414 42142 34466 42194
rect 8318 42030 8370 42082
rect 22766 42030 22818 42082
rect 22878 42030 22930 42082
rect 30270 42030 30322 42082
rect 30606 42030 30658 42082
rect 31278 42030 31330 42082
rect 14814 41918 14866 41970
rect 16606 41918 16658 41970
rect 18286 41918 18338 41970
rect 18622 41918 18674 41970
rect 18734 41918 18786 41970
rect 18958 41918 19010 41970
rect 19630 41918 19682 41970
rect 19854 41918 19906 41970
rect 19966 41918 20018 41970
rect 22542 41918 22594 41970
rect 25230 41918 25282 41970
rect 27806 41918 27858 41970
rect 28254 41918 28306 41970
rect 28366 41918 28418 41970
rect 29262 41918 29314 41970
rect 29486 41918 29538 41970
rect 31054 41918 31106 41970
rect 31502 41918 31554 41970
rect 31726 41918 31778 41970
rect 31950 41918 32002 41970
rect 32286 41918 32338 41970
rect 32958 41918 33010 41970
rect 33294 41918 33346 41970
rect 33630 41918 33682 41970
rect 34190 41918 34242 41970
rect 34526 41918 34578 41970
rect 34638 41918 34690 41970
rect 34750 41918 34802 41970
rect 35422 41918 35474 41970
rect 17502 41806 17554 41858
rect 25678 41806 25730 41858
rect 29710 41806 29762 41858
rect 36094 41806 36146 41858
rect 38222 41806 38274 41858
rect 14926 41694 14978 41746
rect 25454 41694 25506 41746
rect 25902 41694 25954 41746
rect 26350 41694 26402 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 22542 41358 22594 41410
rect 29374 41358 29426 41410
rect 34974 41358 35026 41410
rect 20078 41246 20130 41298
rect 20638 41246 20690 41298
rect 29598 41246 29650 41298
rect 30606 41246 30658 41298
rect 31390 41246 31442 41298
rect 1822 41134 1874 41186
rect 10894 41134 10946 41186
rect 11230 41134 11282 41186
rect 11566 41134 11618 41186
rect 11902 41134 11954 41186
rect 19182 41134 19234 41186
rect 19854 41134 19906 41186
rect 21646 41134 21698 41186
rect 22094 41134 22146 41186
rect 22990 41134 23042 41186
rect 24110 41134 24162 41186
rect 26238 41134 26290 41186
rect 28702 41134 28754 41186
rect 31054 41134 31106 41186
rect 31278 41134 31330 41186
rect 31726 41134 31778 41186
rect 32622 41134 32674 41186
rect 33182 41134 33234 41186
rect 36318 41134 36370 41186
rect 2494 41022 2546 41074
rect 14142 41022 14194 41074
rect 19630 41022 19682 41074
rect 20190 41022 20242 41074
rect 21758 41022 21810 41074
rect 21870 41022 21922 41074
rect 24782 41022 24834 41074
rect 26798 41022 26850 41074
rect 28366 41022 28418 41074
rect 29262 41022 29314 41074
rect 31838 41022 31890 41074
rect 32734 41022 32786 41074
rect 33518 41022 33570 41074
rect 2046 40910 2098 40962
rect 11342 40910 11394 40962
rect 23102 40910 23154 40962
rect 23214 40910 23266 40962
rect 23438 40910 23490 40962
rect 27806 40910 27858 40962
rect 28478 40910 28530 40962
rect 31502 40910 31554 40962
rect 32958 40910 33010 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 9774 40574 9826 40626
rect 10334 40574 10386 40626
rect 14254 40574 14306 40626
rect 18846 40574 18898 40626
rect 19854 40574 19906 40626
rect 20190 40574 20242 40626
rect 22430 40574 22482 40626
rect 30158 40574 30210 40626
rect 30382 40574 30434 40626
rect 30718 40574 30770 40626
rect 31950 40574 32002 40626
rect 32398 40574 32450 40626
rect 2046 40462 2098 40514
rect 9662 40462 9714 40514
rect 20078 40462 20130 40514
rect 20414 40462 20466 40514
rect 23326 40462 23378 40514
rect 32510 40462 32562 40514
rect 33854 40462 33906 40514
rect 1710 40350 1762 40402
rect 2494 40350 2546 40402
rect 13246 40350 13298 40402
rect 13470 40350 13522 40402
rect 19518 40350 19570 40402
rect 21310 40350 21362 40402
rect 24334 40350 24386 40402
rect 30046 40350 30098 40402
rect 30606 40350 30658 40402
rect 30942 40350 30994 40402
rect 31390 40350 31442 40402
rect 32062 40350 32114 40402
rect 33182 40350 33234 40402
rect 13694 40238 13746 40290
rect 20974 40238 21026 40290
rect 21534 40238 21586 40290
rect 21758 40238 21810 40290
rect 23662 40238 23714 40290
rect 23998 40238 24050 40290
rect 35982 40238 36034 40290
rect 9774 40126 9826 40178
rect 20638 40126 20690 40178
rect 21982 40126 22034 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 18846 39790 18898 39842
rect 12910 39678 12962 39730
rect 19070 39678 19122 39730
rect 19630 39678 19682 39730
rect 20190 39678 20242 39730
rect 25566 39678 25618 39730
rect 29598 39678 29650 39730
rect 33182 39678 33234 39730
rect 8542 39566 8594 39618
rect 8766 39566 8818 39618
rect 9214 39566 9266 39618
rect 9774 39566 9826 39618
rect 10110 39566 10162 39618
rect 16382 39566 16434 39618
rect 18510 39566 18562 39618
rect 19518 39566 19570 39618
rect 19966 39566 20018 39618
rect 20302 39566 20354 39618
rect 22766 39566 22818 39618
rect 22990 39566 23042 39618
rect 24782 39566 24834 39618
rect 30830 39566 30882 39618
rect 1710 39454 1762 39506
rect 8206 39454 8258 39506
rect 9326 39454 9378 39506
rect 10782 39454 10834 39506
rect 14926 39454 14978 39506
rect 17390 39454 17442 39506
rect 19294 39454 19346 39506
rect 20638 39454 20690 39506
rect 25790 39454 25842 39506
rect 2046 39342 2098 39394
rect 2494 39342 2546 39394
rect 8430 39342 8482 39394
rect 9438 39342 9490 39394
rect 15038 39342 15090 39394
rect 19742 39342 19794 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 8206 39006 8258 39058
rect 9662 39006 9714 39058
rect 10334 39006 10386 39058
rect 10670 39006 10722 39058
rect 11118 39006 11170 39058
rect 18398 39006 18450 39058
rect 26238 39006 26290 39058
rect 26910 39006 26962 39058
rect 7534 38894 7586 38946
rect 7646 38894 7698 38946
rect 8094 38894 8146 38946
rect 8766 38894 8818 38946
rect 9550 38894 9602 38946
rect 9886 38894 9938 38946
rect 11342 38894 11394 38946
rect 11454 38894 11506 38946
rect 12574 38894 12626 38946
rect 12686 38894 12738 38946
rect 13022 38894 13074 38946
rect 14030 38894 14082 38946
rect 15710 38894 15762 38946
rect 17838 38894 17890 38946
rect 19070 38894 19122 38946
rect 19182 38894 19234 38946
rect 23326 38894 23378 38946
rect 25342 38894 25394 38946
rect 26126 38894 26178 38946
rect 34190 38894 34242 38946
rect 7870 38782 7922 38834
rect 8430 38782 8482 38834
rect 8654 38782 8706 38834
rect 8990 38782 9042 38834
rect 15150 38782 15202 38834
rect 17390 38782 17442 38834
rect 18286 38782 18338 38834
rect 18846 38782 18898 38834
rect 19630 38782 19682 38834
rect 20414 38782 20466 38834
rect 20638 38782 20690 38834
rect 21646 38782 21698 38834
rect 23662 38782 23714 38834
rect 24334 38782 24386 38834
rect 25230 38782 25282 38834
rect 26462 38782 26514 38834
rect 33406 38782 33458 38834
rect 13694 38670 13746 38722
rect 21534 38670 21586 38722
rect 22094 38670 22146 38722
rect 22766 38670 22818 38722
rect 23550 38670 23602 38722
rect 36318 38670 36370 38722
rect 13134 38558 13186 38610
rect 22542 38558 22594 38610
rect 22878 38558 22930 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 23774 38222 23826 38274
rect 24446 38222 24498 38274
rect 24782 38222 24834 38274
rect 25678 38222 25730 38274
rect 26014 38222 26066 38274
rect 26910 38222 26962 38274
rect 27582 38222 27634 38274
rect 34974 38222 35026 38274
rect 6974 38110 7026 38162
rect 9102 38110 9154 38162
rect 14926 38110 14978 38162
rect 22094 38110 22146 38162
rect 24222 38110 24274 38162
rect 25454 38110 25506 38162
rect 26574 38110 26626 38162
rect 28030 38110 28082 38162
rect 29486 38110 29538 38162
rect 31614 38110 31666 38162
rect 9886 37998 9938 38050
rect 14030 37998 14082 38050
rect 15038 37998 15090 38050
rect 20078 37998 20130 38050
rect 21646 37998 21698 38050
rect 22654 37998 22706 38050
rect 22878 37998 22930 38050
rect 23550 37998 23602 38050
rect 26238 37998 26290 38050
rect 27246 37998 27298 38050
rect 32398 37998 32450 38050
rect 36318 37998 36370 38050
rect 14702 37886 14754 37938
rect 16942 37886 16994 37938
rect 21310 37886 21362 37938
rect 26686 37886 26738 37938
rect 10334 37774 10386 37826
rect 21422 37774 21474 37826
rect 27470 37774 27522 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 16270 37438 16322 37490
rect 28478 37438 28530 37490
rect 19742 37326 19794 37378
rect 19854 37326 19906 37378
rect 25342 37326 25394 37378
rect 26462 37326 26514 37378
rect 28030 37326 28082 37378
rect 25454 37214 25506 37266
rect 25902 37214 25954 37266
rect 26686 37214 26738 37266
rect 27134 37214 27186 37266
rect 27358 37214 27410 37266
rect 16158 37102 16210 37154
rect 28926 37102 28978 37154
rect 19854 36990 19906 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 8766 36542 8818 36594
rect 10894 36542 10946 36594
rect 17950 36542 18002 36594
rect 24670 36542 24722 36594
rect 8094 36430 8146 36482
rect 16382 36430 16434 36482
rect 18622 36430 18674 36482
rect 27582 36430 27634 36482
rect 16046 36318 16098 36370
rect 17726 36318 17778 36370
rect 18286 36318 18338 36370
rect 26798 36318 26850 36370
rect 38222 36318 38274 36370
rect 11342 36206 11394 36258
rect 14590 36206 14642 36258
rect 28030 36206 28082 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 22542 35870 22594 35922
rect 25790 35870 25842 35922
rect 14926 35758 14978 35810
rect 15262 35758 15314 35810
rect 22654 35758 22706 35810
rect 27694 35758 27746 35810
rect 11566 35646 11618 35698
rect 17726 35646 17778 35698
rect 21870 35646 21922 35698
rect 25678 35646 25730 35698
rect 26910 35646 26962 35698
rect 12238 35534 12290 35586
rect 14366 35534 14418 35586
rect 15822 35534 15874 35586
rect 17614 35534 17666 35586
rect 22094 35534 22146 35586
rect 29822 35534 29874 35586
rect 17390 35422 17442 35474
rect 22206 35422 22258 35474
rect 25454 35422 25506 35474
rect 25790 35422 25842 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 13470 35086 13522 35138
rect 15150 34974 15202 35026
rect 19182 34974 19234 35026
rect 22654 34974 22706 35026
rect 23102 34974 23154 35026
rect 14366 34862 14418 34914
rect 14814 34862 14866 34914
rect 15262 34862 15314 34914
rect 15598 34862 15650 34914
rect 16382 34862 16434 34914
rect 21758 34862 21810 34914
rect 22206 34862 22258 34914
rect 13582 34750 13634 34802
rect 14254 34750 14306 34802
rect 15038 34750 15090 34802
rect 17054 34750 17106 34802
rect 14142 34638 14194 34690
rect 19630 34638 19682 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 15150 34302 15202 34354
rect 17502 34302 17554 34354
rect 21086 34302 21138 34354
rect 22766 34302 22818 34354
rect 24670 34302 24722 34354
rect 16270 34190 16322 34242
rect 16382 34190 16434 34242
rect 20302 34190 20354 34242
rect 22318 34190 22370 34242
rect 11790 34078 11842 34130
rect 16046 34078 16098 34130
rect 17390 34078 17442 34130
rect 17614 34078 17666 34130
rect 20078 34078 20130 34130
rect 20526 34078 20578 34130
rect 20638 34078 20690 34130
rect 21646 34078 21698 34130
rect 21982 34078 22034 34130
rect 24446 34078 24498 34130
rect 25342 34078 25394 34130
rect 25566 34078 25618 34130
rect 12574 33966 12626 34018
rect 14702 33966 14754 34018
rect 16606 33966 16658 34018
rect 21422 33966 21474 34018
rect 26238 33966 26290 34018
rect 15598 33854 15650 33906
rect 17838 33854 17890 33906
rect 19742 33854 19794 33906
rect 21982 33854 22034 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 13918 33518 13970 33570
rect 14366 33518 14418 33570
rect 17166 33518 17218 33570
rect 18734 33518 18786 33570
rect 19070 33518 19122 33570
rect 21422 33518 21474 33570
rect 21646 33518 21698 33570
rect 26014 33518 26066 33570
rect 13694 33406 13746 33458
rect 14030 33406 14082 33458
rect 17390 33406 17442 33458
rect 22318 33406 22370 33458
rect 23998 33406 24050 33458
rect 24894 33406 24946 33458
rect 26798 33406 26850 33458
rect 14254 33294 14306 33346
rect 14814 33294 14866 33346
rect 15150 33294 15202 33346
rect 15374 33294 15426 33346
rect 16830 33294 16882 33346
rect 18958 33294 19010 33346
rect 19966 33294 20018 33346
rect 20190 33294 20242 33346
rect 20302 33294 20354 33346
rect 20526 33294 20578 33346
rect 21758 33294 21810 33346
rect 26350 33294 26402 33346
rect 14926 33182 14978 33234
rect 18622 33182 18674 33234
rect 21310 33182 21362 33234
rect 1710 33070 1762 33122
rect 26126 33070 26178 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 24222 32734 24274 32786
rect 21086 32622 21138 32674
rect 23550 32622 23602 32674
rect 23774 32622 23826 32674
rect 27470 32622 27522 32674
rect 14030 32510 14082 32562
rect 14702 32510 14754 32562
rect 14926 32510 14978 32562
rect 21870 32510 21922 32562
rect 23214 32510 23266 32562
rect 24334 32510 24386 32562
rect 28142 32510 28194 32562
rect 14366 32398 14418 32450
rect 18622 32398 18674 32450
rect 18958 32398 19010 32450
rect 23326 32398 23378 32450
rect 25342 32398 25394 32450
rect 14030 32286 14082 32338
rect 15262 32286 15314 32338
rect 24222 32286 24274 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 14702 31950 14754 32002
rect 23438 31838 23490 31890
rect 14478 31726 14530 31778
rect 14926 31726 14978 31778
rect 15486 31726 15538 31778
rect 22542 31726 22594 31778
rect 22766 31726 22818 31778
rect 23214 31726 23266 31778
rect 26350 31726 26402 31778
rect 14366 31614 14418 31666
rect 25566 31614 25618 31666
rect 22654 31502 22706 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 20750 31166 20802 31218
rect 22878 31166 22930 31218
rect 25454 31166 25506 31218
rect 26126 31166 26178 31218
rect 12126 31054 12178 31106
rect 18174 31054 18226 31106
rect 21870 31054 21922 31106
rect 38222 31054 38274 31106
rect 11454 30942 11506 30994
rect 14702 30942 14754 30994
rect 17502 30942 17554 30994
rect 23214 30942 23266 30994
rect 23998 30942 24050 30994
rect 24670 30942 24722 30994
rect 25230 30942 25282 30994
rect 14254 30830 14306 30882
rect 20302 30830 20354 30882
rect 24222 30830 24274 30882
rect 25566 30830 25618 30882
rect 21982 30718 22034 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 20862 30270 20914 30322
rect 22094 30270 22146 30322
rect 24222 30270 24274 30322
rect 21310 30158 21362 30210
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 38222 23214 38274 23266
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 2942 3278 2994 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 3360 99200 3472 100000
rect 3388 95956 3444 99200
rect 4476 96460 4740 96470
rect 4532 96404 4580 96460
rect 4636 96404 4684 96460
rect 4476 96394 4740 96404
rect 35196 96460 35460 96470
rect 35252 96404 35300 96460
rect 35356 96404 35404 96460
rect 35196 96394 35460 96404
rect 3612 95956 3668 95966
rect 3388 95954 3668 95956
rect 3388 95902 3614 95954
rect 3666 95902 3668 95954
rect 3388 95900 3668 95902
rect 3612 95890 3668 95900
rect 19836 95676 20100 95686
rect 19892 95620 19940 95676
rect 19996 95620 20044 95676
rect 19836 95610 20100 95620
rect 4476 94892 4740 94902
rect 4532 94836 4580 94892
rect 4636 94836 4684 94892
rect 4476 94826 4740 94836
rect 35196 94892 35460 94902
rect 35252 94836 35300 94892
rect 35356 94836 35404 94892
rect 35196 94826 35460 94836
rect 19836 94108 20100 94118
rect 19892 94052 19940 94108
rect 19996 94052 20044 94108
rect 19836 94042 20100 94052
rect 4476 93324 4740 93334
rect 4532 93268 4580 93324
rect 4636 93268 4684 93324
rect 4476 93258 4740 93268
rect 35196 93324 35460 93334
rect 35252 93268 35300 93324
rect 35356 93268 35404 93324
rect 35196 93258 35460 93268
rect 19836 92540 20100 92550
rect 19892 92484 19940 92540
rect 19996 92484 20044 92540
rect 19836 92474 20100 92484
rect 4476 91756 4740 91766
rect 4532 91700 4580 91756
rect 4636 91700 4684 91756
rect 4476 91690 4740 91700
rect 35196 91756 35460 91766
rect 35252 91700 35300 91756
rect 35356 91700 35404 91756
rect 35196 91690 35460 91700
rect 19836 90972 20100 90982
rect 19892 90916 19940 90972
rect 19996 90916 20044 90972
rect 19836 90906 20100 90916
rect 4476 90188 4740 90198
rect 4532 90132 4580 90188
rect 4636 90132 4684 90188
rect 4476 90122 4740 90132
rect 35196 90188 35460 90198
rect 35252 90132 35300 90188
rect 35356 90132 35404 90188
rect 35196 90122 35460 90132
rect 19836 89404 20100 89414
rect 19892 89348 19940 89404
rect 19996 89348 20044 89404
rect 19836 89338 20100 89348
rect 4476 88620 4740 88630
rect 4532 88564 4580 88620
rect 4636 88564 4684 88620
rect 4476 88554 4740 88564
rect 35196 88620 35460 88630
rect 35252 88564 35300 88620
rect 35356 88564 35404 88620
rect 35196 88554 35460 88564
rect 19836 87836 20100 87846
rect 19892 87780 19940 87836
rect 19996 87780 20044 87836
rect 19836 87770 20100 87780
rect 4476 87052 4740 87062
rect 4532 86996 4580 87052
rect 4636 86996 4684 87052
rect 4476 86986 4740 86996
rect 35196 87052 35460 87062
rect 35252 86996 35300 87052
rect 35356 86996 35404 87052
rect 35196 86986 35460 86996
rect 19836 86268 20100 86278
rect 19892 86212 19940 86268
rect 19996 86212 20044 86268
rect 19836 86202 20100 86212
rect 4476 85484 4740 85494
rect 4532 85428 4580 85484
rect 4636 85428 4684 85484
rect 4476 85418 4740 85428
rect 35196 85484 35460 85494
rect 35252 85428 35300 85484
rect 35356 85428 35404 85484
rect 35196 85418 35460 85428
rect 19836 84700 20100 84710
rect 19892 84644 19940 84700
rect 19996 84644 20044 84700
rect 19836 84634 20100 84644
rect 4476 83916 4740 83926
rect 4532 83860 4580 83916
rect 4636 83860 4684 83916
rect 4476 83850 4740 83860
rect 35196 83916 35460 83926
rect 35252 83860 35300 83916
rect 35356 83860 35404 83916
rect 35196 83850 35460 83860
rect 19836 83132 20100 83142
rect 19892 83076 19940 83132
rect 19996 83076 20044 83132
rect 19836 83066 20100 83076
rect 4476 82348 4740 82358
rect 4532 82292 4580 82348
rect 4636 82292 4684 82348
rect 4476 82282 4740 82292
rect 35196 82348 35460 82358
rect 35252 82292 35300 82348
rect 35356 82292 35404 82348
rect 35196 82282 35460 82292
rect 19836 81564 20100 81574
rect 19892 81508 19940 81564
rect 19996 81508 20044 81564
rect 19836 81498 20100 81508
rect 4476 80780 4740 80790
rect 4532 80724 4580 80780
rect 4636 80724 4684 80780
rect 4476 80714 4740 80724
rect 35196 80780 35460 80790
rect 35252 80724 35300 80780
rect 35356 80724 35404 80780
rect 35196 80714 35460 80724
rect 19836 79996 20100 80006
rect 19892 79940 19940 79996
rect 19996 79940 20044 79996
rect 19836 79930 20100 79940
rect 4476 79212 4740 79222
rect 4532 79156 4580 79212
rect 4636 79156 4684 79212
rect 4476 79146 4740 79156
rect 35196 79212 35460 79222
rect 35252 79156 35300 79212
rect 35356 79156 35404 79212
rect 35196 79146 35460 79156
rect 19836 78428 20100 78438
rect 19892 78372 19940 78428
rect 19996 78372 20044 78428
rect 19836 78362 20100 78372
rect 4476 77644 4740 77654
rect 4532 77588 4580 77644
rect 4636 77588 4684 77644
rect 4476 77578 4740 77588
rect 35196 77644 35460 77654
rect 35252 77588 35300 77644
rect 35356 77588 35404 77644
rect 35196 77578 35460 77588
rect 19836 76860 20100 76870
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 19836 76794 20100 76804
rect 4476 76076 4740 76086
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4476 76010 4740 76020
rect 35196 76076 35460 76086
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35196 76010 35460 76020
rect 19836 75292 20100 75302
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 19836 75226 20100 75236
rect 4476 74508 4740 74518
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4476 74442 4740 74452
rect 35196 74508 35460 74518
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35196 74442 35460 74452
rect 19836 73724 20100 73734
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 19836 73658 20100 73668
rect 4476 72940 4740 72950
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4476 72874 4740 72884
rect 35196 72940 35460 72950
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35196 72874 35460 72884
rect 19836 72156 20100 72166
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 19836 72090 20100 72100
rect 4476 71372 4740 71382
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4476 71306 4740 71316
rect 35196 71372 35460 71382
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35196 71306 35460 71316
rect 19836 70588 20100 70598
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 19836 70522 20100 70532
rect 25340 70308 25396 70318
rect 25340 70306 25508 70308
rect 25340 70254 25342 70306
rect 25394 70254 25508 70306
rect 25340 70252 25508 70254
rect 25340 70242 25396 70252
rect 17948 70196 18004 70206
rect 17388 70194 18116 70196
rect 17388 70142 17950 70194
rect 18002 70142 18116 70194
rect 17388 70140 18116 70142
rect 4476 69804 4740 69814
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4476 69738 4740 69748
rect 13020 69412 13076 69422
rect 2044 68740 2100 68750
rect 2044 68646 2100 68684
rect 9660 68740 9716 68750
rect 9660 68646 9716 68684
rect 9772 68738 9828 68750
rect 9772 68686 9774 68738
rect 9826 68686 9828 68738
rect 1708 68626 1764 68638
rect 1708 68574 1710 68626
rect 1762 68574 1764 68626
rect 1708 68516 1764 68574
rect 8316 68628 8372 68638
rect 1708 67956 1764 68460
rect 2492 68516 2548 68526
rect 2492 68422 2548 68460
rect 4476 68236 4740 68246
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4476 68170 4740 68180
rect 1708 67890 1764 67900
rect 7644 67956 7700 67966
rect 7644 67862 7700 67900
rect 1708 67730 1764 67742
rect 1708 67678 1710 67730
rect 1762 67678 1764 67730
rect 1708 67284 1764 67678
rect 2044 67618 2100 67630
rect 2044 67566 2046 67618
rect 2098 67566 2100 67618
rect 2044 67396 2100 67566
rect 2044 67330 2100 67340
rect 2492 67618 2548 67630
rect 2492 67566 2494 67618
rect 2546 67566 2548 67618
rect 1708 67218 1764 67228
rect 2492 67284 2548 67566
rect 2492 67218 2548 67228
rect 8204 67396 8260 67406
rect 2044 67172 2100 67182
rect 2044 67078 2100 67116
rect 8204 67170 8260 67340
rect 8204 67118 8206 67170
rect 8258 67118 8260 67170
rect 8204 67106 8260 67118
rect 8316 67170 8372 68572
rect 9772 68628 9828 68686
rect 9772 68562 9828 68572
rect 10332 68626 10388 68638
rect 10332 68574 10334 68626
rect 10386 68574 10388 68626
rect 9772 68404 9828 68414
rect 9772 68310 9828 68348
rect 10332 68068 10388 68574
rect 11004 68514 11060 68526
rect 11004 68462 11006 68514
rect 11058 68462 11060 68514
rect 10332 68012 10948 68068
rect 8764 67956 8820 67966
rect 8316 67118 8318 67170
rect 8370 67118 8372 67170
rect 1708 67058 1764 67070
rect 1708 67006 1710 67058
rect 1762 67006 1764 67058
rect 1708 66612 1764 67006
rect 1708 66546 1764 66556
rect 2492 66946 2548 66958
rect 2492 66894 2494 66946
rect 2546 66894 2548 66946
rect 2492 66612 2548 66894
rect 4476 66668 4740 66678
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4476 66602 4740 66612
rect 2492 66546 2548 66556
rect 2156 65378 2212 65390
rect 2156 65326 2158 65378
rect 2210 65326 2212 65378
rect 1820 64706 1876 64718
rect 1820 64654 1822 64706
rect 1874 64654 1876 64706
rect 1820 64484 1876 64654
rect 2156 64596 2212 65326
rect 8316 65156 8372 67118
rect 8540 67172 8596 67182
rect 8540 67170 8708 67172
rect 8540 67118 8542 67170
rect 8594 67118 8708 67170
rect 8540 67116 8708 67118
rect 8540 67106 8596 67116
rect 8652 67060 8708 67116
rect 8764 67170 8820 67900
rect 10556 67842 10612 68012
rect 10780 67844 10836 67854
rect 10556 67790 10558 67842
rect 10610 67790 10612 67842
rect 10556 67778 10612 67790
rect 10668 67842 10836 67844
rect 10668 67790 10782 67842
rect 10834 67790 10836 67842
rect 10668 67788 10836 67790
rect 9772 67730 9828 67742
rect 9772 67678 9774 67730
rect 9826 67678 9828 67730
rect 9772 67282 9828 67678
rect 9772 67230 9774 67282
rect 9826 67230 9828 67282
rect 9772 67218 9828 67230
rect 10108 67732 10164 67742
rect 8764 67118 8766 67170
rect 8818 67118 8820 67170
rect 8764 67106 8820 67118
rect 8876 67170 8932 67182
rect 8876 67118 8878 67170
rect 8930 67118 8932 67170
rect 8652 66994 8708 67004
rect 4476 65100 4740 65110
rect 8316 65100 8820 65156
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4476 65034 4740 65044
rect 2380 64596 2436 64606
rect 2156 64540 2380 64596
rect 2380 64502 2436 64540
rect 2716 64596 2772 64606
rect 2716 64502 2772 64540
rect 8652 64596 8708 64606
rect 8652 64502 8708 64540
rect 8764 64596 8820 65100
rect 8876 64820 8932 67118
rect 9884 67172 9940 67182
rect 9100 67058 9156 67070
rect 9100 67006 9102 67058
rect 9154 67006 9156 67058
rect 9100 66836 9156 67006
rect 9436 67060 9492 67070
rect 9436 66966 9492 67004
rect 9772 67058 9828 67070
rect 9772 67006 9774 67058
rect 9826 67006 9828 67058
rect 9772 66836 9828 67006
rect 9100 66780 9828 66836
rect 9884 66274 9940 67116
rect 9884 66222 9886 66274
rect 9938 66222 9940 66274
rect 9884 66210 9940 66222
rect 10108 67170 10164 67676
rect 10668 67172 10724 67788
rect 10780 67778 10836 67788
rect 10108 67118 10110 67170
rect 10162 67118 10164 67170
rect 9660 66050 9716 66062
rect 9660 65998 9662 66050
rect 9714 65998 9716 66050
rect 9660 65940 9716 65998
rect 9996 66050 10052 66062
rect 9996 65998 9998 66050
rect 10050 65998 10052 66050
rect 9996 65940 10052 65998
rect 9660 65884 10052 65940
rect 9660 65828 9716 65884
rect 8876 64754 8932 64764
rect 9212 65772 9716 65828
rect 8764 64594 8932 64596
rect 8764 64542 8766 64594
rect 8818 64542 8932 64594
rect 8764 64540 8932 64542
rect 8764 64530 8820 64540
rect 1708 63922 1764 63934
rect 1708 63870 1710 63922
rect 1762 63870 1764 63922
rect 1708 63252 1764 63870
rect 1820 63924 1876 64428
rect 2044 64484 2100 64494
rect 3164 64484 3220 64494
rect 2044 64482 2212 64484
rect 2044 64430 2046 64482
rect 2098 64430 2212 64482
rect 2044 64428 2212 64430
rect 2044 64418 2100 64428
rect 1820 63858 1876 63868
rect 2044 64034 2100 64046
rect 2044 63982 2046 64034
rect 2098 63982 2100 64034
rect 2044 63812 2100 63982
rect 2044 63746 2100 63756
rect 2156 63364 2212 64428
rect 3164 64390 3220 64428
rect 2156 63298 2212 63308
rect 2492 63922 2548 63934
rect 2492 63870 2494 63922
rect 2546 63870 2548 63922
rect 1708 63186 1764 63196
rect 2492 63252 2548 63870
rect 8876 63588 8932 64540
rect 8988 64482 9044 64494
rect 8988 64430 8990 64482
rect 9042 64430 9044 64482
rect 8988 64036 9044 64430
rect 9212 64484 9268 65772
rect 9436 65604 9492 65614
rect 9324 64708 9380 64718
rect 9436 64708 9492 65548
rect 10108 65492 10164 67118
rect 10220 67116 10724 67172
rect 10220 66274 10276 67116
rect 10220 66222 10222 66274
rect 10274 66222 10276 66274
rect 10220 66210 10276 66222
rect 10892 67058 10948 68012
rect 11004 67954 11060 68462
rect 11004 67902 11006 67954
rect 11058 67902 11060 67954
rect 11004 67890 11060 67902
rect 11788 68404 11844 68414
rect 11788 67842 11844 68348
rect 11788 67790 11790 67842
rect 11842 67790 11844 67842
rect 11788 67778 11844 67790
rect 12124 67900 12516 67956
rect 12124 67842 12180 67900
rect 12124 67790 12126 67842
rect 12178 67790 12180 67842
rect 12124 67778 12180 67790
rect 12460 67844 12516 67900
rect 12572 67844 12628 67854
rect 12460 67842 12628 67844
rect 12460 67790 12574 67842
rect 12626 67790 12628 67842
rect 12460 67788 12628 67790
rect 12572 67778 12628 67788
rect 10892 67006 10894 67058
rect 10946 67006 10948 67058
rect 10892 65604 10948 67006
rect 11228 67730 11284 67742
rect 11228 67678 11230 67730
rect 11282 67678 11284 67730
rect 11228 66500 11284 67678
rect 11452 67732 11508 67742
rect 11452 67638 11508 67676
rect 12348 67732 12404 67742
rect 12348 67638 12404 67676
rect 12908 67732 12964 67742
rect 12908 67638 12964 67676
rect 11900 67618 11956 67630
rect 11900 67566 11902 67618
rect 11954 67566 11956 67618
rect 11900 67284 11956 67566
rect 11676 67228 11956 67284
rect 12796 67620 12852 67630
rect 11676 67170 11732 67228
rect 11676 67118 11678 67170
rect 11730 67118 11732 67170
rect 11676 67106 11732 67118
rect 11228 66434 11284 66444
rect 12572 66500 12628 66510
rect 12572 66274 12628 66444
rect 12572 66222 12574 66274
rect 12626 66222 12628 66274
rect 12572 66210 12628 66222
rect 12348 66052 12404 66062
rect 12796 66052 12852 67564
rect 12908 66276 12964 66286
rect 13020 66276 13076 69356
rect 15260 69412 15316 69422
rect 15260 69318 15316 69356
rect 16604 69410 16660 69422
rect 16604 69358 16606 69410
rect 16658 69358 16660 69410
rect 15820 69186 15876 69198
rect 15820 69134 15822 69186
rect 15874 69134 15876 69186
rect 13692 68626 13748 68638
rect 13692 68574 13694 68626
rect 13746 68574 13748 68626
rect 13244 68516 13300 68526
rect 13244 68422 13300 68460
rect 13580 67620 13636 67630
rect 13580 67526 13636 67564
rect 12908 66274 13076 66276
rect 12908 66222 12910 66274
rect 12962 66222 13076 66274
rect 12908 66220 13076 66222
rect 12908 66210 12964 66220
rect 12348 66050 12852 66052
rect 12348 65998 12350 66050
rect 12402 65998 12798 66050
rect 12850 65998 12852 66050
rect 12348 65996 12852 65998
rect 12348 65986 12404 65996
rect 10892 65538 10948 65548
rect 9324 64706 9492 64708
rect 9324 64654 9326 64706
rect 9378 64654 9492 64706
rect 9324 64652 9492 64654
rect 9324 64642 9380 64652
rect 9212 64428 9380 64484
rect 8988 63970 9044 63980
rect 4476 63532 4740 63542
rect 8876 63532 9044 63588
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4476 63466 4740 63476
rect 2492 63186 2548 63196
rect 1708 63026 1764 63038
rect 1708 62974 1710 63026
rect 1762 62974 1764 63026
rect 1708 62580 1764 62974
rect 2044 63028 2100 63038
rect 2044 62934 2100 62972
rect 8876 63028 8932 63038
rect 8876 62934 8932 62972
rect 8988 63026 9044 63532
rect 8988 62974 8990 63026
rect 9042 62974 9044 63026
rect 1708 62514 1764 62524
rect 2492 62914 2548 62926
rect 2492 62862 2494 62914
rect 2546 62862 2548 62914
rect 2492 62580 2548 62862
rect 2492 62514 2548 62524
rect 8092 62580 8148 62590
rect 8092 62486 8148 62524
rect 8988 62580 9044 62974
rect 9212 62916 9268 62926
rect 8988 62514 9044 62524
rect 9100 62914 9268 62916
rect 9100 62862 9214 62914
rect 9266 62862 9268 62914
rect 9100 62860 9268 62862
rect 7868 62354 7924 62366
rect 7868 62302 7870 62354
rect 7922 62302 7924 62354
rect 7868 62188 7924 62302
rect 8540 62354 8596 62366
rect 8540 62302 8542 62354
rect 8594 62302 8596 62354
rect 7868 62132 8484 62188
rect 4476 61964 4740 61974
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4476 61898 4740 61908
rect 8428 61572 8484 62132
rect 8316 61570 8484 61572
rect 8316 61518 8430 61570
rect 8482 61518 8484 61570
rect 8316 61516 8484 61518
rect 6076 60452 6132 60462
rect 4476 60396 4740 60406
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4476 60330 4740 60340
rect 6076 60002 6132 60396
rect 6076 59950 6078 60002
rect 6130 59950 6132 60002
rect 6076 59938 6132 59950
rect 1708 59892 1764 59902
rect 1708 59220 1764 59836
rect 2492 59892 2548 59902
rect 2492 59798 2548 59836
rect 6748 59892 6804 59902
rect 6748 59890 8036 59892
rect 6748 59838 6750 59890
rect 6802 59838 8036 59890
rect 6748 59836 8036 59838
rect 6748 59826 6804 59836
rect 2044 59780 2100 59790
rect 2044 59686 2100 59724
rect 7980 59442 8036 59836
rect 7980 59390 7982 59442
rect 8034 59390 8036 59442
rect 7980 59378 8036 59390
rect 1708 59154 1764 59164
rect 7868 59218 7924 59230
rect 7868 59166 7870 59218
rect 7922 59166 7924 59218
rect 4476 58828 4740 58838
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4476 58762 4740 58772
rect 1708 58322 1764 58334
rect 1708 58270 1710 58322
rect 1762 58270 1764 58322
rect 1708 57876 1764 58270
rect 7868 58324 7924 59166
rect 8204 59220 8260 59230
rect 8204 59126 8260 59164
rect 7868 58268 8148 58324
rect 2044 58212 2100 58222
rect 2044 58118 2100 58156
rect 2492 58210 2548 58222
rect 2492 58158 2494 58210
rect 2546 58158 2548 58210
rect 1708 57810 1764 57820
rect 2492 57876 2548 58158
rect 2492 57810 2548 57820
rect 7756 58212 7812 58222
rect 2044 57764 2100 57774
rect 2044 57670 2100 57708
rect 7756 57762 7812 58156
rect 8092 57874 8148 58268
rect 8092 57822 8094 57874
rect 8146 57822 8148 57874
rect 8092 57810 8148 57822
rect 7756 57710 7758 57762
rect 7810 57710 7812 57762
rect 7756 57698 7812 57710
rect 7868 57762 7924 57774
rect 7868 57710 7870 57762
rect 7922 57710 7924 57762
rect 1708 57650 1764 57662
rect 1708 57598 1710 57650
rect 1762 57598 1764 57650
rect 1708 57204 1764 57598
rect 1708 57138 1764 57148
rect 2492 57538 2548 57550
rect 2492 57486 2494 57538
rect 2546 57486 2548 57538
rect 2492 57204 2548 57486
rect 4476 57260 4740 57270
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4476 57194 4740 57204
rect 2492 57138 2548 57148
rect 7868 56980 7924 57710
rect 7644 56924 7924 56980
rect 8316 56980 8372 61516
rect 8428 61506 8484 61516
rect 8540 61348 8596 62302
rect 8764 62354 8820 62366
rect 8764 62302 8766 62354
rect 8818 62302 8820 62354
rect 8764 61796 8820 62302
rect 9100 62354 9156 62860
rect 9212 62850 9268 62860
rect 9100 62302 9102 62354
rect 9154 62302 9156 62354
rect 9100 62290 9156 62302
rect 8876 62244 8932 62282
rect 8876 62178 8932 62188
rect 8764 61730 8820 61740
rect 8876 61572 8932 61582
rect 9324 61572 9380 64428
rect 8876 61570 9380 61572
rect 8876 61518 8878 61570
rect 8930 61518 9380 61570
rect 8876 61516 9380 61518
rect 8876 61506 8932 61516
rect 9212 61348 9268 61358
rect 8540 61346 9268 61348
rect 8540 61294 9214 61346
rect 9266 61294 9268 61346
rect 8540 61292 9268 61294
rect 8428 59220 8484 59230
rect 8540 59220 8596 61292
rect 9212 61282 9268 61292
rect 8988 59780 9044 59790
rect 9212 59780 9268 59790
rect 8988 59778 9212 59780
rect 8988 59726 8990 59778
rect 9042 59726 9212 59778
rect 8988 59724 9212 59726
rect 8988 59714 9044 59724
rect 9212 59714 9268 59724
rect 8428 59218 8596 59220
rect 8428 59166 8430 59218
rect 8482 59166 8596 59218
rect 8428 59164 8596 59166
rect 8428 59154 8484 59164
rect 8316 56924 8484 56980
rect 1708 56754 1764 56766
rect 1708 56702 1710 56754
rect 1762 56702 1764 56754
rect 1708 56532 1764 56702
rect 7420 56754 7476 56766
rect 7420 56702 7422 56754
rect 7474 56702 7476 56754
rect 2044 56644 2100 56654
rect 2044 56642 2212 56644
rect 2044 56590 2046 56642
rect 2098 56590 2212 56642
rect 2044 56588 2212 56590
rect 2044 56578 2100 56588
rect 1708 56466 1764 56476
rect 2044 56308 2100 56318
rect 2044 56214 2100 56252
rect 2156 56196 2212 56588
rect 2492 56642 2548 56654
rect 2492 56590 2494 56642
rect 2546 56590 2548 56642
rect 2492 56532 2548 56590
rect 2492 56466 2548 56476
rect 7420 56308 7476 56702
rect 7420 56242 7476 56252
rect 7532 56644 7588 56654
rect 7644 56644 7700 56924
rect 7756 56756 7812 56766
rect 7980 56756 8036 56766
rect 7756 56754 8036 56756
rect 7756 56702 7758 56754
rect 7810 56702 7982 56754
rect 8034 56702 8036 56754
rect 7756 56700 8036 56702
rect 7756 56690 7812 56700
rect 7980 56690 8036 56700
rect 8316 56754 8372 56766
rect 8316 56702 8318 56754
rect 8370 56702 8372 56754
rect 7532 56642 7700 56644
rect 7532 56590 7534 56642
rect 7586 56590 7700 56642
rect 7532 56588 7700 56590
rect 8092 56642 8148 56654
rect 8092 56590 8094 56642
rect 8146 56590 8148 56642
rect 2156 56130 2212 56140
rect 1708 56082 1764 56094
rect 1708 56030 1710 56082
rect 1762 56030 1764 56082
rect 1708 55860 1764 56030
rect 5964 56082 6020 56094
rect 5964 56030 5966 56082
rect 6018 56030 6020 56082
rect 1708 55794 1764 55804
rect 2492 55970 2548 55982
rect 2492 55918 2494 55970
rect 2546 55918 2548 55970
rect 2492 55860 2548 55918
rect 2492 55794 2548 55804
rect 4476 55692 4740 55702
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4476 55626 4740 55636
rect 2044 55300 2100 55310
rect 5964 55300 6020 56030
rect 7532 56084 7588 56588
rect 7532 56028 7924 56084
rect 6636 55972 6692 55982
rect 6636 55878 6692 55916
rect 7644 55748 7700 55758
rect 6300 55524 6356 55534
rect 6300 55300 6356 55468
rect 5964 55298 6356 55300
rect 5964 55246 6302 55298
rect 6354 55246 6356 55298
rect 5964 55244 6356 55246
rect 1708 55188 1764 55198
rect 1708 55094 1764 55132
rect 2044 55186 2100 55244
rect 2044 55134 2046 55186
rect 2098 55134 2100 55186
rect 2044 55122 2100 55134
rect 2492 55188 2548 55198
rect 2492 55094 2548 55132
rect 4476 54124 4740 54134
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4476 54058 4740 54068
rect 1708 53506 1764 53518
rect 1708 53454 1710 53506
rect 1762 53454 1764 53506
rect 1708 53172 1764 53454
rect 2044 53508 2100 53518
rect 2044 53506 2212 53508
rect 2044 53454 2046 53506
rect 2098 53454 2212 53506
rect 2044 53452 2212 53454
rect 2044 53442 2100 53452
rect 1708 53106 1764 53116
rect 1708 52162 1764 52174
rect 1708 52110 1710 52162
rect 1762 52110 1764 52162
rect 1708 51828 1764 52110
rect 2044 52164 2100 52174
rect 2044 52050 2100 52108
rect 2044 51998 2046 52050
rect 2098 51998 2100 52050
rect 2044 51986 2100 51998
rect 2156 52052 2212 53452
rect 2492 53506 2548 53518
rect 2492 53454 2494 53506
rect 2546 53454 2548 53506
rect 2492 53172 2548 53454
rect 2492 53106 2548 53116
rect 4476 52556 4740 52566
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4476 52490 4740 52500
rect 2156 51986 2212 51996
rect 2492 52162 2548 52174
rect 2492 52110 2494 52162
rect 2546 52110 2548 52162
rect 1708 51762 1764 51772
rect 2492 51828 2548 52110
rect 2492 51762 2548 51772
rect 2044 51492 2100 51502
rect 2044 51398 2100 51436
rect 1708 51378 1764 51390
rect 6188 51380 6244 55244
rect 6300 55234 6356 55244
rect 6972 55188 7028 55198
rect 6972 55094 7028 55132
rect 7644 54628 7700 55692
rect 7756 54628 7812 54638
rect 7644 54626 7812 54628
rect 7644 54574 7758 54626
rect 7810 54574 7812 54626
rect 7644 54572 7812 54574
rect 7756 54562 7812 54572
rect 7868 54626 7924 56028
rect 8092 55188 8148 56590
rect 8092 55122 8148 55132
rect 8204 56084 8260 56094
rect 8092 54740 8148 54750
rect 8204 54740 8260 56028
rect 8316 55412 8372 56702
rect 8316 55346 8372 55356
rect 8428 55188 8484 56924
rect 8540 56754 8596 59164
rect 8540 56702 8542 56754
rect 8594 56702 8596 56754
rect 8540 56196 8596 56702
rect 8540 56130 8596 56140
rect 8652 58212 8708 58222
rect 8092 54738 8260 54740
rect 8092 54686 8094 54738
rect 8146 54686 8260 54738
rect 8092 54684 8260 54686
rect 8316 55132 8484 55188
rect 8652 55300 8708 58156
rect 8092 54674 8148 54684
rect 7868 54574 7870 54626
rect 7922 54574 7924 54626
rect 7868 53732 7924 54574
rect 7868 53666 7924 53676
rect 1708 51326 1710 51378
rect 1762 51326 1764 51378
rect 1708 51156 1764 51326
rect 5852 51378 6244 51380
rect 5852 51326 6190 51378
rect 6242 51326 6244 51378
rect 5852 51324 6244 51326
rect 1708 51090 1764 51100
rect 2492 51266 2548 51278
rect 2492 51214 2494 51266
rect 2546 51214 2548 51266
rect 2492 51156 2548 51214
rect 2492 51090 2548 51100
rect 4476 50988 4740 50998
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4476 50922 4740 50932
rect 2716 50596 2772 50606
rect 1708 50484 1764 50494
rect 1708 50390 1764 50428
rect 2380 50482 2436 50494
rect 2380 50430 2382 50482
rect 2434 50430 2436 50482
rect 2044 50372 2100 50382
rect 2044 50278 2100 50316
rect 2044 49924 2100 49934
rect 2044 49830 2100 49868
rect 1708 49810 1764 49822
rect 1708 49758 1710 49810
rect 1762 49758 1764 49810
rect 1708 49700 1764 49758
rect 2380 49812 2436 50430
rect 2492 50484 2548 50494
rect 2492 50034 2548 50428
rect 2716 50482 2772 50540
rect 2716 50430 2718 50482
rect 2770 50430 2772 50482
rect 2716 50418 2772 50430
rect 3164 50482 3220 50494
rect 3164 50430 3166 50482
rect 3218 50430 3220 50482
rect 2492 49982 2494 50034
rect 2546 49982 2548 50034
rect 2492 49970 2548 49982
rect 2380 49746 2436 49756
rect 3164 49812 3220 50430
rect 3164 49746 3220 49756
rect 5292 49812 5348 49822
rect 5852 49812 5908 51324
rect 6188 51314 6244 51324
rect 6860 51268 6916 51278
rect 6860 51266 7476 51268
rect 6860 51214 6862 51266
rect 6914 51214 7476 51266
rect 6860 51212 7476 51214
rect 6860 51202 6916 51212
rect 7420 50594 7476 51212
rect 7420 50542 7422 50594
rect 7474 50542 7476 50594
rect 7420 50530 7476 50542
rect 7756 50484 7812 50522
rect 8316 50482 8372 55132
rect 8652 54516 8708 55244
rect 8652 54450 8708 54460
rect 8764 55970 8820 55982
rect 8764 55918 8766 55970
rect 8818 55918 8820 55970
rect 8764 54514 8820 55918
rect 9100 55860 9156 55870
rect 8988 55804 9100 55860
rect 9324 55860 9380 61516
rect 9436 62356 9492 64652
rect 9884 65436 10164 65492
rect 9884 64148 9940 65436
rect 11340 64820 11396 64830
rect 9996 64596 10052 64606
rect 9996 64594 10500 64596
rect 9996 64542 9998 64594
rect 10050 64542 10500 64594
rect 9996 64540 10500 64542
rect 9996 64530 10052 64540
rect 10108 64372 10164 64382
rect 9996 64148 10052 64158
rect 9884 64146 10052 64148
rect 9884 64094 9998 64146
rect 10050 64094 10052 64146
rect 9884 64092 10052 64094
rect 9772 63924 9828 63934
rect 9996 63924 10052 64092
rect 9772 63922 9940 63924
rect 9772 63870 9774 63922
rect 9826 63870 9940 63922
rect 9772 63868 9940 63870
rect 9772 63858 9828 63868
rect 9884 63138 9940 63868
rect 9996 63858 10052 63868
rect 9884 63086 9886 63138
rect 9938 63086 9940 63138
rect 9548 62356 9604 62366
rect 9436 62354 9604 62356
rect 9436 62302 9550 62354
rect 9602 62302 9604 62354
rect 9436 62300 9604 62302
rect 9436 60452 9492 62300
rect 9548 62290 9604 62300
rect 9884 62188 9940 63086
rect 9436 60386 9492 60396
rect 9548 62132 9940 62188
rect 10108 62188 10164 64316
rect 10444 64146 10500 64540
rect 11116 64148 11172 64158
rect 10444 64094 10446 64146
rect 10498 64094 10500 64146
rect 10444 64082 10500 64094
rect 10780 64146 11172 64148
rect 10780 64094 11118 64146
rect 11170 64094 11172 64146
rect 10780 64092 11172 64094
rect 10220 64036 10276 64046
rect 10220 63922 10276 63980
rect 10668 64036 10724 64046
rect 10780 64036 10836 64092
rect 11116 64082 11172 64092
rect 11340 64146 11396 64764
rect 11340 64094 11342 64146
rect 11394 64094 11396 64146
rect 11340 64082 11396 64094
rect 10668 64034 10836 64036
rect 10668 63982 10670 64034
rect 10722 63982 10836 64034
rect 10668 63980 10836 63982
rect 10668 63970 10724 63980
rect 10220 63870 10222 63922
rect 10274 63870 10276 63922
rect 10220 63858 10276 63870
rect 10892 63924 10948 63934
rect 10892 63830 10948 63868
rect 11452 63922 11508 63934
rect 11452 63870 11454 63922
rect 11506 63870 11508 63922
rect 10220 62914 10276 62926
rect 10220 62862 10222 62914
rect 10274 62862 10276 62914
rect 10220 62468 10276 62862
rect 11452 62580 11508 63870
rect 11452 62514 11508 62524
rect 10220 62402 10276 62412
rect 11004 62468 11060 62478
rect 10332 62244 10388 62282
rect 11004 62188 11060 62412
rect 10108 62132 10276 62188
rect 10332 62178 10388 62188
rect 9548 61570 9604 62132
rect 9548 61518 9550 61570
rect 9602 61518 9604 61570
rect 9548 59444 9604 61518
rect 10108 61796 10164 61806
rect 10108 61570 10164 61740
rect 10108 61518 10110 61570
rect 10162 61518 10164 61570
rect 10108 61506 10164 61518
rect 9548 59378 9604 59388
rect 9660 61348 9716 61358
rect 10220 61348 10276 62132
rect 10780 62132 11060 62188
rect 12460 62242 12516 62254
rect 12460 62190 12462 62242
rect 12514 62190 12516 62242
rect 10444 61460 10500 61470
rect 10444 61366 10500 61404
rect 10332 61348 10388 61358
rect 10220 61292 10332 61348
rect 9660 59330 9716 61292
rect 10332 61254 10388 61292
rect 9660 59278 9662 59330
rect 9714 59278 9716 59330
rect 9436 59220 9492 59230
rect 9660 59220 9716 59278
rect 9436 59126 9492 59164
rect 9548 59164 9716 59220
rect 9772 59780 9828 59790
rect 9772 59220 9828 59724
rect 10332 59444 10388 59454
rect 9772 59218 9940 59220
rect 9772 59166 9774 59218
rect 9826 59166 9940 59218
rect 9772 59164 9940 59166
rect 9548 57764 9604 59164
rect 9772 59154 9828 59164
rect 9772 58212 9828 58250
rect 9772 58146 9828 58156
rect 9884 58100 9940 59164
rect 10108 58434 10164 58446
rect 10108 58382 10110 58434
rect 10162 58382 10164 58434
rect 10108 58212 10164 58382
rect 10332 58322 10388 59388
rect 10332 58270 10334 58322
rect 10386 58270 10388 58322
rect 10332 58258 10388 58270
rect 10108 58146 10164 58156
rect 9884 58044 10052 58100
rect 9884 57764 9940 57774
rect 9548 57762 9940 57764
rect 9548 57710 9886 57762
rect 9938 57710 9940 57762
rect 9548 57708 9940 57710
rect 9884 57698 9940 57708
rect 9436 56084 9492 56094
rect 9436 55990 9492 56028
rect 9772 56082 9828 56094
rect 9772 56030 9774 56082
rect 9826 56030 9828 56082
rect 9660 55972 9716 55982
rect 9660 55878 9716 55916
rect 9772 55860 9828 56030
rect 9996 56084 10052 58044
rect 10220 57652 10276 57662
rect 10220 57650 10388 57652
rect 10220 57598 10222 57650
rect 10274 57598 10388 57650
rect 10220 57596 10388 57598
rect 10220 57586 10276 57596
rect 10108 56196 10164 56206
rect 10108 56102 10164 56140
rect 9996 56018 10052 56028
rect 9324 55804 9492 55860
rect 8764 54462 8766 54514
rect 8818 54462 8820 54514
rect 8764 53620 8820 54462
rect 8764 53554 8820 53564
rect 8876 54740 8932 54750
rect 8988 54740 9044 55804
rect 9100 55794 9156 55804
rect 9100 55410 9156 55422
rect 9100 55358 9102 55410
rect 9154 55358 9156 55410
rect 9100 55300 9156 55358
rect 9324 55412 9380 55422
rect 9212 55300 9268 55310
rect 9100 55244 9212 55300
rect 9212 55234 9268 55244
rect 9324 55298 9380 55356
rect 9324 55246 9326 55298
rect 9378 55246 9380 55298
rect 9324 55234 9380 55246
rect 9100 54740 9156 54750
rect 9436 54740 9492 55804
rect 9772 55794 9828 55804
rect 9660 55300 9716 55310
rect 9716 55244 9940 55300
rect 9660 55206 9716 55244
rect 9548 55076 9604 55086
rect 9548 55074 9716 55076
rect 9548 55022 9550 55074
rect 9602 55022 9716 55074
rect 9548 55020 9716 55022
rect 9548 55010 9604 55020
rect 8988 54738 9156 54740
rect 8988 54686 9102 54738
rect 9154 54686 9156 54738
rect 8988 54684 9156 54686
rect 8876 54626 8932 54684
rect 9100 54674 9156 54684
rect 9324 54684 9492 54740
rect 9660 54740 9716 55020
rect 9772 54740 9828 54750
rect 9660 54684 9772 54740
rect 8876 54574 8878 54626
rect 8930 54574 8932 54626
rect 8540 52052 8596 52062
rect 8540 51380 8596 51996
rect 8540 50594 8596 51324
rect 8540 50542 8542 50594
rect 8594 50542 8596 50594
rect 8540 50530 8596 50542
rect 8316 50430 8318 50482
rect 8370 50430 8372 50482
rect 8316 50428 8372 50430
rect 7756 50418 7812 50428
rect 7644 50370 7700 50382
rect 7644 50318 7646 50370
rect 7698 50318 7700 50370
rect 5292 49810 5908 49812
rect 5292 49758 5294 49810
rect 5346 49758 5908 49810
rect 5292 49756 5908 49758
rect 7196 49924 7252 49934
rect 5292 49746 5348 49756
rect 1708 49140 1764 49644
rect 2940 49700 2996 49710
rect 2940 49606 2996 49644
rect 5964 49698 6020 49710
rect 5964 49646 5966 49698
rect 6018 49646 6020 49698
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 1708 49074 1764 49084
rect 1708 48914 1764 48926
rect 1708 48862 1710 48914
rect 1762 48862 1764 48914
rect 1708 48468 1764 48862
rect 2044 48916 2100 48926
rect 2044 48822 2100 48860
rect 1708 48402 1764 48412
rect 2492 48802 2548 48814
rect 2492 48750 2494 48802
rect 2546 48750 2548 48802
rect 2492 48468 2548 48750
rect 2492 48402 2548 48412
rect 5964 48468 6020 49646
rect 7196 49026 7252 49868
rect 7196 48974 7198 49026
rect 7250 48974 7252 49026
rect 7196 48962 7252 48974
rect 7532 49028 7588 49038
rect 7644 49028 7700 50318
rect 7532 49026 7700 49028
rect 7532 48974 7534 49026
rect 7586 48974 7700 49026
rect 7532 48972 7700 48974
rect 7868 50372 8372 50428
rect 7532 48962 7588 48972
rect 6636 48916 6692 48926
rect 7868 48916 7924 50372
rect 8764 50260 8820 50270
rect 8652 50204 8764 50260
rect 8204 49812 8260 49822
rect 8204 49698 8260 49756
rect 8204 49646 8206 49698
rect 8258 49646 8260 49698
rect 8204 49026 8260 49646
rect 8204 48974 8206 49026
rect 8258 48974 8260 49026
rect 8204 48962 8260 48974
rect 8652 49026 8708 50204
rect 8764 50194 8820 50204
rect 8876 50036 8932 54574
rect 9100 54516 9156 54526
rect 8988 51828 9044 51838
rect 8988 51266 9044 51772
rect 8988 51214 8990 51266
rect 9042 51214 9044 51266
rect 8988 51202 9044 51214
rect 8652 48974 8654 49026
rect 8706 48974 8708 49026
rect 6636 48822 6692 48860
rect 7644 48860 8148 48916
rect 6748 48802 6804 48814
rect 6972 48804 7028 48814
rect 6748 48750 6750 48802
rect 6802 48750 6804 48802
rect 5964 48402 6020 48412
rect 6636 48468 6692 48478
rect 6636 48374 6692 48412
rect 2044 48356 2100 48366
rect 2044 48262 2100 48300
rect 1708 48242 1764 48254
rect 1708 48190 1710 48242
rect 1762 48190 1764 48242
rect 1708 47796 1764 48190
rect 1708 47730 1764 47740
rect 2492 48130 2548 48142
rect 2492 48078 2494 48130
rect 2546 48078 2548 48130
rect 2492 47796 2548 48078
rect 6748 48132 6804 48750
rect 6860 48802 7028 48804
rect 6860 48750 6974 48802
rect 7026 48750 7028 48802
rect 6860 48748 7028 48750
rect 6860 48466 6916 48748
rect 6972 48738 7028 48748
rect 7084 48804 7140 48814
rect 6860 48414 6862 48466
rect 6914 48414 6916 48466
rect 6860 48402 6916 48414
rect 6972 48356 7028 48366
rect 7084 48356 7140 48748
rect 7308 48802 7364 48814
rect 7308 48750 7310 48802
rect 7362 48750 7364 48802
rect 7308 48356 7364 48750
rect 7644 48466 7700 48860
rect 7644 48414 7646 48466
rect 7698 48414 7700 48466
rect 7644 48402 7700 48414
rect 6972 48354 7140 48356
rect 6972 48302 6974 48354
rect 7026 48302 7140 48354
rect 6972 48300 7140 48302
rect 7196 48354 7364 48356
rect 7196 48302 7310 48354
rect 7362 48302 7364 48354
rect 7196 48300 7364 48302
rect 6972 48290 7028 48300
rect 7196 48132 7252 48300
rect 7308 48290 7364 48300
rect 7980 48356 8036 48366
rect 6748 48076 7252 48132
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 2492 47730 2548 47740
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 6524 45890 6580 45902
rect 6524 45838 6526 45890
rect 6578 45838 6580 45890
rect 2044 45220 2100 45230
rect 2044 45126 2100 45164
rect 1708 45106 1764 45118
rect 1708 45054 1710 45106
rect 1762 45054 1764 45106
rect 1708 44996 1764 45054
rect 1708 44436 1764 44940
rect 2492 44996 2548 45006
rect 2492 44902 2548 44940
rect 5964 44884 6020 44894
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 1708 44370 1764 44380
rect 1708 44210 1764 44222
rect 1708 44158 1710 44210
rect 1762 44158 1764 44210
rect 1708 43764 1764 44158
rect 2044 44100 2100 44110
rect 2044 44006 2100 44044
rect 2492 44098 2548 44110
rect 2492 44046 2494 44098
rect 2546 44046 2548 44098
rect 1708 43698 1764 43708
rect 2492 43764 2548 44046
rect 2492 43698 2548 43708
rect 5964 43650 6020 44828
rect 5964 43598 5966 43650
rect 6018 43598 6020 43650
rect 5964 43586 6020 43598
rect 5292 43540 5348 43550
rect 5292 43446 5348 43484
rect 6524 43540 6580 45838
rect 6636 45220 6692 45230
rect 6860 45220 6916 45230
rect 6636 44322 6692 45164
rect 6748 45218 6916 45220
rect 6748 45166 6862 45218
rect 6914 45166 6916 45218
rect 6748 45164 6916 45166
rect 6748 44546 6804 45164
rect 6860 45154 6916 45164
rect 6972 45106 7028 45118
rect 6972 45054 6974 45106
rect 7026 45054 7028 45106
rect 6860 44884 6916 44894
rect 6860 44790 6916 44828
rect 6972 44772 7028 45054
rect 6972 44706 7028 44716
rect 6748 44494 6750 44546
rect 6802 44494 6804 44546
rect 6748 44482 6804 44494
rect 6636 44270 6638 44322
rect 6690 44270 6692 44322
rect 6636 44258 6692 44270
rect 6748 44212 6804 44222
rect 7196 44212 7252 48076
rect 7980 47458 8036 48300
rect 7980 47406 7982 47458
rect 8034 47406 8036 47458
rect 7980 47394 8036 47406
rect 8092 47346 8148 48860
rect 8428 48804 8484 48814
rect 8428 48710 8484 48748
rect 8092 47294 8094 47346
rect 8146 47294 8148 47346
rect 8092 47282 8148 47294
rect 8316 47234 8372 47246
rect 8316 47182 8318 47234
rect 8370 47182 8372 47234
rect 8316 46788 8372 47182
rect 8428 46788 8484 46798
rect 8316 46786 8484 46788
rect 8316 46734 8430 46786
rect 8482 46734 8484 46786
rect 8316 46732 8484 46734
rect 8428 46722 8484 46732
rect 7308 46564 7364 46574
rect 7308 46002 7364 46508
rect 8540 46564 8596 46574
rect 8540 46470 8596 46508
rect 7308 45950 7310 46002
rect 7362 45950 7364 46002
rect 7308 45938 7364 45950
rect 8092 44772 8148 44782
rect 8148 44716 8372 44772
rect 8092 44706 8148 44716
rect 8316 44434 8372 44716
rect 8316 44382 8318 44434
rect 8370 44382 8372 44434
rect 8316 44370 8372 44382
rect 8540 44324 8596 44334
rect 8652 44324 8708 48974
rect 8764 49980 8932 50036
rect 8764 47012 8820 49980
rect 9100 49812 9156 54460
rect 9100 49746 9156 49756
rect 8876 48914 8932 48926
rect 8876 48862 8878 48914
rect 8930 48862 8932 48914
rect 8876 47348 8932 48862
rect 8876 47282 8932 47292
rect 9212 47236 9268 47246
rect 8988 47234 9268 47236
rect 8988 47182 9214 47234
rect 9266 47182 9268 47234
rect 8988 47180 9268 47182
rect 8876 47012 8932 47022
rect 8764 46956 8876 47012
rect 8876 46946 8932 46956
rect 8764 46788 8820 46798
rect 8764 46694 8820 46732
rect 8988 46676 9044 47180
rect 9212 47170 9268 47180
rect 8988 46582 9044 46620
rect 8988 45332 9044 45342
rect 9212 45332 9268 45342
rect 8988 45330 9212 45332
rect 8988 45278 8990 45330
rect 9042 45278 9212 45330
rect 8988 45276 9212 45278
rect 8988 45266 9044 45276
rect 9212 45266 9268 45276
rect 8540 44322 8708 44324
rect 8540 44270 8542 44322
rect 8594 44270 8708 44322
rect 8540 44268 8708 44270
rect 8764 45220 8820 45230
rect 8764 44322 8820 45164
rect 8764 44270 8766 44322
rect 8818 44270 8820 44322
rect 7532 44212 7588 44222
rect 6748 44210 7588 44212
rect 6748 44158 6750 44210
rect 6802 44158 7534 44210
rect 7586 44158 7588 44210
rect 6748 44156 7588 44158
rect 6748 44146 6804 44156
rect 7532 44146 7588 44156
rect 8204 44210 8260 44222
rect 8204 44158 8206 44210
rect 8258 44158 8260 44210
rect 7644 44100 7700 44110
rect 7644 44006 7700 44044
rect 7868 44098 7924 44110
rect 7868 44046 7870 44098
rect 7922 44046 7924 44098
rect 7868 43708 7924 44046
rect 8204 43764 8260 44158
rect 7868 43652 8148 43708
rect 8204 43698 8260 43708
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 6524 42756 6580 43484
rect 6524 42690 6580 42700
rect 7084 42756 7140 42766
rect 7084 42662 7140 42700
rect 7756 42644 7812 42654
rect 7756 42642 8036 42644
rect 7756 42590 7758 42642
rect 7810 42590 8036 42642
rect 7756 42588 8036 42590
rect 7756 42578 7812 42588
rect 7980 42194 8036 42588
rect 7980 42142 7982 42194
rect 8034 42142 8036 42194
rect 7980 42130 8036 42142
rect 8092 42196 8148 43652
rect 8316 42532 8372 42542
rect 8204 42196 8260 42206
rect 8092 42194 8260 42196
rect 8092 42142 8206 42194
rect 8258 42142 8260 42194
rect 8092 42140 8260 42142
rect 8204 42130 8260 42140
rect 8316 42082 8372 42476
rect 8316 42030 8318 42082
rect 8370 42030 8372 42082
rect 8316 42018 8372 42030
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 1820 41186 1876 41198
rect 1820 41134 1822 41186
rect 1874 41134 1876 41186
rect 1820 41076 1876 41134
rect 1708 40402 1764 40414
rect 1708 40350 1710 40402
rect 1762 40350 1764 40402
rect 1708 40292 1764 40350
rect 1820 40404 1876 41020
rect 2492 41076 2548 41086
rect 2492 40982 2548 41020
rect 2044 40964 2100 40974
rect 2044 40870 2100 40908
rect 1820 40338 1876 40348
rect 2044 40514 2100 40526
rect 2044 40462 2046 40514
rect 2098 40462 2100 40514
rect 1708 39732 1764 40236
rect 1708 39666 1764 39676
rect 2044 39620 2100 40462
rect 2492 40402 2548 40414
rect 2492 40350 2494 40402
rect 2546 40350 2548 40402
rect 2492 40292 2548 40350
rect 2492 40226 2548 40236
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 2044 39554 2100 39564
rect 8540 39620 8596 44268
rect 8764 44258 8820 44270
rect 9324 43708 9380 54684
rect 9772 54646 9828 54684
rect 9548 53732 9604 53742
rect 9436 51828 9492 51838
rect 9436 50594 9492 51772
rect 9548 51490 9604 53676
rect 9548 51438 9550 51490
rect 9602 51438 9604 51490
rect 9548 51156 9604 51438
rect 9772 51940 9828 51950
rect 9772 51380 9828 51884
rect 9884 51716 9940 55244
rect 10332 55188 10388 57596
rect 10108 55186 10388 55188
rect 10108 55134 10334 55186
rect 10386 55134 10388 55186
rect 10108 55132 10388 55134
rect 10108 54738 10164 55132
rect 10332 55122 10388 55132
rect 10556 55298 10612 55310
rect 10556 55246 10558 55298
rect 10610 55246 10612 55298
rect 10108 54686 10110 54738
rect 10162 54686 10164 54738
rect 9996 51716 10052 51726
rect 9884 51660 9996 51716
rect 9996 51650 10052 51660
rect 10108 51492 10164 54686
rect 10556 55076 10612 55246
rect 10332 53172 10388 53182
rect 10556 53172 10612 55020
rect 10332 53170 10612 53172
rect 10332 53118 10334 53170
rect 10386 53118 10612 53170
rect 10332 53116 10612 53118
rect 10332 53106 10388 53116
rect 10220 52834 10276 52846
rect 10220 52782 10222 52834
rect 10274 52782 10276 52834
rect 10220 51940 10276 52782
rect 10220 51874 10276 51884
rect 10220 51602 10276 51614
rect 10220 51550 10222 51602
rect 10274 51550 10276 51602
rect 10220 51492 10276 51550
rect 10556 51492 10612 51502
rect 10108 51436 10500 51492
rect 9828 51324 10276 51380
rect 9772 51286 9828 51324
rect 9548 51100 9940 51156
rect 9436 50542 9438 50594
rect 9490 50542 9492 50594
rect 9436 50530 9492 50542
rect 9660 50596 9716 50606
rect 9548 50484 9604 50522
rect 9548 50418 9604 50428
rect 9660 50148 9716 50540
rect 9772 50484 9828 50522
rect 9772 50418 9828 50428
rect 9884 50148 9940 51100
rect 9548 50092 9716 50148
rect 9772 50092 9940 50148
rect 9996 50482 10052 50494
rect 9996 50430 9998 50482
rect 10050 50430 10052 50482
rect 9548 49922 9604 50092
rect 9548 49870 9550 49922
rect 9602 49870 9604 49922
rect 9548 49858 9604 49870
rect 9660 49924 9716 49934
rect 9772 49924 9828 50092
rect 9660 49922 9828 49924
rect 9660 49870 9662 49922
rect 9714 49870 9828 49922
rect 9660 49868 9828 49870
rect 9996 49924 10052 50430
rect 10220 50036 10276 51324
rect 10444 50596 10500 51436
rect 10556 51490 10724 51492
rect 10556 51438 10558 51490
rect 10610 51438 10724 51490
rect 10556 51436 10724 51438
rect 10556 51426 10612 51436
rect 10556 50596 10612 50606
rect 10444 50594 10612 50596
rect 10444 50542 10558 50594
rect 10610 50542 10612 50594
rect 10444 50540 10612 50542
rect 10556 50530 10612 50540
rect 10668 50484 10724 51436
rect 10668 50418 10724 50428
rect 10332 50370 10388 50382
rect 10332 50318 10334 50370
rect 10386 50318 10388 50370
rect 10332 50260 10388 50318
rect 10332 50194 10388 50204
rect 10444 50036 10500 50046
rect 10220 50034 10500 50036
rect 10220 49982 10446 50034
rect 10498 49982 10500 50034
rect 10220 49980 10500 49982
rect 10444 49970 10500 49980
rect 9996 49868 10164 49924
rect 9660 49858 9716 49868
rect 9884 49812 9940 49822
rect 9884 49810 10052 49812
rect 9884 49758 9886 49810
rect 9938 49758 10052 49810
rect 9884 49756 10052 49758
rect 9884 49746 9940 49756
rect 9772 49700 9828 49710
rect 9772 49140 9828 49644
rect 9884 49140 9940 49150
rect 9772 49138 9940 49140
rect 9772 49086 9886 49138
rect 9938 49086 9940 49138
rect 9772 49084 9940 49086
rect 9660 47012 9716 47022
rect 9436 46788 9492 46798
rect 9436 46694 9492 46732
rect 9660 46786 9716 46956
rect 9660 46734 9662 46786
rect 9714 46734 9716 46786
rect 9436 46002 9492 46014
rect 9436 45950 9438 46002
rect 9490 45950 9492 46002
rect 9436 45556 9492 45950
rect 9660 45780 9716 46734
rect 9660 45714 9716 45724
rect 9772 46674 9828 46686
rect 9772 46622 9774 46674
rect 9826 46622 9828 46674
rect 9772 45556 9828 46622
rect 9436 45500 9828 45556
rect 9436 44212 9492 45500
rect 9436 44146 9492 44156
rect 9884 45332 9940 49084
rect 9996 47460 10052 49756
rect 10108 48580 10164 49868
rect 10220 49812 10276 49822
rect 10220 49718 10276 49756
rect 10556 49586 10612 49598
rect 10556 49534 10558 49586
rect 10610 49534 10612 49586
rect 10108 48524 10276 48580
rect 9996 47404 10164 47460
rect 10108 46674 10164 47404
rect 10108 46622 10110 46674
rect 10162 46622 10164 46674
rect 10108 46610 10164 46622
rect 10220 47348 10276 48524
rect 10556 48468 10612 49534
rect 10556 48402 10612 48412
rect 9884 43762 9940 45276
rect 10108 45890 10164 45902
rect 10108 45838 10110 45890
rect 10162 45838 10164 45890
rect 10108 44324 10164 45838
rect 10220 45220 10276 47292
rect 10444 46900 10500 46910
rect 10780 46900 10836 62132
rect 12460 61348 12516 62190
rect 12460 61282 12516 61292
rect 11788 60674 11844 60686
rect 11788 60622 11790 60674
rect 11842 60622 11844 60674
rect 11788 60452 11844 60622
rect 11788 60386 11844 60396
rect 12236 60452 12292 60462
rect 11116 59444 11172 59454
rect 11116 59350 11172 59388
rect 11452 59330 11508 59342
rect 11452 59278 11454 59330
rect 11506 59278 11508 59330
rect 11452 58660 11508 59278
rect 12236 59218 12292 60396
rect 12236 59166 12238 59218
rect 12290 59166 12292 59218
rect 12236 59154 12292 59166
rect 11452 58594 11508 58604
rect 12572 57652 12628 65996
rect 12796 65986 12852 65996
rect 13692 64820 13748 68574
rect 14476 68516 14532 68526
rect 14252 68514 14532 68516
rect 14252 68462 14478 68514
rect 14530 68462 14532 68514
rect 14252 68460 14532 68462
rect 14140 67844 14196 67854
rect 13916 67788 14140 67844
rect 13916 67282 13972 67788
rect 14140 67750 14196 67788
rect 13916 67230 13918 67282
rect 13970 67230 13972 67282
rect 13916 67218 13972 67230
rect 13916 66836 13972 66846
rect 13580 64764 13748 64820
rect 13804 66780 13916 66836
rect 13356 64708 13412 64718
rect 12684 64482 12740 64494
rect 12684 64430 12686 64482
rect 12738 64430 12740 64482
rect 12684 62804 12740 64430
rect 13356 64148 13412 64652
rect 12684 62738 12740 62748
rect 13244 64146 13412 64148
rect 13244 64094 13358 64146
rect 13410 64094 13412 64146
rect 13244 64092 13412 64094
rect 13244 62578 13300 64092
rect 13356 64082 13412 64092
rect 13244 62526 13246 62578
rect 13298 62526 13300 62578
rect 13244 62468 13300 62526
rect 13244 62402 13300 62412
rect 13580 63138 13636 64764
rect 13804 64708 13860 66780
rect 13916 66770 13972 66780
rect 13692 64652 13860 64708
rect 14028 64706 14084 64718
rect 14028 64654 14030 64706
rect 14082 64654 14084 64706
rect 13692 64594 13748 64652
rect 13692 64542 13694 64594
rect 13746 64542 13748 64594
rect 13692 64530 13748 64542
rect 13916 64034 13972 64046
rect 13916 63982 13918 64034
rect 13970 63982 13972 64034
rect 13916 63924 13972 63982
rect 13692 63812 13748 63822
rect 13692 63718 13748 63756
rect 13804 63810 13860 63822
rect 13804 63758 13806 63810
rect 13858 63758 13860 63810
rect 13804 63252 13860 63758
rect 13580 63086 13582 63138
rect 13634 63086 13636 63138
rect 13580 62188 13636 63086
rect 13692 63196 13860 63252
rect 13916 63252 13972 63868
rect 14028 63700 14084 64654
rect 14140 64708 14196 64746
rect 14140 64642 14196 64652
rect 14140 64484 14196 64494
rect 14252 64484 14308 68460
rect 14476 68450 14532 68460
rect 15820 68516 15876 69134
rect 15484 67844 15540 67854
rect 15484 67750 15540 67788
rect 15820 67844 15876 68460
rect 15820 67778 15876 67788
rect 16604 68514 16660 69358
rect 16604 68462 16606 68514
rect 16658 68462 16660 68514
rect 14476 67732 14532 67742
rect 14476 67618 14532 67676
rect 16604 67732 16660 68462
rect 16828 69188 16884 69198
rect 17388 69188 17444 70140
rect 17948 70130 18004 70140
rect 16828 69186 17444 69188
rect 16828 69134 16830 69186
rect 16882 69134 17444 69186
rect 16828 69132 17444 69134
rect 16604 67666 16660 67676
rect 16716 67956 16772 67966
rect 16716 67730 16772 67900
rect 16716 67678 16718 67730
rect 16770 67678 16772 67730
rect 16716 67666 16772 67678
rect 14476 67566 14478 67618
rect 14530 67566 14532 67618
rect 14476 67554 14532 67566
rect 16268 67618 16324 67630
rect 16268 67566 16270 67618
rect 16322 67566 16324 67618
rect 14140 64482 14308 64484
rect 14140 64430 14142 64482
rect 14194 64430 14308 64482
rect 14140 64428 14308 64430
rect 14476 64706 14532 64718
rect 14476 64654 14478 64706
rect 14530 64654 14532 64706
rect 14140 64418 14196 64428
rect 14476 64146 14532 64654
rect 14476 64094 14478 64146
rect 14530 64094 14532 64146
rect 14476 64082 14532 64094
rect 14588 64034 14644 64046
rect 14588 63982 14590 64034
rect 14642 63982 14644 64034
rect 14588 63924 14644 63982
rect 14588 63858 14644 63868
rect 14028 63644 14196 63700
rect 13916 63196 14084 63252
rect 13692 62354 13748 63196
rect 13692 62302 13694 62354
rect 13746 62302 13748 62354
rect 13692 62290 13748 62302
rect 13916 62468 13972 62478
rect 13244 62132 13636 62188
rect 13804 62132 13860 62142
rect 13244 60452 13300 62132
rect 13580 61570 13636 61582
rect 13580 61518 13582 61570
rect 13634 61518 13636 61570
rect 13580 61348 13636 61518
rect 13804 61460 13860 62076
rect 13916 62130 13972 62412
rect 13916 62078 13918 62130
rect 13970 62078 13972 62130
rect 13916 62066 13972 62078
rect 13804 61366 13860 61404
rect 13580 61282 13636 61292
rect 13244 60386 13300 60396
rect 13468 59892 13524 59902
rect 13468 59798 13524 59836
rect 13356 59780 13412 59790
rect 12908 59106 12964 59118
rect 12908 59054 12910 59106
rect 12962 59054 12964 59106
rect 12908 58212 12964 59054
rect 12908 58146 12964 58156
rect 13020 57764 13076 57774
rect 13020 57670 13076 57708
rect 13356 57652 13412 59724
rect 13580 59778 13636 59790
rect 13580 59726 13582 59778
rect 13634 59726 13636 59778
rect 13580 58434 13636 59726
rect 13692 59780 13748 59790
rect 14028 59780 14084 63196
rect 13748 59724 14084 59780
rect 14140 62466 14196 63644
rect 14364 63698 14420 63710
rect 14364 63646 14366 63698
rect 14418 63646 14420 63698
rect 14364 63364 14420 63646
rect 14364 63298 14420 63308
rect 14252 63026 14308 63038
rect 14252 62974 14254 63026
rect 14306 62974 14308 63026
rect 14252 62578 14308 62974
rect 15708 63028 15764 63038
rect 14924 62804 14980 62814
rect 14252 62526 14254 62578
rect 14306 62526 14308 62578
rect 14252 62514 14308 62526
rect 14700 62580 14756 62590
rect 14700 62486 14756 62524
rect 14140 62414 14142 62466
rect 14194 62414 14196 62466
rect 13692 59686 13748 59724
rect 13580 58382 13582 58434
rect 13634 58382 13636 58434
rect 13580 58370 13636 58382
rect 13692 58660 13748 58670
rect 13468 58212 13524 58222
rect 13468 58118 13524 58156
rect 12236 57596 12628 57652
rect 13132 57650 13412 57652
rect 13132 57598 13358 57650
rect 13410 57598 13412 57650
rect 13132 57596 13412 57598
rect 12012 56644 12068 56654
rect 11900 56642 12068 56644
rect 11900 56590 12014 56642
rect 12066 56590 12068 56642
rect 11900 56588 12068 56590
rect 11564 55412 11620 55422
rect 11116 55356 11564 55412
rect 11004 55076 11060 55086
rect 11004 54982 11060 55020
rect 11116 49700 11172 55356
rect 11564 55318 11620 55356
rect 11900 55186 11956 56588
rect 12012 56578 12068 56588
rect 11900 55134 11902 55186
rect 11954 55134 11956 55186
rect 11900 55076 11956 55134
rect 11900 55010 11956 55020
rect 12012 55970 12068 55982
rect 12012 55918 12014 55970
rect 12066 55918 12068 55970
rect 12012 55524 12068 55918
rect 12012 54514 12068 55468
rect 12236 55412 12292 57596
rect 13132 57540 13188 57596
rect 13356 57586 13412 57596
rect 12348 57484 13188 57540
rect 12348 56754 12404 57484
rect 13356 57426 13412 57438
rect 13356 57374 13358 57426
rect 13410 57374 13412 57426
rect 12348 56702 12350 56754
rect 12402 56702 12404 56754
rect 12348 56690 12404 56702
rect 12908 56868 12964 56878
rect 13356 56868 13412 57374
rect 13692 57090 13748 58604
rect 13692 57038 13694 57090
rect 13746 57038 13748 57090
rect 13468 56868 13524 56878
rect 13356 56866 13524 56868
rect 13356 56814 13470 56866
rect 13522 56814 13524 56866
rect 13356 56812 13524 56814
rect 12236 55346 12292 55356
rect 12684 56644 12740 56654
rect 12012 54462 12014 54514
rect 12066 54462 12068 54514
rect 11788 52274 11844 52286
rect 11788 52222 11790 52274
rect 11842 52222 11844 52274
rect 11452 52164 11508 52174
rect 11452 52070 11508 52108
rect 11788 52164 11844 52222
rect 11788 52098 11844 52108
rect 11676 51940 11732 51950
rect 11564 51884 11676 51940
rect 11452 51492 11508 51502
rect 11452 50818 11508 51436
rect 11452 50766 11454 50818
rect 11506 50766 11508 50818
rect 11452 50754 11508 50766
rect 11452 50484 11508 50494
rect 11228 50372 11284 50382
rect 11228 49922 11284 50316
rect 11228 49870 11230 49922
rect 11282 49870 11284 49922
rect 11228 49858 11284 49870
rect 11116 49644 11284 49700
rect 11116 48468 11172 48478
rect 10444 46898 10724 46900
rect 10444 46846 10446 46898
rect 10498 46846 10724 46898
rect 10444 46844 10724 46846
rect 10444 46834 10500 46844
rect 10556 46674 10612 46686
rect 10556 46622 10558 46674
rect 10610 46622 10612 46674
rect 10556 45330 10612 46622
rect 10556 45278 10558 45330
rect 10610 45278 10612 45330
rect 10556 45266 10612 45278
rect 10220 45126 10276 45164
rect 10668 44436 10724 46844
rect 10780 46786 10836 46844
rect 10780 46734 10782 46786
rect 10834 46734 10836 46786
rect 10780 46676 10836 46734
rect 10780 46610 10836 46620
rect 10892 48466 11172 48468
rect 10892 48414 11118 48466
rect 11170 48414 11172 48466
rect 10892 48412 11172 48414
rect 10780 46004 10836 46014
rect 10892 46004 10948 48412
rect 11116 48402 11172 48412
rect 10780 46002 10948 46004
rect 10780 45950 10782 46002
rect 10834 45950 10948 46002
rect 10780 45948 10948 45950
rect 10780 45938 10836 45948
rect 10780 45780 10836 45790
rect 10780 45330 10836 45724
rect 10780 45278 10782 45330
rect 10834 45278 10836 45330
rect 10780 45266 10836 45278
rect 10892 45108 10948 45118
rect 10892 45014 10948 45052
rect 10780 44436 10836 44446
rect 10668 44434 10836 44436
rect 10668 44382 10782 44434
rect 10834 44382 10836 44434
rect 10668 44380 10836 44382
rect 10780 44370 10836 44380
rect 10108 44322 10276 44324
rect 10108 44270 10110 44322
rect 10162 44270 10276 44322
rect 10108 44268 10276 44270
rect 10108 44258 10164 44268
rect 9884 43710 9886 43762
rect 9938 43710 9940 43762
rect 9884 43708 9940 43710
rect 9324 43652 9828 43708
rect 9884 43652 10164 43708
rect 9212 41300 9268 41310
rect 8764 39620 8820 39630
rect 9212 39620 9268 41244
rect 9660 40964 9716 40974
rect 9660 40514 9716 40908
rect 9772 40628 9828 43652
rect 10108 43650 10164 43652
rect 10108 43598 10110 43650
rect 10162 43598 10164 43650
rect 10108 43586 10164 43598
rect 9884 42868 9940 42878
rect 10220 42868 10276 44268
rect 9884 42774 9940 42812
rect 10108 42812 10276 42868
rect 10444 43650 10500 43662
rect 10444 43598 10446 43650
rect 10498 43598 10500 43650
rect 9772 40534 9828 40572
rect 10108 42756 10164 42812
rect 10108 41076 10164 42700
rect 10332 42756 10388 42766
rect 10444 42756 10500 43598
rect 10332 42754 10500 42756
rect 10332 42702 10334 42754
rect 10386 42702 10500 42754
rect 10332 42700 10500 42702
rect 10332 42690 10388 42700
rect 10444 41300 10500 42700
rect 10556 42868 10612 42878
rect 10556 42754 10612 42812
rect 10556 42702 10558 42754
rect 10610 42702 10612 42754
rect 10556 42690 10612 42702
rect 10892 42754 10948 42766
rect 10892 42702 10894 42754
rect 10946 42702 10948 42754
rect 10556 42532 10612 42542
rect 10892 42532 10948 42702
rect 11228 42532 11284 49644
rect 11340 49698 11396 49710
rect 11340 49646 11342 49698
rect 11394 49646 11396 49698
rect 11340 48242 11396 49646
rect 11340 48190 11342 48242
rect 11394 48190 11396 48242
rect 11340 48178 11396 48190
rect 11452 48244 11508 50428
rect 11564 50428 11620 51884
rect 11676 51846 11732 51884
rect 11788 51380 11844 51390
rect 12012 51380 12068 54462
rect 12236 55076 12292 55086
rect 12572 55076 12628 55086
rect 12236 55074 12628 55076
rect 12236 55022 12238 55074
rect 12290 55022 12574 55074
rect 12626 55022 12628 55074
rect 12236 55020 12628 55022
rect 12124 52164 12180 52174
rect 12124 52070 12180 52108
rect 12236 51940 12292 55020
rect 12572 55010 12628 55020
rect 12460 54852 12516 54862
rect 12460 52388 12516 54796
rect 12684 54626 12740 56588
rect 12908 55186 12964 56812
rect 13468 56802 13524 56812
rect 13468 56644 13524 56654
rect 13468 56550 13524 56588
rect 12908 55134 12910 55186
rect 12962 55134 12964 55186
rect 12908 55122 12964 55134
rect 13692 54852 13748 57038
rect 14028 58436 14084 58446
rect 14140 58436 14196 62414
rect 14364 62356 14420 62366
rect 14364 62262 14420 62300
rect 14924 62354 14980 62748
rect 15708 62466 15764 62972
rect 15708 62414 15710 62466
rect 15762 62414 15764 62466
rect 15708 62402 15764 62414
rect 16044 62804 16100 62814
rect 16044 62578 16100 62748
rect 16044 62526 16046 62578
rect 16098 62526 16100 62578
rect 14924 62302 14926 62354
rect 14978 62302 14980 62354
rect 14924 62290 14980 62302
rect 15596 62356 15652 62366
rect 15596 62262 15652 62300
rect 14812 61348 14868 61358
rect 14812 60002 14868 61292
rect 14812 59950 14814 60002
rect 14866 59950 14868 60002
rect 14812 59938 14868 59950
rect 14476 59892 14532 59902
rect 14476 59798 14532 59836
rect 15036 59892 15092 59902
rect 14364 59780 14420 59790
rect 14028 58434 14196 58436
rect 14028 58382 14030 58434
rect 14082 58382 14196 58434
rect 14028 58380 14196 58382
rect 14252 59778 14420 59780
rect 14252 59726 14366 59778
rect 14418 59726 14420 59778
rect 14252 59724 14420 59726
rect 14252 58436 14308 59724
rect 14364 59714 14420 59724
rect 15036 59106 15092 59836
rect 15932 59892 15988 59902
rect 16044 59892 16100 62526
rect 15932 59890 16100 59892
rect 15932 59838 15934 59890
rect 15986 59838 16100 59890
rect 15932 59836 16100 59838
rect 15932 59826 15988 59836
rect 15036 59054 15038 59106
rect 15090 59054 15092 59106
rect 15036 59042 15092 59054
rect 15820 59778 15876 59790
rect 15820 59726 15822 59778
rect 15874 59726 15876 59778
rect 14028 56868 14084 58380
rect 14252 58342 14308 58380
rect 15820 57764 15876 59726
rect 16268 59442 16324 67566
rect 16828 67170 16884 69132
rect 17388 68738 17444 69132
rect 17388 68686 17390 68738
rect 17442 68686 17444 68738
rect 17388 68674 17444 68686
rect 17612 69412 17668 69422
rect 17612 68850 17668 69356
rect 17612 68798 17614 68850
rect 17666 68798 17668 68850
rect 17612 68404 17668 68798
rect 17836 69410 17892 69422
rect 17836 69358 17838 69410
rect 17890 69358 17892 69410
rect 17724 68516 17780 68526
rect 17724 68422 17780 68460
rect 17612 68338 17668 68348
rect 16828 67118 16830 67170
rect 16882 67118 16884 67170
rect 16828 67106 16884 67118
rect 17388 67956 17444 67966
rect 17388 67170 17444 67900
rect 17836 67956 17892 69358
rect 17836 67890 17892 67900
rect 17724 67844 17780 67854
rect 17724 67228 17780 67788
rect 17948 67620 18004 67630
rect 17724 67172 17892 67228
rect 17388 67118 17390 67170
rect 17442 67118 17444 67170
rect 17388 67106 17444 67118
rect 17836 67058 17892 67172
rect 17836 67006 17838 67058
rect 17890 67006 17892 67058
rect 17836 66994 17892 67006
rect 16716 66836 16772 66846
rect 16716 66742 16772 66780
rect 17612 66836 17668 66846
rect 17948 66836 18004 67564
rect 18060 67058 18116 70140
rect 19852 70194 19908 70206
rect 19852 70142 19854 70194
rect 19906 70142 19908 70194
rect 18172 69970 18228 69982
rect 18172 69918 18174 69970
rect 18226 69918 18228 69970
rect 18172 69412 18228 69918
rect 18396 69970 18452 69982
rect 18396 69918 18398 69970
rect 18450 69918 18452 69970
rect 18396 69636 18452 69918
rect 18508 69972 18564 69982
rect 18508 69970 19124 69972
rect 18508 69918 18510 69970
rect 18562 69918 19124 69970
rect 18508 69916 19124 69918
rect 18508 69906 18564 69916
rect 18396 69580 18564 69636
rect 18172 69346 18228 69356
rect 18396 69410 18452 69422
rect 18396 69358 18398 69410
rect 18450 69358 18452 69410
rect 18172 67732 18228 67742
rect 18172 67638 18228 67676
rect 18060 67006 18062 67058
rect 18114 67006 18116 67058
rect 18060 66994 18116 67006
rect 18396 66948 18452 69358
rect 18508 68626 18564 69580
rect 19068 69410 19124 69916
rect 19068 69358 19070 69410
rect 19122 69358 19124 69410
rect 19068 69346 19124 69358
rect 19516 69636 19572 69646
rect 18508 68574 18510 68626
rect 18562 68574 18564 68626
rect 18508 67620 18564 68574
rect 18956 68628 19012 68638
rect 18956 68534 19012 68572
rect 18508 67554 18564 67564
rect 18396 66882 18452 66892
rect 18620 66948 18676 66958
rect 18620 66946 19012 66948
rect 18620 66894 18622 66946
rect 18674 66894 19012 66946
rect 18620 66892 19012 66894
rect 18620 66882 18676 66892
rect 17612 66834 18004 66836
rect 17612 66782 17614 66834
rect 17666 66782 18004 66834
rect 17612 66780 18004 66782
rect 17612 66770 17668 66780
rect 17948 64034 18004 64046
rect 17948 63982 17950 64034
rect 18002 63982 18004 64034
rect 17836 63252 17892 63262
rect 17388 63138 17444 63150
rect 17388 63086 17390 63138
rect 17442 63086 17444 63138
rect 16492 63028 16548 63038
rect 16492 62914 16548 62972
rect 17276 63028 17332 63038
rect 17276 62934 17332 62972
rect 16492 62862 16494 62914
rect 16546 62862 16548 62914
rect 16492 62850 16548 62862
rect 17388 62916 17444 63086
rect 16828 62580 16884 62590
rect 16828 62486 16884 62524
rect 17388 62356 17444 62860
rect 17836 63138 17892 63196
rect 17836 63086 17838 63138
rect 17890 63086 17892 63138
rect 17836 62692 17892 63086
rect 17836 62626 17892 62636
rect 17500 62580 17556 62590
rect 17948 62580 18004 63982
rect 18284 63922 18340 63934
rect 18284 63870 18286 63922
rect 18338 63870 18340 63922
rect 18284 63812 18340 63870
rect 18284 63746 18340 63756
rect 18956 63922 19012 66892
rect 19516 66836 19572 69580
rect 19852 69636 19908 70142
rect 19852 69570 19908 69580
rect 20076 70194 20132 70206
rect 20076 70142 20078 70194
rect 20130 70142 20132 70194
rect 20076 69524 20132 70142
rect 20076 69458 20132 69468
rect 20188 70194 20244 70206
rect 20188 70142 20190 70194
rect 20242 70142 20244 70194
rect 20188 69410 20244 70142
rect 20636 69972 20692 69982
rect 24444 69972 24500 69982
rect 20636 69970 21476 69972
rect 20636 69918 20638 69970
rect 20690 69918 21476 69970
rect 20636 69916 21476 69918
rect 20636 69906 20692 69916
rect 20636 69636 20692 69646
rect 20636 69542 20692 69580
rect 20412 69524 20468 69534
rect 20412 69430 20468 69468
rect 20188 69358 20190 69410
rect 20242 69358 20244 69410
rect 19628 69298 19684 69310
rect 19628 69246 19630 69298
rect 19682 69246 19684 69298
rect 19628 68852 19684 69246
rect 19836 69020 20100 69030
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 19836 68954 20100 68964
rect 20188 68852 20244 69358
rect 20748 69298 20804 69310
rect 20748 69246 20750 69298
rect 20802 69246 20804 69298
rect 19628 68786 19684 68796
rect 19740 68796 20244 68852
rect 20412 68852 20468 68862
rect 19628 68626 19684 68638
rect 19628 68574 19630 68626
rect 19682 68574 19684 68626
rect 19628 68516 19684 68574
rect 19628 68450 19684 68460
rect 19628 67956 19684 67966
rect 19740 67956 19796 68796
rect 19628 67954 19796 67956
rect 19628 67902 19630 67954
rect 19682 67902 19796 67954
rect 19628 67900 19796 67902
rect 20076 68404 20132 68414
rect 19628 67890 19684 67900
rect 20076 67842 20132 68348
rect 20076 67790 20078 67842
rect 20130 67790 20132 67842
rect 20076 67778 20132 67790
rect 20188 68402 20244 68414
rect 20188 68350 20190 68402
rect 20242 68350 20244 68402
rect 19836 67452 20100 67462
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 19836 67386 20100 67396
rect 20188 67170 20244 68350
rect 20188 67118 20190 67170
rect 20242 67118 20244 67170
rect 20188 67106 20244 67118
rect 20412 67058 20468 68796
rect 20524 68516 20580 68526
rect 20524 67954 20580 68460
rect 20524 67902 20526 67954
rect 20578 67902 20580 67954
rect 20524 67890 20580 67902
rect 20748 67228 20804 69246
rect 21084 68516 21140 68526
rect 21084 68422 21140 68460
rect 20748 67172 21364 67228
rect 20412 67006 20414 67058
rect 20466 67006 20468 67058
rect 20412 66994 20468 67006
rect 21308 67058 21364 67172
rect 21308 67006 21310 67058
rect 21362 67006 21364 67058
rect 21308 66994 21364 67006
rect 21420 66946 21476 69916
rect 22316 69524 22372 69534
rect 22316 69430 22372 69468
rect 23548 69524 23604 69534
rect 23212 68514 23268 68526
rect 23212 68462 23214 68514
rect 23266 68462 23268 68514
rect 23212 67282 23268 68462
rect 23212 67230 23214 67282
rect 23266 67230 23268 67282
rect 23212 67218 23268 67230
rect 23548 67842 23604 69468
rect 24444 69522 24500 69916
rect 25228 69972 25284 69982
rect 25228 69878 25284 69916
rect 24444 69470 24446 69522
rect 24498 69470 24500 69522
rect 24444 69458 24500 69470
rect 25228 69410 25284 69422
rect 25228 69358 25230 69410
rect 25282 69358 25284 69410
rect 25228 69076 25284 69358
rect 25452 69412 25508 70252
rect 25564 70084 25620 70094
rect 25564 69990 25620 70028
rect 26124 70084 26180 70094
rect 26124 69990 26180 70028
rect 27692 70084 27748 70094
rect 25564 69412 25620 69422
rect 25452 69410 25620 69412
rect 25452 69358 25566 69410
rect 25618 69358 25620 69410
rect 25452 69356 25620 69358
rect 25116 69020 25284 69076
rect 24668 68740 24724 68750
rect 24556 68684 24668 68740
rect 23996 68626 24052 68638
rect 23996 68574 23998 68626
rect 24050 68574 24052 68626
rect 23996 68180 24052 68574
rect 24332 68626 24388 68638
rect 24332 68574 24334 68626
rect 24386 68574 24388 68626
rect 24332 68516 24388 68574
rect 24332 68450 24388 68460
rect 23996 68114 24052 68124
rect 24556 67956 24612 68684
rect 24668 68646 24724 68684
rect 24556 67862 24612 67900
rect 24668 68516 24724 68526
rect 23548 67790 23550 67842
rect 23602 67790 23604 67842
rect 21420 66894 21422 66946
rect 21474 66894 21476 66946
rect 21420 66882 21476 66894
rect 22988 67058 23044 67070
rect 22988 67006 22990 67058
rect 23042 67006 23044 67058
rect 21196 66836 21252 66846
rect 19516 66770 19572 66780
rect 21084 66834 21252 66836
rect 21084 66782 21198 66834
rect 21250 66782 21252 66834
rect 21084 66780 21252 66782
rect 19836 65884 20100 65894
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 19836 65818 20100 65828
rect 19836 64316 20100 64326
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 19836 64250 20100 64260
rect 18956 63870 18958 63922
rect 19010 63870 19012 63922
rect 18060 63364 18116 63374
rect 18060 63270 18116 63308
rect 18956 63364 19012 63870
rect 20188 64034 20244 64046
rect 20188 63982 20190 64034
rect 20242 63982 20244 64034
rect 18956 63298 19012 63308
rect 19628 63810 19684 63822
rect 19628 63758 19630 63810
rect 19682 63758 19684 63810
rect 19404 63140 19460 63150
rect 19404 63046 19460 63084
rect 18396 63028 18452 63038
rect 17500 62578 17780 62580
rect 17500 62526 17502 62578
rect 17554 62526 17780 62578
rect 17500 62524 17780 62526
rect 17500 62514 17556 62524
rect 17612 62356 17668 62366
rect 17388 62354 17668 62356
rect 17388 62302 17614 62354
rect 17666 62302 17668 62354
rect 17388 62300 17668 62302
rect 17612 62244 17668 62300
rect 17612 62178 17668 62188
rect 17724 62356 17780 62524
rect 17612 61460 17668 61470
rect 16828 60786 16884 60798
rect 16828 60734 16830 60786
rect 16882 60734 16884 60786
rect 16828 60564 16884 60734
rect 17500 60674 17556 60686
rect 17500 60622 17502 60674
rect 17554 60622 17556 60674
rect 17500 60564 17556 60622
rect 16828 60508 17556 60564
rect 16268 59390 16270 59442
rect 16322 59390 16324 59442
rect 16268 58434 16324 59390
rect 16828 59220 16884 59230
rect 16828 59126 16884 59164
rect 16268 58382 16270 58434
rect 16322 58382 16324 58434
rect 16156 57764 16212 57774
rect 16268 57764 16324 58382
rect 16716 58322 16772 58334
rect 16716 58270 16718 58322
rect 16770 58270 16772 58322
rect 15820 57762 16100 57764
rect 15820 57710 15822 57762
rect 15874 57710 16100 57762
rect 15820 57708 16100 57710
rect 15820 57698 15876 57708
rect 14028 56774 14084 56812
rect 15036 57538 15092 57550
rect 15036 57486 15038 57538
rect 15090 57486 15092 57538
rect 15036 57428 15092 57486
rect 16044 57428 16100 57708
rect 16156 57762 16660 57764
rect 16156 57710 16158 57762
rect 16210 57710 16660 57762
rect 16156 57708 16660 57710
rect 16156 57698 16212 57708
rect 16380 57428 16436 57438
rect 16044 57426 16436 57428
rect 16044 57374 16382 57426
rect 16434 57374 16436 57426
rect 16044 57372 16436 57374
rect 14252 56756 14308 56766
rect 14252 56662 14308 56700
rect 13692 54786 13748 54796
rect 15036 55298 15092 57372
rect 16380 57362 16436 57372
rect 16604 57204 16660 57708
rect 16716 57652 16772 58270
rect 16716 57586 16772 57596
rect 16716 57426 16772 57438
rect 16716 57374 16718 57426
rect 16770 57374 16772 57426
rect 16716 57316 16772 57374
rect 16716 57260 16884 57316
rect 16604 57148 16772 57204
rect 16604 56980 16660 56990
rect 15596 56754 15652 56766
rect 15596 56702 15598 56754
rect 15650 56702 15652 56754
rect 15484 56644 15540 56654
rect 15484 56550 15540 56588
rect 15596 55524 15652 56702
rect 15036 55246 15038 55298
rect 15090 55246 15092 55298
rect 12684 54574 12686 54626
rect 12738 54574 12740 54626
rect 12684 54562 12740 54574
rect 14924 54738 14980 54750
rect 14924 54686 14926 54738
rect 14978 54686 14980 54738
rect 14924 54628 14980 54686
rect 14924 54562 14980 54572
rect 15036 53508 15092 55246
rect 15484 55468 15652 55524
rect 16268 56754 16324 56766
rect 16268 56702 16270 56754
rect 16322 56702 16324 56754
rect 15260 55074 15316 55086
rect 15260 55022 15262 55074
rect 15314 55022 15316 55074
rect 15036 53452 15204 53508
rect 15148 53060 15204 53452
rect 15260 53284 15316 55022
rect 15484 54628 15540 55468
rect 15484 54562 15540 54572
rect 15596 55300 15652 55310
rect 16268 55300 16324 56702
rect 16604 56082 16660 56924
rect 16716 56866 16772 57148
rect 16716 56814 16718 56866
rect 16770 56814 16772 56866
rect 16716 56802 16772 56814
rect 16604 56030 16606 56082
rect 16658 56030 16660 56082
rect 16604 56018 16660 56030
rect 15596 55298 16324 55300
rect 15596 55246 15598 55298
rect 15650 55246 16324 55298
rect 15596 55244 16324 55246
rect 16604 55860 16660 55870
rect 16828 55860 16884 57260
rect 17276 56980 17332 60508
rect 17612 60452 17668 61404
rect 17500 60396 17668 60452
rect 17388 59892 17444 59902
rect 17388 59798 17444 59836
rect 17500 59330 17556 60396
rect 17500 59278 17502 59330
rect 17554 59278 17556 59330
rect 17500 59266 17556 59278
rect 17724 59330 17780 62300
rect 17948 62354 18004 62524
rect 17948 62302 17950 62354
rect 18002 62302 18004 62354
rect 17948 62290 18004 62302
rect 18172 62914 18228 62926
rect 18172 62862 18174 62914
rect 18226 62862 18228 62914
rect 18172 61572 18228 62862
rect 18172 61506 18228 61516
rect 18396 60898 18452 62972
rect 18844 63026 18900 63038
rect 18844 62974 18846 63026
rect 18898 62974 18900 63026
rect 18844 62916 18900 62974
rect 18844 62850 18900 62860
rect 18732 62468 18788 62478
rect 18732 61460 18788 62412
rect 19516 62468 19572 62478
rect 19516 62374 19572 62412
rect 18956 62356 19012 62366
rect 19012 62300 19236 62356
rect 18956 62262 19012 62300
rect 18956 61908 19012 61918
rect 18956 61460 19012 61852
rect 19180 61572 19236 62300
rect 19292 62354 19348 62366
rect 19292 62302 19294 62354
rect 19346 62302 19348 62354
rect 19292 61908 19348 62302
rect 19628 62356 19684 63758
rect 19964 63698 20020 63710
rect 19964 63646 19966 63698
rect 20018 63646 20020 63698
rect 19964 63364 20020 63646
rect 19964 63298 20020 63308
rect 20188 63252 20244 63982
rect 20188 63186 20244 63196
rect 20300 63698 20356 63710
rect 20300 63646 20302 63698
rect 20354 63646 20356 63698
rect 20300 63138 20356 63646
rect 20300 63086 20302 63138
rect 20354 63086 20356 63138
rect 20300 63074 20356 63086
rect 20412 62916 20468 62926
rect 20300 62914 20468 62916
rect 20300 62862 20414 62914
rect 20466 62862 20468 62914
rect 20300 62860 20468 62862
rect 19836 62748 20100 62758
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 19836 62682 20100 62692
rect 19628 62290 19684 62300
rect 20188 62466 20244 62478
rect 20188 62414 20190 62466
rect 20242 62414 20244 62466
rect 19964 62244 20020 62254
rect 19852 62242 20020 62244
rect 19852 62190 19966 62242
rect 20018 62190 20020 62242
rect 19852 62188 20020 62190
rect 19628 62132 19684 62142
rect 19852 62132 20132 62188
rect 19628 62038 19684 62076
rect 19292 61842 19348 61852
rect 19964 61908 20020 61918
rect 19740 61796 19796 61806
rect 19740 61702 19796 61740
rect 19292 61628 19684 61684
rect 19292 61572 19348 61628
rect 19180 61570 19348 61572
rect 19180 61518 19294 61570
rect 19346 61518 19348 61570
rect 19180 61516 19348 61518
rect 19292 61506 19348 61516
rect 19628 61570 19684 61628
rect 19964 61572 20020 61852
rect 19628 61518 19630 61570
rect 19682 61518 19684 61570
rect 19628 61506 19684 61518
rect 19740 61516 20020 61572
rect 18732 61366 18788 61404
rect 18844 61458 19012 61460
rect 18844 61406 18958 61458
rect 19010 61406 19012 61458
rect 18844 61404 19012 61406
rect 18396 60846 18398 60898
rect 18450 60846 18452 60898
rect 17724 59278 17726 59330
rect 17778 59278 17780 59330
rect 17724 59266 17780 59278
rect 18172 60004 18228 60014
rect 18396 60004 18452 60846
rect 18732 60788 18788 60798
rect 18732 60694 18788 60732
rect 18508 60004 18564 60014
rect 18396 60002 18564 60004
rect 18396 59950 18510 60002
rect 18562 59950 18564 60002
rect 18396 59948 18564 59950
rect 18172 59442 18228 59948
rect 18508 59938 18564 59948
rect 18172 59390 18174 59442
rect 18226 59390 18228 59442
rect 17612 59220 17668 59230
rect 17500 58434 17556 58446
rect 17500 58382 17502 58434
rect 17554 58382 17556 58434
rect 17500 58212 17556 58382
rect 17500 58146 17556 58156
rect 17612 57988 17668 59164
rect 18172 58546 18228 59390
rect 18844 59442 18900 61404
rect 18956 61394 19012 61404
rect 19740 61402 19796 61516
rect 19068 61346 19124 61358
rect 19068 61294 19070 61346
rect 19122 61294 19124 61346
rect 19068 60226 19124 61294
rect 19068 60174 19070 60226
rect 19122 60174 19124 60226
rect 19068 60162 19124 60174
rect 19404 61348 19460 61358
rect 19740 61350 19742 61402
rect 19794 61350 19796 61402
rect 19740 61338 19796 61350
rect 20076 61348 20132 62132
rect 20188 61908 20244 62414
rect 20188 61842 20244 61852
rect 20188 61572 20244 61582
rect 20188 61478 20244 61516
rect 20076 61292 20244 61348
rect 19404 60788 19460 61292
rect 19628 61236 19684 61246
rect 19292 60004 19348 60014
rect 19404 60004 19460 60732
rect 19516 60900 19572 60910
rect 19516 60786 19572 60844
rect 19516 60734 19518 60786
rect 19570 60734 19572 60786
rect 19516 60722 19572 60734
rect 19628 60676 19684 61180
rect 19836 61180 20100 61190
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 19836 61114 20100 61124
rect 20076 60676 20132 60686
rect 19628 60620 19908 60676
rect 19740 60226 19796 60238
rect 19740 60174 19742 60226
rect 19794 60174 19796 60226
rect 19628 60004 19684 60014
rect 19404 60002 19684 60004
rect 19404 59950 19630 60002
rect 19682 59950 19684 60002
rect 19404 59948 19684 59950
rect 19740 60004 19796 60174
rect 19852 60226 19908 60620
rect 20076 60582 20132 60620
rect 19852 60174 19854 60226
rect 19906 60174 19908 60226
rect 19852 60162 19908 60174
rect 19964 60564 20020 60574
rect 19964 60004 20020 60508
rect 20188 60452 20244 61292
rect 20300 60788 20356 62860
rect 20412 62850 20468 62860
rect 20412 62132 20468 62142
rect 20412 61570 20468 62076
rect 20412 61518 20414 61570
rect 20466 61518 20468 61570
rect 20412 61506 20468 61518
rect 20748 61460 20804 61470
rect 20748 61366 20804 61404
rect 20412 61346 20468 61358
rect 20412 61294 20414 61346
rect 20466 61294 20468 61346
rect 20412 61012 20468 61294
rect 21084 61012 21140 66780
rect 21196 66770 21252 66780
rect 22988 65492 23044 67006
rect 23548 67060 23604 67790
rect 24668 67842 24724 68460
rect 25116 68180 25172 69020
rect 25228 68852 25284 68862
rect 25228 68738 25284 68796
rect 25228 68686 25230 68738
rect 25282 68686 25284 68738
rect 25228 68180 25284 68686
rect 25452 68628 25508 68638
rect 25564 68628 25620 69356
rect 25788 69298 25844 69310
rect 25788 69246 25790 69298
rect 25842 69246 25844 69298
rect 25788 68740 25844 69246
rect 25900 69298 25956 69310
rect 25900 69246 25902 69298
rect 25954 69246 25956 69298
rect 25900 68852 25956 69246
rect 26348 69186 26404 69198
rect 26348 69134 26350 69186
rect 26402 69134 26404 69186
rect 26124 68852 26180 68862
rect 25900 68796 26124 68852
rect 25788 68646 25844 68684
rect 25452 68626 25620 68628
rect 25452 68574 25454 68626
rect 25506 68574 25620 68626
rect 25452 68572 25620 68574
rect 25452 68516 25508 68572
rect 25452 68450 25508 68460
rect 25676 68514 25732 68526
rect 25676 68462 25678 68514
rect 25730 68462 25732 68514
rect 25676 68404 25732 68462
rect 26124 68514 26180 68796
rect 26124 68462 26126 68514
rect 26178 68462 26180 68514
rect 26124 68450 26180 68462
rect 25676 68348 26068 68404
rect 25788 68180 25844 68190
rect 25228 68124 25620 68180
rect 25116 68114 25172 68124
rect 24668 67790 24670 67842
rect 24722 67790 24724 67842
rect 23884 67732 23940 67742
rect 23884 67638 23940 67676
rect 24220 67730 24276 67742
rect 24220 67678 24222 67730
rect 24274 67678 24276 67730
rect 24220 67228 24276 67678
rect 24668 67732 24724 67790
rect 24668 67666 24724 67676
rect 25452 67956 25508 67966
rect 24220 67172 24388 67228
rect 23548 66994 23604 67004
rect 24332 65602 24388 67172
rect 25452 67170 25508 67900
rect 25452 67118 25454 67170
rect 25506 67118 25508 67170
rect 25452 67106 25508 67118
rect 25564 67170 25620 68124
rect 25788 67842 25844 68124
rect 25788 67790 25790 67842
rect 25842 67790 25844 67842
rect 25788 67228 25844 67790
rect 26012 67228 26068 68348
rect 25788 67172 25956 67228
rect 26012 67172 26180 67228
rect 25564 67118 25566 67170
rect 25618 67118 25620 67170
rect 25564 67106 25620 67118
rect 25228 67060 25284 67070
rect 25228 66966 25284 67004
rect 25676 67060 25732 67070
rect 24332 65550 24334 65602
rect 24386 65550 24388 65602
rect 24332 65538 24388 65550
rect 22988 65426 23044 65436
rect 23884 65492 23940 65502
rect 23884 65398 23940 65436
rect 24444 65490 24500 65502
rect 24444 65438 24446 65490
rect 24498 65438 24500 65490
rect 24444 64484 24500 65438
rect 24668 65492 24724 65502
rect 24668 65398 24724 65436
rect 25340 65492 25396 65502
rect 25340 65380 25396 65436
rect 25340 65378 25508 65380
rect 25340 65326 25342 65378
rect 25394 65326 25508 65378
rect 25340 65324 25508 65326
rect 25340 65314 25396 65324
rect 24444 64418 24500 64428
rect 25340 64484 25396 64494
rect 24332 63924 24388 63934
rect 24332 63830 24388 63868
rect 21420 63812 21476 63822
rect 21420 63140 21476 63756
rect 23548 63810 23604 63822
rect 23548 63758 23550 63810
rect 23602 63758 23604 63810
rect 21420 63074 21476 63084
rect 21532 63252 21588 63262
rect 21532 62466 21588 63196
rect 22764 63140 22820 63150
rect 22764 63046 22820 63084
rect 23324 63138 23380 63150
rect 23324 63086 23326 63138
rect 23378 63086 23380 63138
rect 21532 62414 21534 62466
rect 21586 62414 21588 62466
rect 21532 62402 21588 62414
rect 22092 62468 22148 62478
rect 22092 62242 22148 62412
rect 23324 62468 23380 63086
rect 23548 63028 23604 63758
rect 25228 63700 25284 63710
rect 24668 63698 25284 63700
rect 24668 63646 25230 63698
rect 25282 63646 25284 63698
rect 24668 63644 25284 63646
rect 24332 63140 24388 63150
rect 23660 63028 23716 63038
rect 23548 63026 23716 63028
rect 23548 62974 23662 63026
rect 23714 62974 23716 63026
rect 23548 62972 23716 62974
rect 23660 62962 23716 62972
rect 23996 63028 24052 63038
rect 24220 63028 24276 63038
rect 23996 63026 24276 63028
rect 23996 62974 23998 63026
rect 24050 62974 24222 63026
rect 24274 62974 24276 63026
rect 23996 62972 24276 62974
rect 23996 62962 24052 62972
rect 24220 62962 24276 62972
rect 23324 62402 23380 62412
rect 23884 62916 23940 62926
rect 22092 62190 22094 62242
rect 22146 62190 22148 62242
rect 22092 62178 22148 62190
rect 23884 61682 23940 62860
rect 24332 62578 24388 63084
rect 24668 63138 24724 63644
rect 25228 63634 25284 63644
rect 25340 63476 25396 64428
rect 25116 63420 25396 63476
rect 25452 64036 25508 65324
rect 25676 64708 25732 67004
rect 25788 67058 25844 67070
rect 25788 67006 25790 67058
rect 25842 67006 25844 67058
rect 25788 66948 25844 67006
rect 25788 66882 25844 66892
rect 24668 63086 24670 63138
rect 24722 63086 24724 63138
rect 24668 63074 24724 63086
rect 24892 63140 24948 63150
rect 24332 62526 24334 62578
rect 24386 62526 24388 62578
rect 24332 62514 24388 62526
rect 24668 62916 24724 62926
rect 24556 62468 24612 62478
rect 24556 62374 24612 62412
rect 24668 62466 24724 62860
rect 24668 62414 24670 62466
rect 24722 62414 24724 62466
rect 24668 62402 24724 62414
rect 24220 62356 24276 62366
rect 24220 62262 24276 62300
rect 23884 61630 23886 61682
rect 23938 61630 23940 61682
rect 23884 61618 23940 61630
rect 23996 61572 24052 61582
rect 24668 61572 24724 61582
rect 23996 61570 24724 61572
rect 23996 61518 23998 61570
rect 24050 61518 24670 61570
rect 24722 61518 24724 61570
rect 23996 61516 24724 61518
rect 23996 61506 24052 61516
rect 24668 61506 24724 61516
rect 24892 61570 24948 63084
rect 24892 61518 24894 61570
rect 24946 61518 24948 61570
rect 24892 61506 24948 61518
rect 25004 63028 25060 63038
rect 25116 63028 25172 63420
rect 25004 63026 25172 63028
rect 25004 62974 25006 63026
rect 25058 62974 25172 63026
rect 25004 62972 25172 62974
rect 25228 63138 25284 63150
rect 25228 63086 25230 63138
rect 25282 63086 25284 63138
rect 23324 61460 23380 61470
rect 23324 61366 23380 61404
rect 23212 61348 23268 61358
rect 23212 61254 23268 61292
rect 24444 61348 24500 61358
rect 24444 61254 24500 61292
rect 24780 61346 24836 61358
rect 24780 61294 24782 61346
rect 24834 61294 24836 61346
rect 20412 60956 20916 61012
rect 20636 60788 20692 60798
rect 20300 60786 20692 60788
rect 20300 60734 20638 60786
rect 20690 60734 20692 60786
rect 20300 60732 20692 60734
rect 19740 59948 20020 60004
rect 20076 60396 20244 60452
rect 19292 59910 19348 59948
rect 19628 59938 19684 59948
rect 20076 59780 20132 60396
rect 18844 59390 18846 59442
rect 18898 59390 18900 59442
rect 18844 59378 18900 59390
rect 19628 59724 20132 59780
rect 18508 59220 18564 59230
rect 18508 59126 18564 59164
rect 18172 58494 18174 58546
rect 18226 58494 18228 58546
rect 18172 58482 18228 58494
rect 17836 58436 17892 58446
rect 17836 58342 17892 58380
rect 17276 56914 17332 56924
rect 17388 57932 17668 57988
rect 18396 58322 18452 58334
rect 18396 58270 18398 58322
rect 18450 58270 18452 58322
rect 17164 56644 17220 56654
rect 17164 56550 17220 56588
rect 17388 56642 17444 57932
rect 17612 57762 17668 57774
rect 17612 57710 17614 57762
rect 17666 57710 17668 57762
rect 17612 57428 17668 57710
rect 17724 57652 17780 57662
rect 17724 57558 17780 57596
rect 17388 56590 17390 56642
rect 17442 56590 17444 56642
rect 16660 55804 16884 55860
rect 15260 53218 15316 53228
rect 15148 52994 15204 53004
rect 15260 53060 15316 53070
rect 15596 53060 15652 55244
rect 16604 54626 16660 55804
rect 17276 55410 17332 55422
rect 17276 55358 17278 55410
rect 17330 55358 17332 55410
rect 17164 55188 17220 55198
rect 17164 55094 17220 55132
rect 16604 54574 16606 54626
rect 16658 54574 16660 54626
rect 16604 54562 16660 54574
rect 16044 54290 16100 54302
rect 16044 54238 16046 54290
rect 16098 54238 16100 54290
rect 15260 53058 15652 53060
rect 15260 53006 15262 53058
rect 15314 53006 15652 53058
rect 15260 53004 15652 53006
rect 15260 52994 15316 53004
rect 12236 51874 12292 51884
rect 12348 52386 12516 52388
rect 12348 52334 12462 52386
rect 12514 52334 12516 52386
rect 12348 52332 12516 52334
rect 11788 51378 12068 51380
rect 11788 51326 11790 51378
rect 11842 51326 12068 51378
rect 11788 51324 12068 51326
rect 11788 51314 11844 51324
rect 11676 50706 11732 50718
rect 11676 50654 11678 50706
rect 11730 50654 11732 50706
rect 11676 50596 11732 50654
rect 11676 50530 11732 50540
rect 11564 50372 11732 50428
rect 11676 50370 11732 50372
rect 11676 50318 11678 50370
rect 11730 50318 11732 50370
rect 11564 49812 11620 49822
rect 11676 49812 11732 50318
rect 11564 49810 11732 49812
rect 11564 49758 11566 49810
rect 11618 49758 11732 49810
rect 11564 49756 11732 49758
rect 11900 49810 11956 51324
rect 12348 50818 12404 52332
rect 12460 52322 12516 52332
rect 14812 52946 14868 52958
rect 14812 52894 14814 52946
rect 14866 52894 14868 52946
rect 12684 52050 12740 52062
rect 12684 51998 12686 52050
rect 12738 51998 12740 52050
rect 12460 51938 12516 51950
rect 12460 51886 12462 51938
rect 12514 51886 12516 51938
rect 12460 51490 12516 51886
rect 12460 51438 12462 51490
rect 12514 51438 12516 51490
rect 12460 51426 12516 51438
rect 12348 50766 12350 50818
rect 12402 50766 12404 50818
rect 12348 50754 12404 50766
rect 12124 50596 12180 50606
rect 12124 50502 12180 50540
rect 12684 50594 12740 51998
rect 12908 52052 12964 52062
rect 12908 51958 12964 51996
rect 14812 51492 14868 52894
rect 15036 52948 15092 52958
rect 15036 52854 15092 52892
rect 15372 52724 15428 52734
rect 15596 52724 15652 53004
rect 15372 52722 15540 52724
rect 15372 52670 15374 52722
rect 15426 52670 15540 52722
rect 15372 52668 15540 52670
rect 15372 52658 15428 52668
rect 15484 52162 15540 52668
rect 15596 52658 15652 52668
rect 15932 53506 15988 53518
rect 15932 53454 15934 53506
rect 15986 53454 15988 53506
rect 15484 52110 15486 52162
rect 15538 52110 15540 52162
rect 15484 52098 15540 52110
rect 15708 52274 15764 52286
rect 15708 52222 15710 52274
rect 15762 52222 15764 52274
rect 15596 52052 15652 52062
rect 15596 51602 15652 51996
rect 15596 51550 15598 51602
rect 15650 51550 15652 51602
rect 15596 51538 15652 51550
rect 14812 51426 14868 51436
rect 15708 51378 15764 52222
rect 15932 51604 15988 53454
rect 16044 53172 16100 54238
rect 16940 53730 16996 53742
rect 16940 53678 16942 53730
rect 16994 53678 16996 53730
rect 16044 53106 16100 53116
rect 16380 53620 16436 53630
rect 16380 52948 16436 53564
rect 16940 53620 16996 53678
rect 16940 53554 16996 53564
rect 16380 52882 16436 52892
rect 16492 53508 16548 53518
rect 17276 53508 17332 55358
rect 17388 55300 17444 56590
rect 17500 56978 17556 56990
rect 17500 56926 17502 56978
rect 17554 56926 17556 56978
rect 17500 56308 17556 56926
rect 17612 56866 17668 57372
rect 18396 57092 18452 58270
rect 18956 58212 19012 58222
rect 18620 57540 18676 57550
rect 18956 57540 19012 58156
rect 18620 57538 19012 57540
rect 18620 57486 18622 57538
rect 18674 57486 19012 57538
rect 18620 57484 19012 57486
rect 18620 57428 18676 57484
rect 18620 57362 18676 57372
rect 18396 57026 18452 57036
rect 18060 56980 18116 56990
rect 18060 56886 18116 56924
rect 17612 56814 17614 56866
rect 17666 56814 17668 56866
rect 17612 56802 17668 56814
rect 17612 56308 17668 56318
rect 17500 56306 17668 56308
rect 17500 56254 17614 56306
rect 17666 56254 17668 56306
rect 17500 56252 17668 56254
rect 17612 56242 17668 56252
rect 18732 56196 18788 56206
rect 17500 56084 17556 56094
rect 17556 56028 17668 56084
rect 17500 55990 17556 56028
rect 17388 55234 17444 55244
rect 17612 54514 17668 56028
rect 17836 56082 17892 56094
rect 17836 56030 17838 56082
rect 17890 56030 17892 56082
rect 17724 55970 17780 55982
rect 17724 55918 17726 55970
rect 17778 55918 17780 55970
rect 17724 55412 17780 55918
rect 17836 55860 17892 56030
rect 17836 55794 17892 55804
rect 18060 56082 18116 56094
rect 18060 56030 18062 56082
rect 18114 56030 18116 56082
rect 17724 55346 17780 55356
rect 18060 55188 18116 56030
rect 18396 56082 18452 56094
rect 18396 56030 18398 56082
rect 18450 56030 18452 56082
rect 18396 55860 18452 56030
rect 18396 55794 18452 55804
rect 18396 55298 18452 55310
rect 18396 55246 18398 55298
rect 18450 55246 18452 55298
rect 18172 55188 18228 55198
rect 18060 55186 18228 55188
rect 18060 55134 18174 55186
rect 18226 55134 18228 55186
rect 18060 55132 18228 55134
rect 17612 54462 17614 54514
rect 17666 54462 17668 54514
rect 17388 53732 17444 53742
rect 17612 53732 17668 54462
rect 17388 53730 17668 53732
rect 17388 53678 17390 53730
rect 17442 53678 17668 53730
rect 17388 53676 17668 53678
rect 17724 54628 17780 54638
rect 17724 54402 17780 54572
rect 17724 54350 17726 54402
rect 17778 54350 17780 54402
rect 17388 53666 17444 53676
rect 17724 53620 17780 54350
rect 18172 54402 18228 55132
rect 18172 54350 18174 54402
rect 18226 54350 18228 54402
rect 18172 53732 18228 54350
rect 18172 53666 18228 53676
rect 18284 54516 18340 54526
rect 17836 53620 17892 53630
rect 17724 53618 17892 53620
rect 17724 53566 17838 53618
rect 17890 53566 17892 53618
rect 17724 53564 17892 53566
rect 17836 53554 17892 53564
rect 18172 53508 18228 53518
rect 17276 53452 17556 53508
rect 16268 52836 16324 52846
rect 16268 52742 16324 52780
rect 16492 51940 16548 53452
rect 17500 53170 17556 53452
rect 17500 53118 17502 53170
rect 17554 53118 17556 53170
rect 17500 53106 17556 53118
rect 17724 53170 17780 53182
rect 17724 53118 17726 53170
rect 17778 53118 17780 53170
rect 16604 53060 16660 53070
rect 16604 52946 16660 53004
rect 16604 52894 16606 52946
rect 16658 52894 16660 52946
rect 16604 52882 16660 52894
rect 17388 52948 17444 52958
rect 17388 52854 17444 52892
rect 16716 52274 16772 52286
rect 16716 52222 16718 52274
rect 16770 52222 16772 52274
rect 16716 52164 16772 52222
rect 16716 52098 16772 52108
rect 16492 51874 16548 51884
rect 16716 51940 16772 51950
rect 16044 51604 16100 51614
rect 15932 51602 16100 51604
rect 15932 51550 16046 51602
rect 16098 51550 16100 51602
rect 15932 51548 16100 51550
rect 15708 51326 15710 51378
rect 15762 51326 15764 51378
rect 14588 51268 14644 51278
rect 14588 51174 14644 51212
rect 15708 51268 15764 51326
rect 12684 50542 12686 50594
rect 12738 50542 12740 50594
rect 12684 50484 12740 50542
rect 12684 50418 12740 50428
rect 12908 50484 12964 50522
rect 12908 50418 12964 50428
rect 15148 50484 15204 50522
rect 12796 50370 12852 50382
rect 12796 50318 12798 50370
rect 12850 50318 12852 50370
rect 12684 49924 12740 49934
rect 12796 49924 12852 50318
rect 12684 49922 12852 49924
rect 12684 49870 12686 49922
rect 12738 49870 12852 49922
rect 12684 49868 12852 49870
rect 14812 50260 14868 50270
rect 12684 49858 12740 49868
rect 11900 49758 11902 49810
rect 11954 49758 11956 49810
rect 11564 49746 11620 49756
rect 11900 49746 11956 49758
rect 14812 49698 14868 50204
rect 15148 50036 15204 50428
rect 15260 50482 15316 50494
rect 15260 50430 15262 50482
rect 15314 50430 15316 50482
rect 15260 50260 15316 50430
rect 15708 50484 15764 51212
rect 15708 50418 15764 50428
rect 15820 50594 15876 50606
rect 15820 50542 15822 50594
rect 15874 50542 15876 50594
rect 15260 50194 15316 50204
rect 15148 49980 15428 50036
rect 15372 49924 15428 49980
rect 15596 50034 15652 50046
rect 15596 49982 15598 50034
rect 15650 49982 15652 50034
rect 15372 49922 15540 49924
rect 15372 49870 15374 49922
rect 15426 49870 15540 49922
rect 15372 49868 15540 49870
rect 15372 49858 15428 49868
rect 14812 49646 14814 49698
rect 14866 49646 14868 49698
rect 14812 49364 14868 49646
rect 14812 49298 14868 49308
rect 15484 49026 15540 49868
rect 15484 48974 15486 49026
rect 15538 48974 15540 49026
rect 15484 48962 15540 48974
rect 15596 48468 15652 49982
rect 15708 50036 15764 50046
rect 15820 50036 15876 50542
rect 15764 49980 15876 50036
rect 15708 49970 15764 49980
rect 15932 49924 15988 49934
rect 16044 49924 16100 51548
rect 16604 51492 16660 51502
rect 16716 51492 16772 51884
rect 17724 51716 17780 53118
rect 18172 52836 18228 53452
rect 18172 52162 18228 52780
rect 18172 52110 18174 52162
rect 18226 52110 18228 52162
rect 18172 52098 18228 52110
rect 17948 52050 18004 52062
rect 17948 51998 17950 52050
rect 18002 51998 18004 52050
rect 17948 51940 18004 51998
rect 18004 51884 18116 51940
rect 17948 51874 18004 51884
rect 16660 51436 16772 51492
rect 17164 51660 17780 51716
rect 17836 51828 17892 51838
rect 16604 51398 16660 51436
rect 15820 49922 16100 49924
rect 15820 49870 15934 49922
rect 15986 49870 16100 49922
rect 15820 49868 16100 49870
rect 16268 50596 16324 50606
rect 15708 49028 15764 49038
rect 15820 49028 15876 49868
rect 15932 49858 15988 49868
rect 16268 49812 16324 50540
rect 16380 50484 16436 50522
rect 16380 50418 16436 50428
rect 16044 49810 16324 49812
rect 16044 49758 16270 49810
rect 16322 49758 16324 49810
rect 16044 49756 16324 49758
rect 15708 49026 15876 49028
rect 15708 48974 15710 49026
rect 15762 48974 15876 49026
rect 15708 48972 15876 48974
rect 15932 49028 15988 49038
rect 16044 49028 16100 49756
rect 16268 49746 16324 49756
rect 15932 49026 16100 49028
rect 15932 48974 15934 49026
rect 15986 48974 16100 49026
rect 15932 48972 16100 48974
rect 15708 48962 15764 48972
rect 15932 48962 15988 48972
rect 15148 48412 15652 48468
rect 16268 48802 16324 48814
rect 16268 48750 16270 48802
rect 16322 48750 16324 48802
rect 11564 48244 11620 48254
rect 11452 48242 11620 48244
rect 11452 48190 11566 48242
rect 11618 48190 11620 48242
rect 11452 48188 11620 48190
rect 11564 48178 11620 48188
rect 11900 48244 11956 48254
rect 11900 48150 11956 48188
rect 11340 48018 11396 48030
rect 11340 47966 11342 48018
rect 11394 47966 11396 48018
rect 11340 47348 11396 47966
rect 11340 47282 11396 47292
rect 11340 46900 11396 46910
rect 11340 46806 11396 46844
rect 12908 46002 12964 46014
rect 12908 45950 12910 46002
rect 12962 45950 12964 46002
rect 12908 45668 12964 45950
rect 14924 46004 14980 46014
rect 14924 45910 14980 45948
rect 14252 45892 14308 45902
rect 14252 45778 14308 45836
rect 15036 45892 15092 45902
rect 14252 45726 14254 45778
rect 14306 45726 14308 45778
rect 13916 45668 13972 45678
rect 12908 45602 12964 45612
rect 13804 45612 13916 45668
rect 12572 45108 12628 45118
rect 12572 43650 12628 45052
rect 12908 44434 12964 44446
rect 12908 44382 12910 44434
rect 12962 44382 12964 44434
rect 12908 44324 12964 44382
rect 12908 43762 12964 44268
rect 13580 44324 13636 44334
rect 13580 44230 13636 44268
rect 13692 44212 13748 44222
rect 13804 44212 13860 45612
rect 13916 45574 13972 45612
rect 14028 45106 14084 45118
rect 14028 45054 14030 45106
rect 14082 45054 14084 45106
rect 14028 44324 14084 45054
rect 14252 44994 14308 45726
rect 14588 45778 14644 45790
rect 14588 45726 14590 45778
rect 14642 45726 14644 45778
rect 14588 45668 14644 45726
rect 14812 45668 14868 45678
rect 14588 45602 14644 45612
rect 14700 45666 14868 45668
rect 14700 45614 14814 45666
rect 14866 45614 14868 45666
rect 14700 45612 14868 45614
rect 14476 45108 14532 45118
rect 14700 45108 14756 45612
rect 14812 45602 14868 45612
rect 14812 45332 14868 45342
rect 14812 45238 14868 45276
rect 15036 45218 15092 45836
rect 15036 45166 15038 45218
rect 15090 45166 15092 45218
rect 15036 45154 15092 45166
rect 14532 45052 14756 45108
rect 14476 45014 14532 45052
rect 14252 44942 14254 44994
rect 14306 44942 14308 44994
rect 14252 44930 14308 44942
rect 13692 44210 13860 44212
rect 13692 44158 13694 44210
rect 13746 44158 13860 44210
rect 13692 44156 13860 44158
rect 13916 44212 13972 44222
rect 13692 44146 13748 44156
rect 12908 43710 12910 43762
rect 12962 43710 12964 43762
rect 12908 43698 12964 43710
rect 12572 43598 12574 43650
rect 12626 43598 12628 43650
rect 12572 43586 12628 43598
rect 13916 43538 13972 44156
rect 14028 43764 14084 44268
rect 15148 43708 15204 48412
rect 15484 48244 15540 48254
rect 15484 47348 15540 48188
rect 16268 48244 16324 48750
rect 16268 48178 16324 48188
rect 15484 46898 15540 47292
rect 15484 46846 15486 46898
rect 15538 46846 15540 46898
rect 15484 46834 15540 46846
rect 16604 48020 16660 48030
rect 15372 46562 15428 46574
rect 15372 46510 15374 46562
rect 15426 46510 15428 46562
rect 15372 45892 15428 46510
rect 15820 46562 15876 46574
rect 15820 46510 15822 46562
rect 15874 46510 15876 46562
rect 15820 46228 15876 46510
rect 15932 46452 15988 46462
rect 15932 46450 16100 46452
rect 15932 46398 15934 46450
rect 15986 46398 16100 46450
rect 15932 46396 16100 46398
rect 15932 46386 15988 46396
rect 15372 45798 15428 45836
rect 15484 46172 15876 46228
rect 15484 45220 15540 46172
rect 15820 46004 15876 46014
rect 15484 45154 15540 45164
rect 15596 46002 15876 46004
rect 15596 45950 15822 46002
rect 15874 45950 15876 46002
rect 15596 45948 15876 45950
rect 15596 44882 15652 45948
rect 15820 45938 15876 45948
rect 15932 45890 15988 45902
rect 15932 45838 15934 45890
rect 15986 45838 15988 45890
rect 15932 45108 15988 45838
rect 16044 45892 16100 46396
rect 16044 45836 16324 45892
rect 16044 45108 16100 45118
rect 15932 45106 16100 45108
rect 15932 45054 16046 45106
rect 16098 45054 16100 45106
rect 15932 45052 16100 45054
rect 15596 44830 15598 44882
rect 15650 44830 15652 44882
rect 15372 44100 15428 44110
rect 14028 43698 14084 43708
rect 13916 43486 13918 43538
rect 13970 43486 13972 43538
rect 13916 43474 13972 43486
rect 14700 43652 15204 43708
rect 15260 44044 15372 44100
rect 10892 42530 11284 42532
rect 10892 42478 11230 42530
rect 11282 42478 11284 42530
rect 10892 42476 11284 42478
rect 10556 42438 10612 42476
rect 10500 41244 10948 41300
rect 10444 41206 10500 41244
rect 10892 41186 10948 41244
rect 10892 41134 10894 41186
rect 10946 41134 10948 41186
rect 10892 41122 10948 41134
rect 11228 41188 11284 42476
rect 14028 43426 14084 43438
rect 14028 43374 14030 43426
rect 14082 43374 14084 43426
rect 11228 41094 11284 41132
rect 11564 41186 11620 41198
rect 11564 41134 11566 41186
rect 11618 41134 11620 41186
rect 9660 40462 9662 40514
rect 9714 40462 9716 40514
rect 9660 40450 9716 40462
rect 9772 40180 9828 40190
rect 9772 40086 9828 40124
rect 8540 39618 8708 39620
rect 8540 39566 8542 39618
rect 8594 39566 8708 39618
rect 8540 39564 8708 39566
rect 8540 39554 8596 39564
rect 1708 39506 1764 39518
rect 1708 39454 1710 39506
rect 1762 39454 1764 39506
rect 1708 39060 1764 39454
rect 6972 39508 7028 39518
rect 2044 39396 2100 39406
rect 2044 39302 2100 39340
rect 2492 39394 2548 39406
rect 2492 39342 2494 39394
rect 2546 39342 2548 39394
rect 1708 38994 1764 39004
rect 2492 39060 2548 39342
rect 2492 38994 2548 39004
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 6972 38162 7028 39452
rect 8204 39508 8260 39518
rect 8204 39414 8260 39452
rect 8092 39396 8148 39406
rect 7532 39060 7588 39070
rect 7532 38946 7588 39004
rect 7532 38894 7534 38946
rect 7586 38894 7588 38946
rect 7532 38882 7588 38894
rect 7644 38948 7700 38958
rect 7644 38854 7700 38892
rect 8092 38946 8148 39340
rect 8428 39394 8484 39406
rect 8428 39342 8430 39394
rect 8482 39342 8484 39394
rect 8428 39284 8484 39342
rect 8652 39396 8708 39564
rect 8764 39618 9268 39620
rect 8764 39566 8766 39618
rect 8818 39566 9214 39618
rect 9266 39566 9268 39618
rect 8764 39564 9268 39566
rect 8764 39554 8820 39564
rect 9212 39554 9268 39564
rect 9548 39620 9604 39630
rect 9324 39506 9380 39518
rect 9324 39454 9326 39506
rect 9378 39454 9380 39506
rect 9324 39396 9380 39454
rect 8652 39340 9380 39396
rect 9436 39394 9492 39406
rect 9436 39342 9438 39394
rect 9490 39342 9492 39394
rect 8428 39228 8596 39284
rect 8204 39172 8260 39182
rect 8204 39058 8260 39116
rect 8204 39006 8206 39058
rect 8258 39006 8260 39058
rect 8204 38994 8260 39006
rect 8092 38894 8094 38946
rect 8146 38894 8148 38946
rect 8092 38882 8148 38894
rect 6972 38110 6974 38162
rect 7026 38110 7028 38162
rect 6972 38098 7028 38110
rect 7868 38834 7924 38846
rect 7868 38782 7870 38834
rect 7922 38782 7924 38834
rect 7868 37492 7924 38782
rect 8428 38836 8484 38846
rect 8540 38836 8596 39228
rect 9436 39060 9492 39342
rect 9436 38994 9492 39004
rect 8764 38946 8820 38958
rect 8764 38894 8766 38946
rect 8818 38894 8820 38946
rect 8652 38836 8708 38846
rect 8540 38834 8708 38836
rect 8540 38782 8654 38834
rect 8706 38782 8708 38834
rect 8540 38780 8708 38782
rect 8428 38742 8484 38780
rect 8652 38770 8708 38780
rect 8764 38836 8820 38894
rect 9548 38946 9604 39564
rect 9772 39618 9828 39630
rect 9772 39566 9774 39618
rect 9826 39566 9828 39618
rect 9660 39172 9716 39182
rect 9660 39058 9716 39116
rect 9660 39006 9662 39058
rect 9714 39006 9716 39058
rect 9660 38994 9716 39006
rect 9772 39060 9828 39566
rect 10108 39618 10164 41020
rect 11340 40962 11396 40974
rect 11340 40910 11342 40962
rect 11394 40910 11396 40962
rect 10108 39566 10110 39618
rect 10162 39566 10164 39618
rect 10108 39554 10164 39566
rect 10332 40628 10388 40638
rect 9772 38994 9828 39004
rect 10332 39172 10388 40572
rect 11228 40180 11284 40190
rect 10780 39508 10836 39518
rect 10780 39506 11172 39508
rect 10780 39454 10782 39506
rect 10834 39454 11172 39506
rect 10780 39452 11172 39454
rect 10780 39442 10836 39452
rect 10332 39060 10388 39116
rect 10668 39060 10724 39070
rect 10332 39058 10724 39060
rect 10332 39006 10334 39058
rect 10386 39006 10670 39058
rect 10722 39006 10724 39058
rect 10332 39004 10724 39006
rect 10332 38994 10388 39004
rect 10668 38994 10724 39004
rect 10892 39060 10948 39070
rect 9548 38894 9550 38946
rect 9602 38894 9604 38946
rect 9548 38882 9604 38894
rect 9884 38948 9940 38958
rect 9884 38854 9940 38892
rect 8764 38770 8820 38780
rect 8988 38834 9044 38846
rect 8988 38782 8990 38834
rect 9042 38782 9044 38834
rect 8988 38164 9044 38782
rect 9100 38164 9156 38174
rect 8988 38162 9156 38164
rect 8988 38110 9102 38162
rect 9154 38110 9156 38162
rect 8988 38108 9156 38110
rect 9100 38098 9156 38108
rect 9884 38050 9940 38062
rect 9884 37998 9886 38050
rect 9938 37998 9940 38050
rect 9884 37828 9940 37998
rect 10332 37828 10388 37838
rect 9884 37826 10388 37828
rect 9884 37774 10334 37826
rect 10386 37774 10388 37826
rect 9884 37772 10388 37774
rect 7868 37426 7924 37436
rect 8764 37492 8820 37502
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 8764 36594 8820 37436
rect 8764 36542 8766 36594
rect 8818 36542 8820 36594
rect 8764 36530 8820 36542
rect 8092 36482 8148 36494
rect 8092 36430 8094 36482
rect 8146 36430 8148 36482
rect 8092 36260 8148 36430
rect 8092 36194 8148 36204
rect 10332 36260 10388 37772
rect 10892 36594 10948 39004
rect 11116 39058 11172 39452
rect 11116 39006 11118 39058
rect 11170 39006 11172 39058
rect 11116 38994 11172 39006
rect 11228 38948 11284 40124
rect 11340 39172 11396 40910
rect 11564 40516 11620 41134
rect 11900 41188 11956 41198
rect 11900 41094 11956 41132
rect 11564 40450 11620 40460
rect 12908 40516 12964 40526
rect 12908 39730 12964 40460
rect 13468 40516 13524 40526
rect 12908 39678 12910 39730
rect 12962 39678 12964 39730
rect 11340 39116 11508 39172
rect 11340 38948 11396 38958
rect 11228 38946 11396 38948
rect 11228 38894 11342 38946
rect 11394 38894 11396 38946
rect 11228 38892 11396 38894
rect 11340 38882 11396 38892
rect 11452 38946 11508 39116
rect 11452 38894 11454 38946
rect 11506 38894 11508 38946
rect 11452 38882 11508 38894
rect 12572 39060 12628 39070
rect 12572 38946 12628 39004
rect 12572 38894 12574 38946
rect 12626 38894 12628 38946
rect 12572 38882 12628 38894
rect 12684 38948 12740 38958
rect 12908 38948 12964 39678
rect 13244 40402 13300 40414
rect 13244 40350 13246 40402
rect 13298 40350 13300 40402
rect 13244 39060 13300 40350
rect 13468 40402 13524 40460
rect 13468 40350 13470 40402
rect 13522 40350 13524 40402
rect 13468 40338 13524 40350
rect 13692 40290 13748 40302
rect 13692 40238 13694 40290
rect 13746 40238 13748 40290
rect 13692 39508 13748 40238
rect 13692 39442 13748 39452
rect 14028 39284 14084 43374
rect 14140 43428 14196 43438
rect 14140 42978 14196 43372
rect 14140 42926 14142 42978
rect 14194 42926 14196 42978
rect 14140 42914 14196 42926
rect 14700 42644 14756 43652
rect 15148 42756 15204 42766
rect 15260 42756 15316 44044
rect 15372 44034 15428 44044
rect 15596 43428 15652 44830
rect 15708 44324 15764 44334
rect 15708 43764 15764 44268
rect 15708 43698 15764 43708
rect 16044 43540 16100 45052
rect 16156 44212 16212 44222
rect 16156 44118 16212 44156
rect 16156 43540 16212 43550
rect 16044 43484 16156 43540
rect 16268 43540 16324 45836
rect 16604 45778 16660 47964
rect 16940 46004 16996 46014
rect 16940 45910 16996 45948
rect 16604 45726 16606 45778
rect 16658 45726 16660 45778
rect 16604 45714 16660 45726
rect 17052 45666 17108 45678
rect 17052 45614 17054 45666
rect 17106 45614 17108 45666
rect 16604 45108 16660 45118
rect 16604 45014 16660 45052
rect 16716 44882 16772 44894
rect 16716 44830 16718 44882
rect 16770 44830 16772 44882
rect 16380 43540 16436 43550
rect 16268 43538 16436 43540
rect 16268 43486 16382 43538
rect 16434 43486 16436 43538
rect 16268 43484 16436 43486
rect 15596 43362 15652 43372
rect 15932 43428 15988 43438
rect 15932 43334 15988 43372
rect 16044 42756 16100 42766
rect 14700 42550 14756 42588
rect 14812 42754 15316 42756
rect 14812 42702 15150 42754
rect 15202 42702 15316 42754
rect 14812 42700 15316 42702
rect 15372 42754 16100 42756
rect 15372 42702 16046 42754
rect 16098 42702 16100 42754
rect 15372 42700 16100 42702
rect 14252 42196 14308 42206
rect 14140 41076 14196 41086
rect 14140 40982 14196 41020
rect 14252 40626 14308 42140
rect 14812 41970 14868 42700
rect 15148 42662 15204 42700
rect 15372 42642 15428 42700
rect 16044 42690 16100 42700
rect 15372 42590 15374 42642
rect 15426 42590 15428 42642
rect 15372 42578 15428 42590
rect 16044 42196 16100 42206
rect 16156 42196 16212 43484
rect 16380 43474 16436 43484
rect 16044 42194 16212 42196
rect 16044 42142 16046 42194
rect 16098 42142 16212 42194
rect 16044 42140 16212 42142
rect 16380 42644 16436 42654
rect 16044 42130 16100 42140
rect 14812 41918 14814 41970
rect 14866 41918 14868 41970
rect 14812 41906 14868 41918
rect 14252 40574 14254 40626
rect 14306 40574 14308 40626
rect 14252 40562 14308 40574
rect 14924 41746 14980 41758
rect 14924 41694 14926 41746
rect 14978 41694 14980 41746
rect 14924 39506 14980 41694
rect 14924 39454 14926 39506
rect 14978 39454 14980 39506
rect 14924 39442 14980 39454
rect 15708 40180 15764 40190
rect 15036 39396 15092 39406
rect 15036 39394 15204 39396
rect 15036 39342 15038 39394
rect 15090 39342 15204 39394
rect 15036 39340 15204 39342
rect 15036 39330 15092 39340
rect 14028 39218 14084 39228
rect 13244 38994 13300 39004
rect 13020 38948 13076 38958
rect 12908 38946 13076 38948
rect 12908 38894 13022 38946
rect 13074 38894 13076 38946
rect 12908 38892 13076 38894
rect 12684 38854 12740 38892
rect 13020 38882 13076 38892
rect 14028 38948 14084 38958
rect 14028 38854 14084 38892
rect 14700 38948 14756 38958
rect 13692 38724 13748 38734
rect 13692 38722 13860 38724
rect 13692 38670 13694 38722
rect 13746 38670 13860 38722
rect 13692 38668 13860 38670
rect 13692 38658 13748 38668
rect 13132 38610 13188 38622
rect 13132 38558 13134 38610
rect 13186 38558 13188 38610
rect 13132 38052 13188 38558
rect 13132 37986 13188 37996
rect 10892 36542 10894 36594
rect 10946 36542 10948 36594
rect 10892 36530 10948 36542
rect 10332 36194 10388 36204
rect 11340 36260 11396 36270
rect 11340 35700 11396 36204
rect 11564 35700 11620 35710
rect 11340 35698 11844 35700
rect 11340 35646 11566 35698
rect 11618 35646 11844 35698
rect 11340 35644 11844 35646
rect 11564 35634 11620 35644
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 11788 34130 11844 35644
rect 12236 35586 12292 35598
rect 12236 35534 12238 35586
rect 12290 35534 12292 35586
rect 12236 35140 12292 35534
rect 12236 35074 12292 35084
rect 13468 35140 13524 35150
rect 13468 35046 13524 35084
rect 13804 35028 13860 38668
rect 14028 38052 14084 38062
rect 14028 37958 14084 37996
rect 14700 37938 14756 38892
rect 15148 38836 15204 39340
rect 15708 38946 15764 40124
rect 16380 39618 16436 42588
rect 16604 42642 16660 42654
rect 16604 42590 16606 42642
rect 16658 42590 16660 42642
rect 16604 42196 16660 42590
rect 16604 42130 16660 42140
rect 16604 41970 16660 41982
rect 16604 41918 16606 41970
rect 16658 41918 16660 41970
rect 16604 41748 16660 41918
rect 16716 41860 16772 44830
rect 17052 44548 17108 45614
rect 17052 44482 17108 44492
rect 16716 41794 16772 41804
rect 16604 41682 16660 41692
rect 17164 40516 17220 51660
rect 17836 50932 17892 51772
rect 17612 50876 17892 50932
rect 17948 51490 18004 51502
rect 17948 51438 17950 51490
rect 18002 51438 18004 51490
rect 17612 50706 17668 50876
rect 17612 50654 17614 50706
rect 17666 50654 17668 50706
rect 17612 49810 17668 50654
rect 17724 50708 17780 50718
rect 17948 50708 18004 51438
rect 18060 51378 18116 51884
rect 18060 51326 18062 51378
rect 18114 51326 18116 51378
rect 18060 51314 18116 51326
rect 17724 50706 18004 50708
rect 17724 50654 17726 50706
rect 17778 50654 18004 50706
rect 17724 50652 18004 50654
rect 17724 50596 17780 50652
rect 17724 50530 17780 50540
rect 18284 50428 18340 54460
rect 18396 53508 18452 55246
rect 18732 54402 18788 56140
rect 18956 55970 19012 55982
rect 18956 55918 18958 55970
rect 19010 55918 19012 55970
rect 18844 54628 18900 54638
rect 18844 54534 18900 54572
rect 18956 54516 19012 55918
rect 18956 54450 19012 54460
rect 19068 55300 19124 55310
rect 18732 54350 18734 54402
rect 18786 54350 18788 54402
rect 18732 54338 18788 54350
rect 19068 53508 19124 55244
rect 19180 55186 19236 55198
rect 19180 55134 19182 55186
rect 19234 55134 19236 55186
rect 19180 53956 19236 55134
rect 19292 55188 19348 55198
rect 19292 55074 19348 55132
rect 19292 55022 19294 55074
rect 19346 55022 19348 55074
rect 19292 54404 19348 55022
rect 19628 54740 19684 59724
rect 19836 59612 20100 59622
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 19836 59546 20100 59556
rect 20636 58772 20692 60732
rect 20860 60786 20916 60956
rect 20860 60734 20862 60786
rect 20914 60734 20916 60786
rect 20860 60722 20916 60734
rect 21084 60786 21140 60956
rect 22204 61012 22260 61022
rect 22204 60918 22260 60956
rect 21084 60734 21086 60786
rect 21138 60734 21140 60786
rect 21084 60722 21140 60734
rect 22652 60676 22708 60686
rect 21980 60674 22708 60676
rect 21980 60622 22654 60674
rect 22706 60622 22708 60674
rect 21980 60620 22708 60622
rect 21308 60564 21364 60574
rect 21756 60564 21812 60574
rect 21308 60470 21364 60508
rect 21644 60562 21812 60564
rect 21644 60510 21758 60562
rect 21810 60510 21812 60562
rect 21644 60508 21812 60510
rect 20636 58716 21364 58772
rect 19836 58044 20100 58054
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 19836 57978 20100 57988
rect 19836 56476 20100 56486
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 19836 56410 20100 56420
rect 21084 55972 21140 55982
rect 21084 55970 21252 55972
rect 21084 55918 21086 55970
rect 21138 55918 21252 55970
rect 21084 55916 21252 55918
rect 21084 55906 21140 55916
rect 19836 54908 20100 54918
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 19836 54842 20100 54852
rect 19628 54684 19796 54740
rect 19292 54348 19684 54404
rect 19180 53900 19348 53956
rect 19180 53732 19236 53742
rect 19180 53638 19236 53676
rect 19292 53620 19348 53900
rect 19292 53554 19348 53564
rect 19404 53842 19460 53854
rect 19404 53790 19406 53842
rect 19458 53790 19460 53842
rect 19068 53452 19236 53508
rect 18396 53442 18452 53452
rect 18956 53284 19012 53294
rect 18732 53172 18788 53182
rect 18732 53058 18788 53116
rect 18732 53006 18734 53058
rect 18786 53006 18788 53058
rect 18508 52946 18564 52958
rect 18508 52894 18510 52946
rect 18562 52894 18564 52946
rect 17612 49758 17614 49810
rect 17666 49758 17668 49810
rect 17612 49746 17668 49758
rect 17724 50372 18340 50428
rect 18396 52274 18452 52286
rect 18396 52222 18398 52274
rect 18450 52222 18452 52274
rect 18396 50428 18452 52222
rect 18508 51940 18564 52894
rect 18620 52052 18676 52062
rect 18620 51958 18676 51996
rect 18508 51874 18564 51884
rect 18620 51266 18676 51278
rect 18620 51214 18622 51266
rect 18674 51214 18676 51266
rect 18508 50484 18564 50494
rect 18396 50372 18564 50428
rect 17500 48244 17556 48254
rect 17500 46676 17556 48188
rect 17612 47348 17668 47358
rect 17724 47348 17780 50372
rect 17836 50036 17892 50046
rect 17836 49026 17892 49980
rect 18396 50036 18452 50046
rect 18396 49810 18452 49980
rect 18396 49758 18398 49810
rect 18450 49758 18452 49810
rect 18396 49746 18452 49758
rect 18508 49698 18564 50372
rect 18508 49646 18510 49698
rect 18562 49646 18564 49698
rect 18508 49634 18564 49646
rect 18172 49364 18228 49374
rect 17836 48974 17838 49026
rect 17890 48974 17892 49026
rect 17836 48962 17892 48974
rect 18060 49138 18116 49150
rect 18060 49086 18062 49138
rect 18114 49086 18116 49138
rect 18060 49028 18116 49086
rect 18060 48962 18116 48972
rect 18172 48354 18228 49308
rect 18620 48692 18676 51214
rect 18396 48636 18676 48692
rect 18396 48468 18452 48636
rect 18396 48374 18452 48412
rect 18620 48468 18676 48478
rect 18732 48468 18788 53006
rect 18956 52836 19012 53228
rect 18956 52780 19124 52836
rect 19068 51378 19124 52780
rect 19180 51490 19236 53452
rect 19404 52946 19460 53790
rect 19516 53508 19572 53518
rect 19516 53414 19572 53452
rect 19404 52894 19406 52946
rect 19458 52894 19460 52946
rect 19404 52882 19460 52894
rect 19628 52948 19684 54348
rect 19740 53732 19796 54684
rect 20076 54516 20132 54526
rect 20076 54422 20132 54460
rect 19740 53666 19796 53676
rect 20748 54402 20804 54414
rect 20748 54350 20750 54402
rect 20802 54350 20804 54402
rect 19740 53508 19796 53518
rect 20748 53508 20804 54350
rect 19740 53506 20244 53508
rect 19740 53454 19742 53506
rect 19794 53454 20244 53506
rect 19740 53452 20244 53454
rect 19740 53442 19796 53452
rect 19836 53340 20100 53350
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 19836 53274 20100 53284
rect 20188 53172 20244 53452
rect 20748 53442 20804 53452
rect 20076 53116 20244 53172
rect 19740 52948 19796 52958
rect 19628 52946 19796 52948
rect 19628 52894 19742 52946
rect 19794 52894 19796 52946
rect 19628 52892 19796 52894
rect 19740 52882 19796 52892
rect 20076 52724 20132 53116
rect 20972 52948 21028 52958
rect 20972 52834 21028 52892
rect 20972 52782 20974 52834
rect 21026 52782 21028 52834
rect 20972 52770 21028 52782
rect 20076 52164 20132 52668
rect 20188 52164 20244 52174
rect 20076 52162 20244 52164
rect 20076 52110 20190 52162
rect 20242 52110 20244 52162
rect 20076 52108 20244 52110
rect 20188 52098 20244 52108
rect 20748 52164 20804 52174
rect 20748 51828 20804 52108
rect 19836 51772 20100 51782
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 19836 51706 20100 51716
rect 19180 51438 19182 51490
rect 19234 51438 19236 51490
rect 19180 51426 19236 51438
rect 19068 51326 19070 51378
rect 19122 51326 19124 51378
rect 19068 51314 19124 51326
rect 19740 50820 19796 50830
rect 19740 50706 19796 50764
rect 19740 50654 19742 50706
rect 19794 50654 19796 50706
rect 19740 50642 19796 50654
rect 20748 50594 20804 51772
rect 20748 50542 20750 50594
rect 20802 50542 20804 50594
rect 20748 50530 20804 50542
rect 21084 51492 21140 51502
rect 21084 50820 21140 51436
rect 18956 50484 19012 50494
rect 18956 49028 19012 50428
rect 20636 50484 20692 50522
rect 20636 50418 20692 50428
rect 19836 50204 20100 50214
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 19836 50138 20100 50148
rect 19068 49924 19124 49934
rect 19068 49922 19460 49924
rect 19068 49870 19070 49922
rect 19122 49870 19460 49922
rect 19068 49868 19460 49870
rect 19068 49858 19124 49868
rect 19180 49028 19236 49038
rect 18956 49026 19236 49028
rect 18956 48974 19182 49026
rect 19234 48974 19236 49026
rect 18956 48972 19236 48974
rect 19180 48962 19236 48972
rect 18620 48466 18788 48468
rect 18620 48414 18622 48466
rect 18674 48414 18788 48466
rect 18620 48412 18788 48414
rect 19068 48468 19124 48478
rect 18172 48302 18174 48354
rect 18226 48302 18228 48354
rect 18172 48290 18228 48302
rect 18508 48132 18564 48142
rect 18508 48038 18564 48076
rect 18284 47460 18340 47470
rect 18620 47460 18676 48412
rect 18732 48244 18788 48254
rect 18732 48150 18788 48188
rect 18060 47458 18340 47460
rect 18060 47406 18286 47458
rect 18338 47406 18340 47458
rect 18060 47404 18340 47406
rect 17612 47346 17780 47348
rect 17612 47294 17614 47346
rect 17666 47294 17780 47346
rect 17612 47292 17780 47294
rect 17612 47282 17668 47292
rect 17500 46674 17668 46676
rect 17500 46622 17502 46674
rect 17554 46622 17668 46674
rect 17500 46620 17668 46622
rect 17500 46610 17556 46620
rect 17500 46004 17556 46014
rect 17500 45106 17556 45948
rect 17500 45054 17502 45106
rect 17554 45054 17556 45106
rect 17500 45042 17556 45054
rect 17612 44884 17668 46620
rect 17724 45108 17780 47292
rect 17948 47348 18004 47358
rect 17948 47254 18004 47292
rect 17948 46676 18004 46686
rect 18060 46676 18116 47404
rect 18284 47394 18340 47404
rect 18396 47404 18676 47460
rect 18172 47236 18228 47246
rect 18172 47142 18228 47180
rect 17948 46674 18116 46676
rect 17948 46622 17950 46674
rect 18002 46622 18116 46674
rect 17948 46620 18116 46622
rect 17836 45332 17892 45342
rect 17948 45332 18004 46620
rect 18396 46340 18452 47404
rect 17836 45330 17948 45332
rect 17836 45278 17838 45330
rect 17890 45278 17948 45330
rect 17836 45276 17948 45278
rect 17836 45266 17892 45276
rect 17724 45042 17780 45052
rect 17612 44828 17892 44884
rect 17724 44324 17780 44334
rect 17276 44322 17780 44324
rect 17276 44270 17726 44322
rect 17778 44270 17780 44322
rect 17276 44268 17780 44270
rect 17276 44100 17332 44268
rect 17724 44258 17780 44268
rect 17724 44100 17780 44110
rect 17276 44006 17332 44044
rect 17612 44044 17724 44100
rect 17612 42642 17668 44044
rect 17724 44034 17780 44044
rect 17724 42756 17780 42766
rect 17836 42756 17892 44828
rect 17948 44210 18004 45276
rect 18284 46284 18452 46340
rect 18060 45218 18116 45230
rect 18060 45166 18062 45218
rect 18114 45166 18116 45218
rect 18060 45108 18116 45166
rect 18060 45042 18116 45052
rect 17948 44158 17950 44210
rect 18002 44158 18004 44210
rect 17948 44146 18004 44158
rect 18172 44882 18228 44894
rect 18172 44830 18174 44882
rect 18226 44830 18228 44882
rect 17724 42754 17892 42756
rect 17724 42702 17726 42754
rect 17778 42702 17892 42754
rect 17724 42700 17892 42702
rect 17724 42690 17780 42700
rect 17612 42590 17614 42642
rect 17666 42590 17668 42642
rect 17612 42578 17668 42590
rect 18172 42196 18228 44830
rect 18284 44210 18340 46284
rect 18620 45332 18676 45342
rect 18620 45238 18676 45276
rect 18396 45220 18452 45230
rect 18396 45126 18452 45164
rect 18844 45218 18900 45230
rect 18844 45166 18846 45218
rect 18898 45166 18900 45218
rect 18844 45108 18900 45166
rect 18844 45042 18900 45052
rect 18732 44994 18788 45006
rect 18732 44942 18734 44994
rect 18786 44942 18788 44994
rect 18508 44548 18564 44558
rect 18284 44158 18286 44210
rect 18338 44158 18340 44210
rect 18284 44100 18340 44158
rect 18284 44034 18340 44044
rect 18396 44324 18452 44334
rect 18284 43540 18340 43550
rect 18284 43446 18340 43484
rect 18396 42866 18452 44268
rect 18508 43314 18564 44492
rect 18732 44100 18788 44942
rect 18956 44212 19012 44222
rect 18620 43428 18676 43438
rect 18620 43334 18676 43372
rect 18508 43262 18510 43314
rect 18562 43262 18564 43314
rect 18508 43250 18564 43262
rect 18732 43204 18788 44044
rect 18396 42814 18398 42866
rect 18450 42814 18452 42866
rect 18396 42802 18452 42814
rect 18620 43148 18788 43204
rect 18844 44210 19012 44212
rect 18844 44158 18958 44210
rect 19010 44158 19012 44210
rect 18844 44156 19012 44158
rect 18172 42130 18228 42140
rect 18284 41972 18340 41982
rect 18172 41970 18340 41972
rect 18172 41918 18286 41970
rect 18338 41918 18340 41970
rect 18172 41916 18340 41918
rect 17500 41858 17556 41870
rect 17500 41806 17502 41858
rect 17554 41806 17556 41858
rect 17500 41748 17556 41806
rect 17500 41682 17556 41692
rect 17164 40450 17220 40460
rect 16380 39566 16382 39618
rect 16434 39566 16436 39618
rect 16380 39554 16436 39566
rect 15708 38894 15710 38946
rect 15762 38894 15764 38946
rect 15708 38882 15764 38894
rect 16044 39508 16100 39518
rect 15036 38834 15204 38836
rect 15036 38782 15150 38834
rect 15202 38782 15204 38834
rect 15036 38780 15204 38782
rect 14924 38164 14980 38174
rect 14924 38070 14980 38108
rect 15036 38050 15092 38780
rect 15148 38770 15204 38780
rect 15036 37998 15038 38050
rect 15090 37998 15092 38050
rect 15036 37986 15092 37998
rect 14700 37886 14702 37938
rect 14754 37886 14756 37938
rect 14700 37874 14756 37886
rect 16044 36370 16100 39452
rect 17388 39508 17444 39546
rect 17388 39442 17444 39452
rect 17388 39284 17444 39294
rect 16268 38836 16324 38846
rect 16268 37490 16324 38780
rect 17388 38834 17444 39228
rect 17388 38782 17390 38834
rect 17442 38782 17444 38834
rect 17388 38770 17444 38782
rect 17836 38948 17892 38958
rect 17836 38668 17892 38892
rect 17724 38612 17892 38668
rect 16268 37438 16270 37490
rect 16322 37438 16324 37490
rect 16268 37426 16324 37438
rect 16940 37938 16996 37950
rect 16940 37886 16942 37938
rect 16994 37886 16996 37938
rect 16044 36318 16046 36370
rect 16098 36318 16100 36370
rect 16044 36306 16100 36318
rect 16156 37154 16212 37166
rect 16156 37102 16158 37154
rect 16210 37102 16212 37154
rect 14588 36260 14644 36270
rect 14588 36258 14756 36260
rect 14588 36206 14590 36258
rect 14642 36206 14756 36258
rect 14588 36204 14756 36206
rect 14588 36194 14644 36204
rect 14364 35588 14420 35598
rect 14364 35494 14420 35532
rect 13804 34972 14084 35028
rect 13580 34804 13636 34814
rect 13580 34710 13636 34748
rect 11788 34078 11790 34130
rect 11842 34078 11844 34130
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 11788 33684 11844 34078
rect 4476 33674 4740 33684
rect 11676 33628 11844 33684
rect 12572 34018 12628 34030
rect 12572 33966 12574 34018
rect 12626 33966 12628 34018
rect 1708 33124 1764 33134
rect 1708 33030 1764 33068
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 11452 30996 11508 31006
rect 11676 30996 11732 33628
rect 12572 33572 12628 33966
rect 14028 33796 14084 34972
rect 14364 34916 14420 34926
rect 14364 34822 14420 34860
rect 14252 34804 14308 34814
rect 14252 34710 14308 34748
rect 12572 33506 12628 33516
rect 13804 33740 14084 33796
rect 14140 34692 14196 34702
rect 13692 33460 13748 33470
rect 13692 33366 13748 33404
rect 13804 33236 13860 33740
rect 13916 33572 13972 33582
rect 13916 33478 13972 33516
rect 14028 33460 14084 33470
rect 14028 33366 14084 33404
rect 14140 33348 14196 34636
rect 14700 34356 14756 36204
rect 14924 35810 14980 35822
rect 14924 35758 14926 35810
rect 14978 35758 14980 35810
rect 14924 35252 14980 35758
rect 15260 35812 15316 35822
rect 15260 35718 15316 35756
rect 16156 35812 16212 37102
rect 16380 36484 16436 36494
rect 16156 35746 16212 35756
rect 16268 36482 16436 36484
rect 16268 36430 16382 36482
rect 16434 36430 16436 36482
rect 16268 36428 16436 36430
rect 15820 35588 15876 35598
rect 15596 35532 15820 35588
rect 14924 35196 15316 35252
rect 15148 35028 15204 35038
rect 14812 35026 15204 35028
rect 14812 34974 15150 35026
rect 15202 34974 15204 35026
rect 14812 34972 15204 34974
rect 14812 34914 14868 34972
rect 15148 34962 15204 34972
rect 14812 34862 14814 34914
rect 14866 34862 14868 34914
rect 14812 34850 14868 34862
rect 15260 34916 15316 35196
rect 15596 34916 15652 35532
rect 15820 35494 15876 35532
rect 15316 34860 15428 34916
rect 15260 34850 15316 34860
rect 15036 34802 15092 34814
rect 15036 34750 15038 34802
rect 15090 34750 15092 34802
rect 15036 34692 15092 34750
rect 15036 34626 15092 34636
rect 15260 34692 15316 34702
rect 15148 34356 15204 34366
rect 15260 34356 15316 34636
rect 14700 34354 15316 34356
rect 14700 34302 15150 34354
rect 15202 34302 15316 34354
rect 14700 34300 15316 34302
rect 14700 34020 14756 34030
rect 14700 33926 14756 33964
rect 14476 33908 14532 33918
rect 14364 33852 14476 33908
rect 14364 33570 14420 33852
rect 14476 33842 14532 33852
rect 14364 33518 14366 33570
rect 14418 33518 14420 33570
rect 14140 33282 14196 33292
rect 14252 33346 14308 33358
rect 14252 33294 14254 33346
rect 14306 33294 14308 33346
rect 14252 33236 14308 33294
rect 13804 33180 14084 33236
rect 14028 32676 14084 33180
rect 14252 33170 14308 33180
rect 14364 32788 14420 33518
rect 14812 33348 14868 33358
rect 14812 33254 14868 33292
rect 14924 33236 14980 33246
rect 14924 33142 14980 33180
rect 14364 32732 14980 32788
rect 14028 32620 14756 32676
rect 14028 32564 14084 32620
rect 13916 32562 14084 32564
rect 13916 32510 14030 32562
rect 14082 32510 14084 32562
rect 13916 32508 14084 32510
rect 13916 32116 13972 32508
rect 14028 32498 14084 32508
rect 14700 32562 14756 32620
rect 14700 32510 14702 32562
rect 14754 32510 14756 32562
rect 14700 32498 14756 32510
rect 14364 32450 14420 32462
rect 14364 32398 14366 32450
rect 14418 32398 14420 32450
rect 14028 32338 14084 32350
rect 14028 32286 14030 32338
rect 14082 32286 14084 32338
rect 14028 32228 14084 32286
rect 14364 32340 14420 32398
rect 14812 32340 14868 32732
rect 14924 32562 14980 32732
rect 14924 32510 14926 32562
rect 14978 32510 14980 32562
rect 14924 32498 14980 32510
rect 14364 32284 14868 32340
rect 14028 32172 14756 32228
rect 13916 32060 14308 32116
rect 12124 31668 12180 31678
rect 12124 31106 12180 31612
rect 12124 31054 12126 31106
rect 12178 31054 12180 31106
rect 12124 31042 12180 31054
rect 11508 30940 11732 30996
rect 11452 30902 11508 30940
rect 14252 30882 14308 32060
rect 14700 32002 14756 32172
rect 14700 31950 14702 32002
rect 14754 31950 14756 32002
rect 14700 31938 14756 31950
rect 14924 32004 14980 32014
rect 14476 31780 14532 31790
rect 14476 31686 14532 31724
rect 14924 31778 14980 31948
rect 14924 31726 14926 31778
rect 14978 31726 14980 31778
rect 14924 31714 14980 31726
rect 14364 31668 14420 31678
rect 14364 31574 14420 31612
rect 14700 30996 14756 31006
rect 15036 30996 15092 34300
rect 15148 34290 15204 34300
rect 15372 34244 15428 34860
rect 15260 34188 15372 34244
rect 15260 34132 15316 34188
rect 15372 34150 15428 34188
rect 15484 34914 15652 34916
rect 15484 34862 15598 34914
rect 15650 34862 15652 34914
rect 15484 34860 15652 34862
rect 15148 34076 15316 34132
rect 15148 33346 15204 34076
rect 15148 33294 15150 33346
rect 15202 33294 15204 33346
rect 15148 33282 15204 33294
rect 15372 34020 15428 34030
rect 15372 33346 15428 33964
rect 15372 33294 15374 33346
rect 15426 33294 15428 33346
rect 15372 33282 15428 33294
rect 15484 33460 15540 34860
rect 15596 34850 15652 34860
rect 16268 34242 16324 36428
rect 16380 36418 16436 36428
rect 16380 34914 16436 34926
rect 16380 34862 16382 34914
rect 16434 34862 16436 34914
rect 16380 34692 16436 34862
rect 16380 34626 16436 34636
rect 16828 34916 16884 34926
rect 16268 34190 16270 34242
rect 16322 34190 16324 34242
rect 16044 34132 16100 34142
rect 16044 34038 16100 34076
rect 16268 34020 16324 34190
rect 16380 34244 16436 34254
rect 16380 34150 16436 34188
rect 16828 34132 16884 34860
rect 16940 34692 16996 37886
rect 17724 36370 17780 38612
rect 17948 38500 18004 38510
rect 17948 36594 18004 38444
rect 17948 36542 17950 36594
rect 18002 36542 18004 36594
rect 17948 36530 18004 36542
rect 18172 36372 18228 41916
rect 18284 41906 18340 41916
rect 18620 41970 18676 43148
rect 18620 41918 18622 41970
rect 18674 41918 18676 41970
rect 18620 41906 18676 41918
rect 18732 41972 18788 41982
rect 18732 41878 18788 41916
rect 18732 41748 18788 41758
rect 18732 40516 18788 41692
rect 18844 40852 18900 44156
rect 18956 44146 19012 44156
rect 18956 43316 19012 43326
rect 18956 41970 19012 43260
rect 18956 41918 18958 41970
rect 19010 41918 19012 41970
rect 18956 41906 19012 41918
rect 18844 40796 19012 40852
rect 18844 40626 18900 40638
rect 18844 40574 18846 40626
rect 18898 40574 18900 40626
rect 18844 40516 18900 40574
rect 18508 40460 18900 40516
rect 18508 39618 18564 40460
rect 18956 40404 19012 40796
rect 19068 40740 19124 48412
rect 19180 48132 19236 48142
rect 19236 48076 19348 48132
rect 19180 48066 19236 48076
rect 19180 46676 19236 46686
rect 19180 46582 19236 46620
rect 19292 46562 19348 48076
rect 19292 46510 19294 46562
rect 19346 46510 19348 46562
rect 19292 46498 19348 46510
rect 19404 44436 19460 49868
rect 21084 49922 21140 50764
rect 21196 50428 21252 55916
rect 21308 53730 21364 58716
rect 21532 57538 21588 57550
rect 21532 57486 21534 57538
rect 21586 57486 21588 57538
rect 21420 57092 21476 57102
rect 21420 56978 21476 57036
rect 21420 56926 21422 56978
rect 21474 56926 21476 56978
rect 21420 55970 21476 56926
rect 21532 56868 21588 57486
rect 21532 56802 21588 56812
rect 21420 55918 21422 55970
rect 21474 55918 21476 55970
rect 21420 55906 21476 55918
rect 21308 53678 21310 53730
rect 21362 53678 21364 53730
rect 21308 53666 21364 53678
rect 21420 53732 21476 53742
rect 21644 53732 21700 60508
rect 21756 60498 21812 60508
rect 21868 56868 21924 56878
rect 21868 56774 21924 56812
rect 21980 56644 22036 60620
rect 22652 60610 22708 60620
rect 24780 60452 24836 61294
rect 24780 60386 24836 60396
rect 24780 60004 24836 60014
rect 24780 59910 24836 59948
rect 24892 59892 24948 59902
rect 25004 59892 25060 62972
rect 25228 62580 25284 63086
rect 25452 62580 25508 63980
rect 25564 64652 25732 64708
rect 25788 65378 25844 65390
rect 25788 65326 25790 65378
rect 25842 65326 25844 65378
rect 25564 63810 25620 64652
rect 25676 64484 25732 64494
rect 25788 64484 25844 65326
rect 25732 64428 25844 64484
rect 25676 64390 25732 64428
rect 25564 63758 25566 63810
rect 25618 63758 25620 63810
rect 25564 62916 25620 63758
rect 25788 63922 25844 63934
rect 25788 63870 25790 63922
rect 25842 63870 25844 63922
rect 25788 63028 25844 63870
rect 25900 63924 25956 67172
rect 26124 66276 26180 67172
rect 26236 67060 26292 67070
rect 26236 66966 26292 67004
rect 26348 66836 26404 69134
rect 26684 68516 26740 68526
rect 26460 67730 26516 67742
rect 26460 67678 26462 67730
rect 26514 67678 26516 67730
rect 26460 67170 26516 67678
rect 26460 67118 26462 67170
rect 26514 67118 26516 67170
rect 26460 67106 26516 67118
rect 26460 66836 26516 66846
rect 26348 66780 26460 66836
rect 26460 66498 26516 66780
rect 26460 66446 26462 66498
rect 26514 66446 26516 66498
rect 26460 66434 26516 66446
rect 26572 66834 26628 66846
rect 26572 66782 26574 66834
rect 26626 66782 26628 66834
rect 26236 66276 26292 66286
rect 26124 66274 26292 66276
rect 26124 66222 26238 66274
rect 26290 66222 26292 66274
rect 26124 66220 26292 66222
rect 26236 66210 26292 66220
rect 26236 64036 26292 64046
rect 26236 63942 26292 63980
rect 25900 63858 25956 63868
rect 26012 63140 26068 63150
rect 26012 63046 26068 63084
rect 26236 63138 26292 63150
rect 26236 63086 26238 63138
rect 26290 63086 26292 63138
rect 26236 63028 26292 63086
rect 25788 62972 25956 63028
rect 25620 62860 25844 62916
rect 25564 62850 25620 62860
rect 25228 62524 25620 62580
rect 25452 62356 25508 62366
rect 25228 61570 25284 61582
rect 25228 61518 25230 61570
rect 25282 61518 25284 61570
rect 25228 61460 25284 61518
rect 25228 61394 25284 61404
rect 25340 60452 25396 60462
rect 25340 60002 25396 60396
rect 25340 59950 25342 60002
rect 25394 59950 25396 60002
rect 25340 59938 25396 59950
rect 24892 59890 25060 59892
rect 24892 59838 24894 59890
rect 24946 59838 25060 59890
rect 24892 59836 25060 59838
rect 25116 59890 25172 59902
rect 25116 59838 25118 59890
rect 25170 59838 25172 59890
rect 24444 59780 24500 59790
rect 24892 59780 24948 59836
rect 24332 59778 24948 59780
rect 24332 59726 24446 59778
rect 24498 59726 24948 59778
rect 24332 59724 24948 59726
rect 23660 58212 23716 58222
rect 23660 57762 23716 58156
rect 23660 57710 23662 57762
rect 23714 57710 23716 57762
rect 23660 57698 23716 57710
rect 23212 56980 23268 56990
rect 22652 56868 22708 56878
rect 22652 56774 22708 56812
rect 21868 56588 22036 56644
rect 22316 56754 22372 56766
rect 22316 56702 22318 56754
rect 22370 56702 22372 56754
rect 21756 56084 21812 56094
rect 21756 55990 21812 56028
rect 21756 53732 21812 53742
rect 21644 53676 21756 53732
rect 21308 53060 21364 53070
rect 21420 53060 21476 53676
rect 21756 53666 21812 53676
rect 21308 53058 21476 53060
rect 21308 53006 21310 53058
rect 21362 53006 21476 53058
rect 21308 53004 21476 53006
rect 21532 53618 21588 53630
rect 21532 53566 21534 53618
rect 21586 53566 21588 53618
rect 21532 53060 21588 53566
rect 21308 52994 21364 53004
rect 21532 52994 21588 53004
rect 21756 53506 21812 53518
rect 21756 53454 21758 53506
rect 21810 53454 21812 53506
rect 21756 51156 21812 53454
rect 21868 52946 21924 56588
rect 22204 55522 22260 55534
rect 22204 55470 22206 55522
rect 22258 55470 22260 55522
rect 21980 55412 22036 55422
rect 21980 55318 22036 55356
rect 22092 55300 22148 55310
rect 22092 55206 22148 55244
rect 21868 52894 21870 52946
rect 21922 52894 21924 52946
rect 21868 52882 21924 52894
rect 21980 53730 22036 53742
rect 21980 53678 21982 53730
rect 22034 53678 22036 53730
rect 21980 52948 22036 53678
rect 21980 52882 22036 52892
rect 22092 53508 22148 53518
rect 21868 52164 21924 52174
rect 21868 52070 21924 52108
rect 21756 51090 21812 51100
rect 21980 52050 22036 52062
rect 21980 51998 21982 52050
rect 22034 51998 22036 52050
rect 21196 50372 21364 50428
rect 21084 49870 21086 49922
rect 21138 49870 21140 49922
rect 21084 49858 21140 49870
rect 20412 49028 20468 49038
rect 20412 48934 20468 48972
rect 19964 48914 20020 48926
rect 19964 48862 19966 48914
rect 20018 48862 20020 48914
rect 19964 48804 20020 48862
rect 20860 48916 20916 48926
rect 19964 48748 20244 48804
rect 19836 48636 20100 48646
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 19836 48570 20100 48580
rect 19292 44380 19460 44436
rect 19516 47348 19572 47358
rect 19516 46450 19572 47292
rect 19836 47068 20100 47078
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 19836 47002 20100 47012
rect 20188 47012 20244 48748
rect 20300 48468 20356 48478
rect 20300 48242 20356 48412
rect 20860 48466 20916 48860
rect 20860 48414 20862 48466
rect 20914 48414 20916 48466
rect 20860 48402 20916 48414
rect 21196 48804 21252 48814
rect 21196 48354 21252 48748
rect 21196 48302 21198 48354
rect 21250 48302 21252 48354
rect 21196 48290 21252 48302
rect 20300 48190 20302 48242
rect 20354 48190 20356 48242
rect 20300 47236 20356 48190
rect 20524 48020 20580 48030
rect 20524 47926 20580 47964
rect 20748 47684 20804 47694
rect 20748 47590 20804 47628
rect 20412 47348 20468 47358
rect 20412 47254 20468 47292
rect 20300 47170 20356 47180
rect 20636 47234 20692 47246
rect 20636 47182 20638 47234
rect 20690 47182 20692 47234
rect 20636 47012 20692 47182
rect 20188 46956 20692 47012
rect 19516 46398 19518 46450
rect 19570 46398 19572 46450
rect 19180 44212 19236 44222
rect 19180 44118 19236 44156
rect 19180 41748 19236 41758
rect 19180 41186 19236 41692
rect 19292 41300 19348 44380
rect 19404 44210 19460 44222
rect 19404 44158 19406 44210
rect 19458 44158 19460 44210
rect 19404 44100 19460 44158
rect 19404 44034 19460 44044
rect 19516 42756 19572 46398
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 19964 45332 20020 45342
rect 19852 45108 19908 45118
rect 19852 45014 19908 45052
rect 19964 45106 20020 45276
rect 19964 45054 19966 45106
rect 20018 45054 20020 45106
rect 19964 44546 20020 45054
rect 20188 44884 20244 44894
rect 20188 44790 20244 44828
rect 20300 44882 20356 44894
rect 20300 44830 20302 44882
rect 20354 44830 20356 44882
rect 19964 44494 19966 44546
rect 20018 44494 20020 44546
rect 19964 44482 20020 44494
rect 19628 44210 19684 44222
rect 19628 44158 19630 44210
rect 19682 44158 19684 44210
rect 19628 43316 19684 44158
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 19852 43764 19908 43774
rect 19852 43538 19908 43708
rect 20300 43652 20356 44830
rect 20636 44324 20692 46956
rect 20860 44884 20916 44894
rect 20748 44548 20804 44558
rect 20748 44454 20804 44492
rect 20636 44268 20804 44324
rect 20300 43586 20356 43596
rect 20412 44210 20468 44222
rect 20412 44158 20414 44210
rect 20466 44158 20468 44210
rect 19852 43486 19854 43538
rect 19906 43486 19908 43538
rect 19852 43474 19908 43486
rect 19740 43426 19796 43438
rect 20412 43428 20468 44158
rect 19740 43374 19742 43426
rect 19794 43374 19796 43426
rect 19740 43316 19796 43374
rect 19684 43260 19796 43316
rect 20076 43372 20468 43428
rect 20636 44098 20692 44110
rect 20636 44046 20638 44098
rect 20690 44046 20692 44098
rect 19628 43250 19684 43260
rect 20076 43092 20132 43372
rect 20636 43092 20692 44046
rect 20076 43036 20244 43092
rect 20188 42978 20244 43036
rect 20188 42926 20190 42978
rect 20242 42926 20244 42978
rect 19964 42756 20020 42766
rect 19516 42754 20020 42756
rect 19516 42702 19966 42754
rect 20018 42702 20020 42754
rect 19516 42700 20020 42702
rect 19964 42690 20020 42700
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 19852 42196 19908 42206
rect 19628 41970 19684 41982
rect 19628 41918 19630 41970
rect 19682 41918 19684 41970
rect 19292 41244 19460 41300
rect 19180 41134 19182 41186
rect 19234 41134 19236 41186
rect 19180 41122 19236 41134
rect 19292 41076 19348 41086
rect 19068 40674 19124 40684
rect 19180 40964 19236 40974
rect 18844 40348 19012 40404
rect 18508 39566 18510 39618
rect 18562 39566 18564 39618
rect 18508 39554 18564 39566
rect 18620 40292 18676 40302
rect 18396 39060 18452 39070
rect 18396 38966 18452 39004
rect 18284 38836 18340 38846
rect 18284 38742 18340 38780
rect 18620 36484 18676 40236
rect 18844 39842 18900 40348
rect 19180 40180 19236 40908
rect 18844 39790 18846 39842
rect 18898 39790 18900 39842
rect 18844 39778 18900 39790
rect 18956 40124 19236 40180
rect 18844 38836 18900 38846
rect 18844 38742 18900 38780
rect 18956 36596 19012 40124
rect 19068 39730 19124 39742
rect 19068 39678 19070 39730
rect 19122 39678 19124 39730
rect 19068 38948 19124 39678
rect 19292 39506 19348 41020
rect 19404 40404 19460 41244
rect 19628 41076 19684 41918
rect 19852 41970 19908 42140
rect 19852 41918 19854 41970
rect 19906 41918 19908 41970
rect 19852 41186 19908 41918
rect 19852 41134 19854 41186
rect 19906 41134 19908 41186
rect 19852 41122 19908 41134
rect 19964 41970 20020 41982
rect 19964 41918 19966 41970
rect 20018 41918 20020 41970
rect 19964 41860 20020 41918
rect 19516 41074 19684 41076
rect 19516 41022 19630 41074
rect 19682 41022 19684 41074
rect 19516 41020 19684 41022
rect 19964 41076 20020 41804
rect 20076 41300 20132 41310
rect 20188 41300 20244 42926
rect 20412 43036 20692 43092
rect 20412 42978 20468 43036
rect 20748 42980 20804 44268
rect 20412 42926 20414 42978
rect 20466 42926 20468 42978
rect 20412 42194 20468 42926
rect 20412 42142 20414 42194
rect 20466 42142 20468 42194
rect 20412 42130 20468 42142
rect 20524 42924 20804 42980
rect 20076 41298 20244 41300
rect 20076 41246 20078 41298
rect 20130 41246 20244 41298
rect 20076 41244 20244 41246
rect 20076 41234 20132 41244
rect 20188 41076 20244 41086
rect 19964 41074 20244 41076
rect 19964 41022 20190 41074
rect 20242 41022 20244 41074
rect 19964 41020 20244 41022
rect 19516 40964 19572 41020
rect 19628 41010 19684 41020
rect 20188 41010 20244 41020
rect 19516 40898 19572 40908
rect 19836 40796 20100 40806
rect 19628 40740 19684 40750
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 19628 40628 19684 40684
rect 19852 40628 19908 40638
rect 19628 40626 19908 40628
rect 19628 40574 19854 40626
rect 19906 40574 19908 40626
rect 19628 40572 19908 40574
rect 19516 40404 19572 40414
rect 19404 40402 19796 40404
rect 19404 40350 19518 40402
rect 19570 40350 19796 40402
rect 19404 40348 19796 40350
rect 19516 40338 19572 40348
rect 19628 39956 19684 39966
rect 19516 39844 19572 39854
rect 19516 39618 19572 39788
rect 19628 39730 19684 39900
rect 19628 39678 19630 39730
rect 19682 39678 19684 39730
rect 19628 39666 19684 39678
rect 19516 39566 19518 39618
rect 19570 39566 19572 39618
rect 19516 39554 19572 39566
rect 19740 39620 19796 40348
rect 19852 39844 19908 40572
rect 20188 40628 20244 40638
rect 20188 40534 20244 40572
rect 19852 39778 19908 39788
rect 20076 40514 20132 40526
rect 20076 40462 20078 40514
rect 20130 40462 20132 40514
rect 20076 39844 20132 40462
rect 20412 40516 20468 40526
rect 20524 40516 20580 42924
rect 20860 42868 20916 44828
rect 20636 42812 20916 42868
rect 21196 43538 21252 43550
rect 21196 43486 21198 43538
rect 21250 43486 21252 43538
rect 21196 42868 21252 43486
rect 21308 43316 21364 50372
rect 21644 49812 21700 49822
rect 21644 49718 21700 49756
rect 21420 48916 21476 48926
rect 21420 48466 21476 48860
rect 21756 48804 21812 48814
rect 21756 48710 21812 48748
rect 21420 48414 21422 48466
rect 21474 48414 21476 48466
rect 21420 48402 21476 48414
rect 21532 48244 21588 48254
rect 21532 48150 21588 48188
rect 21644 48242 21700 48254
rect 21644 48190 21646 48242
rect 21698 48190 21700 48242
rect 21644 46116 21700 48190
rect 21868 48242 21924 48254
rect 21868 48190 21870 48242
rect 21922 48190 21924 48242
rect 21868 47124 21924 48190
rect 21868 47058 21924 47068
rect 21868 46900 21924 46910
rect 21980 46900 22036 51998
rect 22092 49810 22148 53452
rect 22204 53396 22260 55470
rect 22316 55076 22372 56702
rect 22764 56644 22820 56654
rect 23100 56644 23156 56654
rect 22764 56642 23156 56644
rect 22764 56590 22766 56642
rect 22818 56590 23102 56642
rect 23154 56590 23156 56642
rect 22764 56588 23156 56590
rect 22764 56084 22820 56588
rect 23100 56578 23156 56588
rect 22764 56018 22820 56028
rect 22316 55020 22596 55076
rect 22428 53730 22484 53742
rect 22428 53678 22430 53730
rect 22482 53678 22484 53730
rect 22204 53340 22372 53396
rect 22316 52946 22372 53340
rect 22316 52894 22318 52946
rect 22370 52894 22372 52946
rect 22204 52836 22260 52846
rect 22204 52742 22260 52780
rect 22316 52052 22372 52894
rect 22428 52052 22484 53678
rect 22540 53618 22596 55020
rect 22540 53566 22542 53618
rect 22594 53566 22596 53618
rect 22540 53554 22596 53566
rect 23100 53620 23156 53630
rect 22988 53060 23044 53070
rect 23100 53060 23156 53564
rect 22988 53058 23156 53060
rect 22988 53006 22990 53058
rect 23042 53006 23156 53058
rect 22988 53004 23156 53006
rect 22988 52994 23044 53004
rect 22428 51996 22820 52052
rect 22316 51986 22372 51996
rect 22428 51380 22484 51418
rect 22092 49758 22094 49810
rect 22146 49758 22148 49810
rect 22092 49746 22148 49758
rect 22316 51324 22428 51380
rect 22204 49698 22260 49710
rect 22204 49646 22206 49698
rect 22258 49646 22260 49698
rect 22204 48354 22260 49646
rect 22316 49026 22372 51324
rect 22428 51314 22484 51324
rect 22428 51156 22484 51166
rect 22428 49140 22484 51100
rect 22652 49924 22708 49934
rect 22652 49830 22708 49868
rect 22764 49812 22820 51996
rect 23100 51492 23156 51502
rect 23100 51398 23156 51436
rect 22988 51380 23044 51390
rect 22428 49084 22596 49140
rect 22316 48974 22318 49026
rect 22370 48974 22372 49026
rect 22316 48468 22372 48974
rect 22316 48412 22484 48468
rect 22204 48302 22206 48354
rect 22258 48302 22260 48354
rect 22204 48290 22260 48302
rect 22316 48244 22372 48254
rect 22316 48150 22372 48188
rect 22428 47236 22484 48412
rect 22540 48242 22596 49084
rect 22764 49138 22820 49756
rect 22764 49086 22766 49138
rect 22818 49086 22820 49138
rect 22764 49074 22820 49086
rect 22876 51378 23044 51380
rect 22876 51326 22990 51378
rect 23042 51326 23044 51378
rect 22876 51324 23044 51326
rect 22764 48914 22820 48926
rect 22764 48862 22766 48914
rect 22818 48862 22820 48914
rect 22764 48468 22820 48862
rect 22876 48916 22932 51324
rect 22988 51314 23044 51324
rect 22876 48850 22932 48860
rect 22988 50484 23044 50494
rect 23212 50484 23268 56924
rect 23660 56866 23716 56878
rect 23660 56814 23662 56866
rect 23714 56814 23716 56866
rect 23660 56532 23716 56814
rect 23660 56466 23716 56476
rect 23884 53732 23940 53742
rect 23772 53060 23828 53070
rect 23436 51938 23492 51950
rect 23436 51886 23438 51938
rect 23490 51886 23492 51938
rect 22988 50482 23268 50484
rect 22988 50430 22990 50482
rect 23042 50430 23268 50482
rect 22988 50428 23268 50430
rect 23324 51602 23380 51614
rect 23324 51550 23326 51602
rect 23378 51550 23380 51602
rect 22764 48402 22820 48412
rect 22540 48190 22542 48242
rect 22594 48190 22596 48242
rect 22540 48178 22596 48190
rect 22764 48242 22820 48254
rect 22764 48190 22766 48242
rect 22818 48190 22820 48242
rect 22764 47684 22820 48190
rect 22764 47618 22820 47628
rect 22428 47180 22820 47236
rect 21868 46898 22036 46900
rect 21868 46846 21870 46898
rect 21922 46846 22036 46898
rect 21868 46844 22036 46846
rect 22204 47012 22260 47022
rect 21868 46834 21924 46844
rect 21644 46022 21700 46060
rect 21756 46674 21812 46686
rect 21756 46622 21758 46674
rect 21810 46622 21812 46674
rect 21644 45892 21700 45902
rect 21532 45780 21588 45790
rect 21644 45780 21700 45836
rect 21532 45778 21700 45780
rect 21532 45726 21534 45778
rect 21586 45726 21700 45778
rect 21532 45724 21700 45726
rect 21532 45714 21588 45724
rect 21420 44548 21476 44558
rect 21476 44492 21588 44548
rect 21420 44482 21476 44492
rect 21420 43652 21476 43662
rect 21420 43558 21476 43596
rect 21532 43538 21588 44492
rect 21532 43486 21534 43538
rect 21586 43486 21588 43538
rect 21532 43474 21588 43486
rect 21644 44322 21700 45724
rect 21644 44270 21646 44322
rect 21698 44270 21700 44322
rect 21308 43260 21588 43316
rect 21196 42812 21476 42868
rect 20636 42754 20692 42812
rect 20636 42702 20638 42754
rect 20690 42702 20692 42754
rect 20636 41972 20692 42702
rect 20748 42644 20804 42654
rect 21308 42644 21364 42654
rect 20748 42642 21364 42644
rect 20748 42590 20750 42642
rect 20802 42590 21310 42642
rect 21362 42590 21364 42642
rect 20748 42588 21364 42590
rect 20748 42578 20804 42588
rect 21308 42578 21364 42588
rect 20636 41906 20692 41916
rect 21420 42530 21476 42812
rect 21420 42478 21422 42530
rect 21474 42478 21476 42530
rect 20636 41748 20692 41758
rect 20636 41300 20692 41692
rect 20636 41298 20804 41300
rect 20636 41246 20638 41298
rect 20690 41246 20804 41298
rect 20636 41244 20804 41246
rect 20636 41234 20692 41244
rect 20412 40514 20580 40516
rect 20412 40462 20414 40514
rect 20466 40462 20580 40514
rect 20412 40460 20580 40462
rect 20412 40450 20468 40460
rect 20636 40180 20692 40190
rect 20524 40178 20692 40180
rect 20524 40126 20638 40178
rect 20690 40126 20692 40178
rect 20524 40124 20692 40126
rect 20524 39844 20580 40124
rect 20636 40114 20692 40124
rect 20076 39778 20132 39788
rect 20188 39788 20580 39844
rect 20636 39844 20692 39854
rect 20188 39730 20244 39788
rect 20188 39678 20190 39730
rect 20242 39678 20244 39730
rect 20188 39666 20244 39678
rect 19964 39620 20020 39630
rect 19740 39618 20020 39620
rect 19740 39566 19966 39618
rect 20018 39566 20020 39618
rect 19740 39564 20020 39566
rect 19292 39454 19294 39506
rect 19346 39454 19348 39506
rect 19068 38854 19124 38892
rect 19180 39284 19236 39294
rect 19180 38946 19236 39228
rect 19180 38894 19182 38946
rect 19234 38894 19236 38946
rect 19180 38882 19236 38894
rect 19180 38500 19236 38510
rect 19292 38500 19348 39454
rect 19236 38444 19348 38500
rect 19404 39508 19460 39518
rect 19180 38434 19236 38444
rect 19404 37380 19460 39452
rect 19852 39508 19908 39564
rect 19964 39554 20020 39564
rect 20300 39620 20356 39630
rect 19852 39442 19908 39452
rect 19740 39396 19796 39434
rect 19740 39330 19796 39340
rect 19836 39228 20100 39238
rect 19628 39172 19684 39182
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 19628 38836 19684 39116
rect 19628 38742 19684 38780
rect 20300 38668 20356 39564
rect 20636 39508 20692 39788
rect 20636 39414 20692 39452
rect 20636 39060 20692 39070
rect 20412 38836 20468 38846
rect 20412 38742 20468 38780
rect 20636 38834 20692 39004
rect 20636 38782 20638 38834
rect 20690 38782 20692 38834
rect 20636 38770 20692 38782
rect 20188 38612 20356 38668
rect 20076 38164 20132 38174
rect 20076 38050 20132 38108
rect 20076 37998 20078 38050
rect 20130 37998 20132 38050
rect 20076 37986 20132 37998
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 19740 37380 19796 37390
rect 19404 37378 19796 37380
rect 19404 37326 19742 37378
rect 19794 37326 19796 37378
rect 19404 37324 19796 37326
rect 19740 37314 19796 37324
rect 19852 37380 19908 37390
rect 19852 37378 20132 37380
rect 19852 37326 19854 37378
rect 19906 37326 20132 37378
rect 19852 37324 20132 37326
rect 19852 37314 19908 37324
rect 20076 37268 20132 37324
rect 20188 37268 20244 38612
rect 20748 38164 20804 41244
rect 21308 40402 21364 40414
rect 21308 40350 21310 40402
rect 21362 40350 21364 40402
rect 20972 40292 21028 40302
rect 20972 40198 21028 40236
rect 21308 39956 21364 40350
rect 21420 40180 21476 42478
rect 21532 40964 21588 43260
rect 21644 42868 21700 44270
rect 21756 45444 21812 46622
rect 21980 46674 22036 46686
rect 21980 46622 21982 46674
rect 22034 46622 22036 46674
rect 21980 45892 22036 46622
rect 22092 46676 22148 46686
rect 22092 46582 22148 46620
rect 21980 45826 22036 45836
rect 22092 45890 22148 45902
rect 22092 45838 22094 45890
rect 22146 45838 22148 45890
rect 22092 45780 22148 45838
rect 22092 45444 22148 45724
rect 21756 45388 22148 45444
rect 21756 44436 21812 45388
rect 22092 45220 22148 45230
rect 21868 44436 21924 44446
rect 21756 44434 21924 44436
rect 21756 44382 21870 44434
rect 21922 44382 21924 44434
rect 21756 44380 21924 44382
rect 21756 44324 21812 44380
rect 21868 44370 21924 44380
rect 21756 44258 21812 44268
rect 21868 43652 21924 43662
rect 21868 43538 21924 43596
rect 21868 43486 21870 43538
rect 21922 43486 21924 43538
rect 21868 43474 21924 43486
rect 21644 42802 21700 42812
rect 21644 42532 21700 42542
rect 21644 42530 21812 42532
rect 21644 42478 21646 42530
rect 21698 42478 21812 42530
rect 21644 42476 21812 42478
rect 21644 42466 21700 42476
rect 21756 41860 21812 42476
rect 21756 41794 21812 41804
rect 22092 41972 22148 45164
rect 22204 43708 22260 46956
rect 22428 46452 22484 46462
rect 22428 46358 22484 46396
rect 22428 46116 22484 46126
rect 22428 45890 22484 46060
rect 22428 45838 22430 45890
rect 22482 45838 22484 45890
rect 22428 45826 22484 45838
rect 22316 44212 22372 44222
rect 22316 44210 22484 44212
rect 22316 44158 22318 44210
rect 22370 44158 22484 44210
rect 22316 44156 22484 44158
rect 22316 44146 22372 44156
rect 22204 43652 22372 43708
rect 22204 43540 22260 43550
rect 22204 43446 22260 43484
rect 22092 41748 22148 41916
rect 22092 41682 22148 41692
rect 21644 41412 21700 41422
rect 21644 41186 21700 41356
rect 21644 41134 21646 41186
rect 21698 41134 21700 41186
rect 21644 41122 21700 41134
rect 22092 41186 22148 41198
rect 22092 41134 22094 41186
rect 22146 41134 22148 41186
rect 21756 41076 21812 41086
rect 21756 40982 21812 41020
rect 21868 41074 21924 41086
rect 21868 41022 21870 41074
rect 21922 41022 21924 41074
rect 21868 40964 21924 41022
rect 21532 40908 21700 40964
rect 21532 40404 21588 40414
rect 21532 40290 21588 40348
rect 21532 40238 21534 40290
rect 21586 40238 21588 40290
rect 21532 40226 21588 40238
rect 21420 40114 21476 40124
rect 21308 39890 21364 39900
rect 21532 39620 21588 39630
rect 21532 38722 21588 39564
rect 21644 38834 21700 40908
rect 21868 40628 21924 40908
rect 21868 40562 21924 40572
rect 21756 40292 21812 40302
rect 21756 40198 21812 40236
rect 21980 40180 22036 40190
rect 21980 40086 22036 40124
rect 22092 39620 22148 41134
rect 22316 39732 22372 43652
rect 22428 43092 22484 44156
rect 22764 43316 22820 47180
rect 22988 45220 23044 50428
rect 23324 49922 23380 51550
rect 23436 50428 23492 51886
rect 23772 51378 23828 53004
rect 23884 52162 23940 53676
rect 23884 52110 23886 52162
rect 23938 52110 23940 52162
rect 23884 52098 23940 52110
rect 23996 53506 24052 53518
rect 23996 53454 23998 53506
rect 24050 53454 24052 53506
rect 23772 51326 23774 51378
rect 23826 51326 23828 51378
rect 23772 51314 23828 51326
rect 23436 50372 23604 50428
rect 23324 49870 23326 49922
rect 23378 49870 23380 49922
rect 23324 49858 23380 49870
rect 23548 49922 23604 50372
rect 23548 49870 23550 49922
rect 23602 49870 23604 49922
rect 23548 49858 23604 49870
rect 23884 50034 23940 50046
rect 23884 49982 23886 50034
rect 23938 49982 23940 50034
rect 23100 49026 23156 49038
rect 23100 48974 23102 49026
rect 23154 48974 23156 49026
rect 23100 48020 23156 48974
rect 23660 49026 23716 49038
rect 23660 48974 23662 49026
rect 23714 48974 23716 49026
rect 23660 48804 23716 48974
rect 23660 48738 23716 48748
rect 23100 47954 23156 47964
rect 23212 48020 23268 48030
rect 23212 48018 23828 48020
rect 23212 47966 23214 48018
rect 23266 47966 23828 48018
rect 23212 47964 23828 47966
rect 23212 47954 23268 47964
rect 23548 45778 23604 45790
rect 23548 45726 23550 45778
rect 23602 45726 23604 45778
rect 22988 45154 23044 45164
rect 23212 45220 23268 45230
rect 23212 45218 23380 45220
rect 23212 45166 23214 45218
rect 23266 45166 23380 45218
rect 23212 45164 23380 45166
rect 23212 45154 23268 45164
rect 22876 45106 22932 45118
rect 22876 45054 22878 45106
rect 22930 45054 22932 45106
rect 22876 44100 22932 45054
rect 23324 44212 23380 45164
rect 23436 44212 23492 44222
rect 23324 44156 23436 44212
rect 23436 44146 23492 44156
rect 22876 44044 23268 44100
rect 22876 43540 22932 44044
rect 22876 43474 22932 43484
rect 23212 43538 23268 44044
rect 23548 43708 23604 45726
rect 23212 43486 23214 43538
rect 23266 43486 23268 43538
rect 23212 43474 23268 43486
rect 23436 43652 23604 43708
rect 23660 44322 23716 44334
rect 23660 44270 23662 44322
rect 23714 44270 23716 44322
rect 22764 43260 23380 43316
rect 22428 43026 22484 43036
rect 22988 43092 23044 43102
rect 23044 43036 23156 43092
rect 22988 43026 23044 43036
rect 22988 42868 23044 42878
rect 22764 42082 22820 42094
rect 22764 42030 22766 42082
rect 22818 42030 22820 42082
rect 22540 41972 22596 41982
rect 22428 41970 22596 41972
rect 22428 41918 22542 41970
rect 22594 41918 22596 41970
rect 22428 41916 22596 41918
rect 22428 41412 22484 41916
rect 22540 41906 22596 41916
rect 22428 41346 22484 41356
rect 22540 41748 22596 41758
rect 22540 41410 22596 41692
rect 22764 41524 22820 42030
rect 22876 42084 22932 42094
rect 22876 41990 22932 42028
rect 22988 41748 23044 42812
rect 22988 41682 23044 41692
rect 22764 41458 22820 41468
rect 22540 41358 22542 41410
rect 22594 41358 22596 41410
rect 22540 41346 22596 41358
rect 22988 41188 23044 41198
rect 23100 41188 23156 43036
rect 22988 41186 23156 41188
rect 22988 41134 22990 41186
rect 23042 41134 23156 41186
rect 22988 41132 23156 41134
rect 22988 41122 23044 41132
rect 23100 40962 23156 40974
rect 23100 40910 23102 40962
rect 23154 40910 23156 40962
rect 22428 40628 22484 40638
rect 22428 40534 22484 40572
rect 23100 40404 23156 40910
rect 23100 40338 23156 40348
rect 23212 40962 23268 40974
rect 23212 40910 23214 40962
rect 23266 40910 23268 40962
rect 22764 40180 22820 40190
rect 22316 39676 22708 39732
rect 21644 38782 21646 38834
rect 21698 38782 21700 38834
rect 21644 38770 21700 38782
rect 21756 39564 22148 39620
rect 21532 38670 21534 38722
rect 21586 38670 21588 38722
rect 21532 38658 21588 38670
rect 21756 38668 21812 39564
rect 22428 39508 22484 39518
rect 20748 38098 20804 38108
rect 21644 38612 21812 38668
rect 22092 38724 22148 38762
rect 22092 38658 22148 38668
rect 21644 38050 21700 38612
rect 22092 38164 22148 38174
rect 22092 38070 22148 38108
rect 21644 37998 21646 38050
rect 21698 37998 21700 38050
rect 21644 37986 21700 37998
rect 21308 37938 21364 37950
rect 21308 37886 21310 37938
rect 21362 37886 21364 37938
rect 21308 37492 21364 37886
rect 21420 37828 21476 37838
rect 21420 37826 21588 37828
rect 21420 37774 21422 37826
rect 21474 37774 21588 37826
rect 21420 37772 21588 37774
rect 21420 37762 21476 37772
rect 21308 37426 21364 37436
rect 20076 37212 20244 37268
rect 19964 37156 20020 37166
rect 19852 37044 19908 37054
rect 19964 37044 20020 37100
rect 19852 37042 20020 37044
rect 19852 36990 19854 37042
rect 19906 36990 20020 37042
rect 19852 36988 20020 36990
rect 19852 36978 19908 36988
rect 18956 36540 19348 36596
rect 18620 36482 19236 36484
rect 18620 36430 18622 36482
rect 18674 36430 19236 36482
rect 18620 36428 19236 36430
rect 18620 36418 18676 36428
rect 18284 36372 18340 36382
rect 17724 36318 17726 36370
rect 17778 36318 17780 36370
rect 17724 36306 17780 36318
rect 17836 36370 18340 36372
rect 17836 36318 18286 36370
rect 18338 36318 18340 36370
rect 17836 36316 18340 36318
rect 17724 35700 17780 35710
rect 17836 35700 17892 36316
rect 18284 36306 18340 36316
rect 17724 35698 17892 35700
rect 17724 35646 17726 35698
rect 17778 35646 17892 35698
rect 17724 35644 17892 35646
rect 17612 35586 17668 35598
rect 17612 35534 17614 35586
rect 17666 35534 17668 35586
rect 17388 35474 17444 35486
rect 17388 35422 17390 35474
rect 17442 35422 17444 35474
rect 17388 34916 17444 35422
rect 17388 34850 17444 34860
rect 16940 34626 16996 34636
rect 17052 34802 17108 34814
rect 17052 34750 17054 34802
rect 17106 34750 17108 34802
rect 17052 34580 17108 34750
rect 17052 34524 17556 34580
rect 17500 34354 17556 34524
rect 17500 34302 17502 34354
rect 17554 34302 17556 34354
rect 17500 34290 17556 34302
rect 17388 34132 17444 34142
rect 16268 33954 16324 33964
rect 16604 34020 16660 34030
rect 16828 34020 16884 34076
rect 17276 34130 17444 34132
rect 17276 34078 17390 34130
rect 17442 34078 17444 34130
rect 17276 34076 17444 34078
rect 16828 33964 17220 34020
rect 16604 33926 16660 33964
rect 15596 33908 15652 33918
rect 15596 33814 15652 33852
rect 17164 33684 17220 33964
rect 17164 33570 17220 33628
rect 17164 33518 17166 33570
rect 17218 33518 17220 33570
rect 17164 33506 17220 33518
rect 15260 32338 15316 32350
rect 15260 32286 15262 32338
rect 15314 32286 15316 32338
rect 15260 32004 15316 32286
rect 15260 31938 15316 31948
rect 15484 31780 15540 33404
rect 16828 33348 16884 33358
rect 17276 33348 17332 34076
rect 17388 34066 17444 34076
rect 17612 34130 17668 35534
rect 17612 34078 17614 34130
rect 17666 34078 17668 34130
rect 17612 34066 17668 34078
rect 17724 34020 17780 35644
rect 19180 35026 19236 36428
rect 19180 34974 19182 35026
rect 19234 34974 19236 35026
rect 19180 34962 19236 34974
rect 17388 33460 17444 33470
rect 17724 33460 17780 33964
rect 19180 34020 19236 34030
rect 17836 33906 17892 33918
rect 17836 33854 17838 33906
rect 17890 33854 17892 33906
rect 17836 33572 17892 33854
rect 19068 33684 19124 33694
rect 17836 33506 17892 33516
rect 18732 33572 18788 33582
rect 18732 33478 18788 33516
rect 19068 33570 19124 33628
rect 19068 33518 19070 33570
rect 19122 33518 19124 33570
rect 19068 33506 19124 33518
rect 17388 33458 17780 33460
rect 17388 33406 17390 33458
rect 17442 33406 17780 33458
rect 17388 33404 17780 33406
rect 17388 33394 17444 33404
rect 16884 33292 17332 33348
rect 18956 33348 19012 33358
rect 16828 33254 16884 33292
rect 18956 33254 19012 33292
rect 18620 33236 18676 33246
rect 15484 31686 15540 31724
rect 18172 33234 18676 33236
rect 18172 33182 18622 33234
rect 18674 33182 18676 33234
rect 18172 33180 18676 33182
rect 18172 31106 18228 33180
rect 18620 33170 18676 33180
rect 19180 33124 19236 33964
rect 19292 33460 19348 36540
rect 21532 36372 21588 37772
rect 21532 36316 21924 36372
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 21868 35924 21924 36316
rect 22428 36260 22484 39452
rect 22652 38836 22708 39676
rect 22764 39618 22820 40124
rect 22764 39566 22766 39618
rect 22818 39566 22820 39618
rect 22764 39508 22820 39566
rect 22988 39620 23044 39630
rect 22988 39526 23044 39564
rect 22764 39442 22820 39452
rect 23212 39172 23268 40910
rect 23324 40740 23380 43260
rect 23436 42084 23492 43652
rect 23548 43538 23604 43550
rect 23548 43486 23550 43538
rect 23602 43486 23604 43538
rect 23548 43204 23604 43486
rect 23548 43138 23604 43148
rect 23660 43538 23716 44270
rect 23772 44212 23828 47964
rect 23884 44324 23940 49982
rect 23996 49810 24052 53454
rect 24108 53060 24164 53070
rect 24108 52946 24164 53004
rect 24108 52894 24110 52946
rect 24162 52894 24164 52946
rect 24108 52882 24164 52894
rect 24220 52948 24276 52958
rect 24220 52834 24276 52892
rect 24220 52782 24222 52834
rect 24274 52782 24276 52834
rect 24108 51492 24164 51502
rect 24220 51492 24276 52782
rect 24108 51490 24276 51492
rect 24108 51438 24110 51490
rect 24162 51438 24276 51490
rect 24108 51436 24276 51438
rect 24108 51426 24164 51436
rect 24332 50428 24388 59724
rect 24444 59714 24500 59724
rect 25116 58436 25172 59838
rect 24780 58380 25172 58436
rect 24780 58322 24836 58380
rect 24780 58270 24782 58322
rect 24834 58270 24836 58322
rect 24780 58258 24836 58270
rect 24444 57652 24500 57662
rect 24444 57558 24500 57596
rect 25004 57092 25060 58380
rect 25116 58210 25172 58222
rect 25116 58158 25118 58210
rect 25170 58158 25172 58210
rect 25116 57428 25172 58158
rect 25452 57540 25508 62300
rect 25564 60004 25620 62524
rect 25676 61460 25732 61470
rect 25676 60674 25732 61404
rect 25788 61458 25844 62860
rect 25900 62468 25956 62972
rect 26236 62962 26292 62972
rect 25900 62402 25956 62412
rect 26572 62188 26628 66782
rect 26684 66500 26740 68460
rect 27580 67170 27636 67182
rect 27580 67118 27582 67170
rect 27634 67118 27636 67170
rect 26796 67060 26852 67070
rect 26796 66966 26852 67004
rect 27020 67060 27076 67070
rect 27468 67060 27524 67070
rect 27020 67058 27524 67060
rect 27020 67006 27022 67058
rect 27074 67006 27470 67058
rect 27522 67006 27524 67058
rect 27020 67004 27524 67006
rect 27020 66994 27076 67004
rect 27468 66994 27524 67004
rect 27580 66948 27636 67118
rect 27580 66882 27636 66892
rect 27356 66836 27412 66846
rect 27356 66742 27412 66780
rect 26796 66500 26852 66510
rect 26684 66498 26852 66500
rect 26684 66446 26798 66498
rect 26850 66446 26852 66498
rect 26684 66444 26852 66446
rect 26796 66434 26852 66444
rect 25788 61406 25790 61458
rect 25842 61406 25844 61458
rect 25788 61394 25844 61406
rect 26348 62132 26628 62188
rect 26684 66274 26740 66286
rect 26684 66222 26686 66274
rect 26738 66222 26740 66274
rect 26684 66052 26740 66222
rect 27244 66052 27300 66062
rect 26684 66050 27300 66052
rect 26684 65998 27246 66050
rect 27298 65998 27300 66050
rect 26684 65996 27300 65998
rect 25676 60622 25678 60674
rect 25730 60622 25732 60674
rect 25676 60610 25732 60622
rect 25676 60004 25732 60014
rect 25564 59948 25676 60004
rect 25676 59108 25732 59948
rect 25788 59892 25844 59902
rect 26236 59892 26292 59902
rect 25788 59890 26292 59892
rect 25788 59838 25790 59890
rect 25842 59838 26238 59890
rect 26290 59838 26292 59890
rect 25788 59836 26292 59838
rect 25788 59826 25844 59836
rect 26236 59826 26292 59836
rect 25900 59108 25956 59118
rect 25676 59052 25900 59108
rect 25900 59014 25956 59052
rect 26348 58996 26404 62132
rect 26572 60676 26628 60686
rect 26572 59890 26628 60620
rect 26572 59838 26574 59890
rect 26626 59838 26628 59890
rect 26572 59826 26628 59838
rect 26012 58940 26404 58996
rect 26460 59108 26516 59118
rect 25900 58660 25956 58670
rect 26012 58660 26068 58940
rect 25900 58658 26068 58660
rect 25900 58606 25902 58658
rect 25954 58606 26068 58658
rect 25900 58604 26068 58606
rect 25900 58594 25956 58604
rect 25564 58548 25620 58558
rect 25564 58454 25620 58492
rect 25676 58436 25732 58446
rect 25676 58342 25732 58380
rect 25564 58212 25620 58222
rect 25564 58118 25620 58156
rect 26012 57650 26068 57662
rect 26012 57598 26014 57650
rect 26066 57598 26068 57650
rect 25676 57540 25732 57550
rect 25452 57538 25732 57540
rect 25452 57486 25678 57538
rect 25730 57486 25732 57538
rect 25452 57484 25732 57486
rect 25116 57362 25172 57372
rect 25676 57426 25732 57484
rect 26012 57538 26068 57598
rect 26012 57486 26014 57538
rect 26066 57486 26068 57538
rect 26012 57474 26068 57486
rect 25676 57374 25678 57426
rect 25730 57374 25732 57426
rect 25340 57092 25396 57102
rect 24668 57090 25620 57092
rect 24668 57038 25342 57090
rect 25394 57038 25620 57090
rect 24668 57036 25620 57038
rect 24444 56866 24500 56878
rect 24444 56814 24446 56866
rect 24498 56814 24500 56866
rect 24444 56532 24500 56814
rect 24668 56866 24724 57036
rect 25340 57026 25396 57036
rect 24668 56814 24670 56866
rect 24722 56814 24724 56866
rect 24668 56802 24724 56814
rect 25116 56866 25172 56878
rect 25116 56814 25118 56866
rect 25170 56814 25172 56866
rect 24780 56756 24836 56766
rect 24780 56662 24836 56700
rect 24444 56466 24500 56476
rect 25116 56532 25172 56814
rect 25116 56466 25172 56476
rect 24556 56196 24612 56206
rect 24556 56102 24612 56140
rect 24444 56082 24500 56094
rect 24444 56030 24446 56082
rect 24498 56030 24500 56082
rect 24444 55300 24500 56030
rect 24780 56084 24836 56094
rect 25340 56084 25396 56094
rect 24780 56082 25396 56084
rect 24780 56030 24782 56082
rect 24834 56030 25342 56082
rect 25394 56030 25396 56082
rect 24780 56028 25396 56030
rect 24780 56018 24836 56028
rect 24444 55234 24500 55244
rect 25340 55186 25396 56028
rect 25564 56082 25620 57036
rect 25676 56980 25732 57374
rect 26236 57092 26292 58940
rect 26236 57026 26292 57036
rect 26348 58772 26404 58782
rect 26348 57428 26404 58716
rect 25676 56914 25732 56924
rect 25676 56644 25732 56654
rect 25676 56550 25732 56588
rect 25564 56030 25566 56082
rect 25618 56030 25620 56082
rect 25564 56018 25620 56030
rect 25788 56532 25844 56542
rect 25788 55860 25844 56476
rect 25900 56084 25956 56094
rect 25900 55990 25956 56028
rect 25788 55766 25844 55804
rect 26348 55298 26404 57372
rect 26348 55246 26350 55298
rect 26402 55246 26404 55298
rect 26348 55234 26404 55246
rect 25340 55134 25342 55186
rect 25394 55134 25396 55186
rect 25340 55122 25396 55134
rect 26460 55076 26516 59052
rect 26124 55020 26516 55076
rect 25452 54626 25508 54638
rect 25452 54574 25454 54626
rect 25506 54574 25508 54626
rect 25340 54402 25396 54414
rect 25340 54350 25342 54402
rect 25394 54350 25396 54402
rect 25228 54290 25284 54302
rect 25228 54238 25230 54290
rect 25282 54238 25284 54290
rect 24444 53730 24500 53742
rect 24444 53678 24446 53730
rect 24498 53678 24500 53730
rect 24444 53508 24500 53678
rect 25004 53620 25060 53630
rect 24444 53442 24500 53452
rect 24668 53618 25060 53620
rect 24668 53566 25006 53618
rect 25058 53566 25060 53618
rect 24668 53564 25060 53566
rect 24668 53060 24724 53564
rect 25004 53554 25060 53564
rect 24556 53058 24724 53060
rect 24556 53006 24670 53058
rect 24722 53006 24724 53058
rect 24556 53004 24724 53006
rect 24444 52052 24500 52062
rect 24444 51958 24500 51996
rect 23996 49758 23998 49810
rect 24050 49758 24052 49810
rect 23996 49746 24052 49758
rect 24108 50372 24388 50428
rect 23996 48468 24052 48478
rect 23996 48354 24052 48412
rect 23996 48302 23998 48354
rect 24050 48302 24052 48354
rect 23996 48290 24052 48302
rect 24108 48354 24164 50372
rect 24556 49924 24612 53004
rect 24668 52994 24724 53004
rect 25228 51828 25284 54238
rect 25340 53620 25396 54350
rect 25340 53554 25396 53564
rect 25228 51762 25284 51772
rect 24668 51380 24724 51390
rect 24668 51286 24724 51324
rect 24556 49858 24612 49868
rect 25228 50484 25284 50494
rect 25452 50484 25508 54574
rect 25900 53732 25956 53742
rect 25900 52946 25956 53676
rect 25900 52894 25902 52946
rect 25954 52894 25956 52946
rect 25900 52882 25956 52894
rect 25676 51492 25732 51502
rect 25676 51398 25732 51436
rect 25284 50428 25508 50484
rect 24220 49138 24276 49150
rect 24220 49086 24222 49138
rect 24274 49086 24276 49138
rect 24220 48804 24276 49086
rect 24220 48738 24276 48748
rect 24108 48302 24110 48354
rect 24162 48302 24164 48354
rect 24108 47572 24164 48302
rect 25004 48468 25060 48478
rect 24220 48244 24276 48254
rect 24668 48244 24724 48254
rect 24220 48242 24500 48244
rect 24220 48190 24222 48242
rect 24274 48190 24500 48242
rect 24220 48188 24500 48190
rect 24220 48178 24276 48188
rect 24108 47506 24164 47516
rect 23996 47012 24052 47022
rect 23996 46114 24052 46956
rect 23996 46062 23998 46114
rect 24050 46062 24052 46114
rect 23996 46050 24052 46062
rect 24108 45780 24164 45790
rect 24108 45686 24164 45724
rect 23884 44268 24164 44324
rect 23772 44210 23940 44212
rect 23772 44158 23774 44210
rect 23826 44158 23940 44210
rect 23772 44156 23940 44158
rect 23772 44146 23828 44156
rect 23660 43486 23662 43538
rect 23714 43486 23716 43538
rect 23660 42868 23716 43486
rect 23884 43538 23940 44156
rect 23884 43486 23886 43538
rect 23938 43486 23940 43538
rect 23884 43474 23940 43486
rect 23660 42802 23716 42812
rect 23548 42084 23604 42094
rect 23436 42028 23548 42084
rect 23436 40964 23492 40974
rect 23436 40870 23492 40908
rect 23324 40684 23492 40740
rect 23324 40516 23380 40526
rect 23324 40422 23380 40460
rect 22652 38780 22820 38836
rect 22764 38722 22820 38780
rect 22764 38670 22766 38722
rect 22818 38670 22820 38722
rect 22540 38612 22596 38622
rect 22540 38610 22708 38612
rect 22540 38558 22542 38610
rect 22594 38558 22708 38610
rect 22540 38556 22708 38558
rect 22540 38546 22596 38556
rect 22652 38052 22708 38556
rect 22764 38052 22820 38670
rect 22876 38612 22932 38622
rect 22876 38610 23044 38612
rect 22876 38558 22878 38610
rect 22930 38558 23044 38610
rect 22876 38556 23044 38558
rect 22876 38546 22932 38556
rect 22876 38052 22932 38062
rect 22764 38050 22932 38052
rect 22764 37998 22878 38050
rect 22930 37998 22932 38050
rect 22764 37996 22932 37998
rect 22652 37958 22708 37996
rect 22876 37986 22932 37996
rect 22428 36204 22708 36260
rect 21868 35698 21924 35868
rect 22540 35924 22596 35934
rect 22540 35830 22596 35868
rect 22652 35812 22708 36204
rect 22652 35810 22820 35812
rect 22652 35758 22654 35810
rect 22706 35758 22820 35810
rect 22652 35756 22820 35758
rect 22652 35746 22708 35756
rect 21868 35646 21870 35698
rect 21922 35646 21924 35698
rect 21868 35634 21924 35646
rect 22092 35586 22148 35598
rect 22092 35534 22094 35586
rect 22146 35534 22148 35586
rect 21756 34914 21812 34926
rect 21756 34862 21758 34914
rect 21810 34862 21812 34914
rect 19292 33394 19348 33404
rect 19628 34692 19684 34702
rect 18956 33068 19236 33124
rect 18172 31054 18174 31106
rect 18226 31054 18228 31106
rect 18172 31042 18228 31054
rect 18620 32452 18676 32462
rect 18620 31892 18676 32396
rect 18956 32450 19012 33068
rect 18956 32398 18958 32450
rect 19010 32398 19012 32450
rect 18956 32386 19012 32398
rect 19628 32452 19684 34636
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 21084 34356 21140 34366
rect 21756 34356 21812 34862
rect 21084 34262 21140 34300
rect 21532 34300 21756 34356
rect 20076 34244 20132 34254
rect 20300 34244 20356 34254
rect 20076 34130 20132 34188
rect 20076 34078 20078 34130
rect 20130 34078 20132 34130
rect 20076 34066 20132 34078
rect 20188 34242 20356 34244
rect 20188 34190 20302 34242
rect 20354 34190 20356 34242
rect 20188 34188 20356 34190
rect 19740 33906 19796 33918
rect 19740 33854 19742 33906
rect 19794 33854 19796 33906
rect 19740 33684 19796 33854
rect 20188 33684 20244 34188
rect 20300 34178 20356 34188
rect 20524 34130 20580 34142
rect 20524 34078 20526 34130
rect 20578 34078 20580 34130
rect 20524 33908 20580 34078
rect 20636 34132 20692 34142
rect 20636 34038 20692 34076
rect 21420 34020 21476 34030
rect 21420 33926 21476 33964
rect 20636 33908 20692 33918
rect 19740 33618 19796 33628
rect 20076 33628 20244 33684
rect 20300 33852 20636 33908
rect 20076 33460 20132 33628
rect 20300 33572 20356 33852
rect 20636 33842 20692 33852
rect 21420 33796 21476 33806
rect 19964 33348 20020 33358
rect 20076 33348 20132 33404
rect 19964 33346 20132 33348
rect 19964 33294 19966 33346
rect 20018 33294 20132 33346
rect 19964 33292 20132 33294
rect 19964 33282 20020 33292
rect 20076 33124 20132 33292
rect 20188 33516 20356 33572
rect 20524 33684 20580 33694
rect 20188 33346 20244 33516
rect 20188 33294 20190 33346
rect 20242 33294 20244 33346
rect 20188 33282 20244 33294
rect 20300 33348 20356 33386
rect 20300 33282 20356 33292
rect 20524 33346 20580 33628
rect 21420 33570 21476 33740
rect 21420 33518 21422 33570
rect 21474 33518 21476 33570
rect 21420 33506 21476 33518
rect 21532 33684 21588 34300
rect 21756 34290 21812 34300
rect 22092 34356 22148 35534
rect 22204 35476 22260 35486
rect 22204 35382 22260 35420
rect 22204 35252 22260 35262
rect 22204 34914 22260 35196
rect 22764 35140 22820 35756
rect 22764 35074 22820 35084
rect 22876 35252 22932 35262
rect 22652 35028 22708 35038
rect 22652 34934 22708 34972
rect 22204 34862 22206 34914
rect 22258 34862 22260 34914
rect 22204 34850 22260 34862
rect 22764 34356 22820 34366
rect 22876 34356 22932 35196
rect 22092 34300 22372 34356
rect 21644 34132 21700 34142
rect 21980 34132 22036 34142
rect 21700 34130 22036 34132
rect 21700 34078 21982 34130
rect 22034 34078 22036 34130
rect 21700 34076 22036 34078
rect 21644 34038 21700 34076
rect 21980 34066 22036 34076
rect 22092 34020 22148 34300
rect 22316 34242 22372 34300
rect 22316 34190 22318 34242
rect 22370 34190 22372 34242
rect 22316 34178 22372 34190
rect 22428 34354 22932 34356
rect 22428 34302 22766 34354
rect 22818 34302 22932 34354
rect 22428 34300 22932 34302
rect 22092 33954 22148 33964
rect 21980 33908 22036 33918
rect 20524 33294 20526 33346
rect 20578 33294 20580 33346
rect 20524 33282 20580 33294
rect 21532 33348 21588 33628
rect 21756 33906 22036 33908
rect 21756 33854 21982 33906
rect 22034 33854 22036 33906
rect 21756 33852 22036 33854
rect 21644 33572 21700 33582
rect 21756 33572 21812 33852
rect 21980 33842 22036 33852
rect 22428 33908 22484 34300
rect 22764 34290 22820 34300
rect 21644 33570 21812 33572
rect 21644 33518 21646 33570
rect 21698 33518 21812 33570
rect 21644 33516 21812 33518
rect 21644 33506 21700 33516
rect 22316 33460 22372 33470
rect 22428 33460 22484 33852
rect 22316 33458 22484 33460
rect 22316 33406 22318 33458
rect 22370 33406 22484 33458
rect 22316 33404 22484 33406
rect 22316 33394 22372 33404
rect 21756 33348 21812 33358
rect 21532 33346 21812 33348
rect 21532 33294 21758 33346
rect 21810 33294 21812 33346
rect 21532 33292 21812 33294
rect 21756 33282 21812 33292
rect 21308 33236 21364 33246
rect 21084 33234 21364 33236
rect 21084 33182 21310 33234
rect 21362 33182 21364 33234
rect 21084 33180 21364 33182
rect 20076 33058 20132 33068
rect 20300 33124 20356 33134
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19628 32386 19684 32396
rect 14756 30940 15092 30996
rect 17500 30996 17556 31006
rect 14700 30902 14756 30940
rect 17500 30902 17556 30940
rect 18620 30996 18676 31836
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 18620 30930 18676 30940
rect 14252 30830 14254 30882
rect 14306 30830 14308 30882
rect 14252 30818 14308 30830
rect 20300 30882 20356 33068
rect 21084 32674 21140 33180
rect 21308 33170 21364 33180
rect 21084 32622 21086 32674
rect 21138 32622 21140 32674
rect 21084 32610 21140 32622
rect 22764 32788 22820 32798
rect 21868 32562 21924 32574
rect 21868 32510 21870 32562
rect 21922 32510 21924 32562
rect 21868 31948 21924 32510
rect 20748 31892 20804 31902
rect 20748 31220 20804 31836
rect 21756 31892 21924 31948
rect 22540 32004 22596 32014
rect 21756 31826 21812 31836
rect 22540 31778 22596 31948
rect 22540 31726 22542 31778
rect 22594 31726 22596 31778
rect 22540 31714 22596 31726
rect 22764 31778 22820 32732
rect 22764 31726 22766 31778
rect 22818 31726 22820 31778
rect 22652 31556 22708 31566
rect 21868 31554 22708 31556
rect 21868 31502 22654 31554
rect 22706 31502 22708 31554
rect 21868 31500 22708 31502
rect 20748 31218 20916 31220
rect 20748 31166 20750 31218
rect 20802 31166 20916 31218
rect 20748 31164 20916 31166
rect 20748 31154 20804 31164
rect 20300 30830 20302 30882
rect 20354 30830 20356 30882
rect 20300 30818 20356 30830
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 20860 30324 20916 31164
rect 21868 31106 21924 31500
rect 22652 31490 22708 31500
rect 22764 31220 22820 31726
rect 22876 31220 22932 31230
rect 22764 31218 22932 31220
rect 22764 31166 22878 31218
rect 22930 31166 22932 31218
rect 22764 31164 22932 31166
rect 22876 31154 22932 31164
rect 21868 31054 21870 31106
rect 21922 31054 21924 31106
rect 21868 31042 21924 31054
rect 22988 30996 23044 38556
rect 23100 35252 23156 35262
rect 23100 35026 23156 35196
rect 23100 34974 23102 35026
rect 23154 34974 23156 35026
rect 23100 34962 23156 34974
rect 23212 34468 23268 39116
rect 23324 39508 23380 39518
rect 23324 38946 23380 39452
rect 23324 38894 23326 38946
rect 23378 38894 23380 38946
rect 23324 38882 23380 38894
rect 23436 35252 23492 40684
rect 23548 38722 23604 42028
rect 24108 41748 24164 44268
rect 24332 43764 24388 43774
rect 24332 43650 24388 43708
rect 24332 43598 24334 43650
rect 24386 43598 24388 43650
rect 24332 43586 24388 43598
rect 24108 41186 24164 41692
rect 24444 41300 24500 48188
rect 24668 48150 24724 48188
rect 24556 47572 24612 47582
rect 24556 45778 24612 47516
rect 25004 47570 25060 48412
rect 25004 47518 25006 47570
rect 25058 47518 25060 47570
rect 25004 47506 25060 47518
rect 25228 46562 25284 50428
rect 26124 48468 26180 55020
rect 26684 54628 26740 65996
rect 27244 65986 27300 65996
rect 26796 63924 26852 63934
rect 26796 63830 26852 63868
rect 27468 63810 27524 63822
rect 27468 63758 27470 63810
rect 27522 63758 27524 63810
rect 27468 63250 27524 63758
rect 27468 63198 27470 63250
rect 27522 63198 27524 63250
rect 27468 63186 27524 63198
rect 27580 63140 27636 63150
rect 27692 63140 27748 70028
rect 35196 69804 35460 69814
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35196 69738 35460 69748
rect 28924 68626 28980 68638
rect 28924 68574 28926 68626
rect 28978 68574 28980 68626
rect 28252 68516 28308 68526
rect 28252 68422 28308 68460
rect 28924 68180 28980 68574
rect 35196 68236 35460 68246
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35196 68170 35460 68180
rect 28924 68114 28980 68124
rect 28588 67954 28644 67966
rect 28588 67902 28590 67954
rect 28642 67902 28644 67954
rect 28588 66948 28644 67902
rect 28588 66882 28644 66892
rect 35196 66668 35460 66678
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35196 66602 35460 66612
rect 35196 65100 35460 65110
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35196 65034 35460 65044
rect 38220 64482 38276 64494
rect 38220 64430 38222 64482
rect 38274 64430 38276 64482
rect 28476 63924 28532 63934
rect 28028 63140 28084 63150
rect 27580 63138 28084 63140
rect 27580 63086 27582 63138
rect 27634 63086 28030 63138
rect 28082 63086 28084 63138
rect 27580 63084 28084 63086
rect 26796 63028 26852 63038
rect 26796 62132 26852 62972
rect 26908 63028 26964 63038
rect 27244 63028 27300 63038
rect 26908 63026 27300 63028
rect 26908 62974 26910 63026
rect 26962 62974 27246 63026
rect 27298 62974 27300 63026
rect 26908 62972 27300 62974
rect 26908 62962 26964 62972
rect 27244 62962 27300 62972
rect 26796 61572 26852 62076
rect 27020 62468 27076 62478
rect 26908 61572 26964 61582
rect 26796 61570 26964 61572
rect 26796 61518 26910 61570
rect 26962 61518 26964 61570
rect 26796 61516 26964 61518
rect 26908 61506 26964 61516
rect 27020 61458 27076 62412
rect 27020 61406 27022 61458
rect 27074 61406 27076 61458
rect 27020 61394 27076 61406
rect 27132 61682 27188 61694
rect 27132 61630 27134 61682
rect 27186 61630 27188 61682
rect 27132 58772 27188 61630
rect 27580 60788 27636 63084
rect 28028 63074 28084 63084
rect 27132 58706 27188 58716
rect 27468 60732 27636 60788
rect 28476 62242 28532 63868
rect 38220 63924 38276 64430
rect 38220 63858 38276 63868
rect 29596 63810 29652 63822
rect 29596 63758 29598 63810
rect 29650 63758 29652 63810
rect 29036 62356 29092 62366
rect 29036 62262 29092 62300
rect 28476 62190 28478 62242
rect 28530 62190 28532 62242
rect 28476 60786 28532 62190
rect 29596 62132 29652 63758
rect 35196 63532 35460 63542
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35196 63466 35460 63476
rect 29596 62066 29652 62076
rect 35196 61964 35460 61974
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35196 61898 35460 61908
rect 28476 60734 28478 60786
rect 28530 60734 28532 60786
rect 26908 58548 26964 58558
rect 27468 58548 27524 60732
rect 28476 60722 28532 60734
rect 27804 60676 27860 60686
rect 27804 60582 27860 60620
rect 35196 60396 35460 60406
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35196 60330 35460 60340
rect 35196 58828 35460 58838
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35196 58762 35460 58772
rect 26908 58546 27524 58548
rect 26908 58494 26910 58546
rect 26962 58494 27524 58546
rect 26908 58492 27524 58494
rect 26908 58482 26964 58492
rect 27244 58322 27300 58334
rect 27244 58270 27246 58322
rect 27298 58270 27300 58322
rect 26236 54572 26740 54628
rect 26796 57092 26852 57102
rect 26236 51378 26292 54572
rect 26796 54516 26852 57036
rect 27244 57090 27300 58270
rect 27244 57038 27246 57090
rect 27298 57038 27300 57090
rect 27244 57026 27300 57038
rect 27468 58322 27524 58492
rect 27580 58548 27636 58558
rect 27580 58546 27860 58548
rect 27580 58494 27582 58546
rect 27634 58494 27860 58546
rect 27580 58492 27860 58494
rect 27580 58482 27636 58492
rect 27468 58270 27470 58322
rect 27522 58270 27524 58322
rect 26908 56866 26964 56878
rect 26908 56814 26910 56866
rect 26962 56814 26964 56866
rect 26908 56196 26964 56814
rect 27356 56866 27412 56878
rect 27356 56814 27358 56866
rect 27410 56814 27412 56866
rect 27356 56756 27412 56814
rect 27356 56690 27412 56700
rect 26908 56130 26964 56140
rect 27132 56082 27188 56094
rect 27132 56030 27134 56082
rect 27186 56030 27188 56082
rect 26572 54460 26852 54516
rect 26908 55298 26964 55310
rect 26908 55246 26910 55298
rect 26962 55246 26964 55298
rect 26572 53508 26628 54460
rect 26908 53956 26964 55246
rect 26796 53900 26964 53956
rect 27132 54514 27188 56030
rect 27356 55860 27412 55870
rect 27356 55186 27412 55804
rect 27356 55134 27358 55186
rect 27410 55134 27412 55186
rect 27356 55122 27412 55134
rect 27132 54462 27134 54514
rect 27186 54462 27188 54514
rect 26572 53452 26740 53508
rect 26572 52834 26628 52846
rect 26572 52782 26574 52834
rect 26626 52782 26628 52834
rect 26572 52386 26628 52782
rect 26572 52334 26574 52386
rect 26626 52334 26628 52386
rect 26572 52322 26628 52334
rect 26684 52386 26740 53452
rect 26796 53506 26852 53900
rect 26796 53454 26798 53506
rect 26850 53454 26852 53506
rect 26796 53060 26852 53454
rect 26908 53730 26964 53742
rect 26908 53678 26910 53730
rect 26962 53678 26964 53730
rect 26908 53508 26964 53678
rect 27132 53732 27188 54462
rect 27132 53666 27188 53676
rect 27244 53842 27300 53854
rect 27244 53790 27246 53842
rect 27298 53790 27300 53842
rect 26908 53442 26964 53452
rect 26796 52994 26852 53004
rect 27244 52836 27300 53790
rect 26684 52334 26686 52386
rect 26738 52334 26740 52386
rect 26572 51604 26628 51614
rect 26684 51604 26740 52334
rect 26908 52780 27300 52836
rect 27356 53508 27412 53518
rect 27356 52836 27412 53452
rect 26908 52386 26964 52780
rect 27356 52770 27412 52780
rect 27356 52388 27412 52398
rect 26908 52334 26910 52386
rect 26962 52334 26964 52386
rect 26908 52322 26964 52334
rect 27132 52386 27412 52388
rect 27132 52334 27358 52386
rect 27410 52334 27412 52386
rect 27132 52332 27412 52334
rect 27132 52162 27188 52332
rect 27356 52322 27412 52332
rect 27132 52110 27134 52162
rect 27186 52110 27188 52162
rect 27132 52098 27188 52110
rect 26572 51602 26740 51604
rect 26572 51550 26574 51602
rect 26626 51550 26740 51602
rect 26572 51548 26740 51550
rect 26572 51538 26628 51548
rect 26908 51492 26964 51502
rect 26964 51436 27412 51492
rect 26908 51398 26964 51436
rect 26236 51326 26238 51378
rect 26290 51326 26292 51378
rect 26236 50428 26292 51326
rect 27356 51266 27412 51436
rect 27356 51214 27358 51266
rect 27410 51214 27412 51266
rect 27356 51154 27412 51214
rect 27356 51102 27358 51154
rect 27410 51102 27412 51154
rect 26572 50594 26628 50606
rect 26572 50542 26574 50594
rect 26626 50542 26628 50594
rect 26572 50484 26628 50542
rect 27020 50484 27076 50494
rect 26572 50482 27076 50484
rect 26572 50430 27022 50482
rect 27074 50430 27076 50482
rect 26572 50428 27076 50430
rect 26236 50372 26516 50428
rect 27020 50372 27188 50428
rect 26460 50316 26964 50372
rect 26460 49028 26516 49038
rect 26348 48916 26404 48926
rect 26124 48374 26180 48412
rect 26236 48914 26404 48916
rect 26236 48862 26350 48914
rect 26402 48862 26404 48914
rect 26236 48860 26404 48862
rect 25564 48354 25620 48366
rect 25564 48302 25566 48354
rect 25618 48302 25620 48354
rect 25340 48244 25396 48254
rect 25564 48244 25620 48302
rect 26236 48244 26292 48860
rect 26348 48850 26404 48860
rect 26460 48692 26516 48972
rect 25564 48188 26292 48244
rect 26348 48636 26516 48692
rect 25340 48150 25396 48188
rect 25340 47572 25396 47582
rect 25340 47478 25396 47516
rect 25228 46510 25230 46562
rect 25282 46510 25284 46562
rect 25228 45890 25284 46510
rect 26124 46564 26180 46574
rect 25228 45838 25230 45890
rect 25282 45838 25284 45890
rect 25228 45826 25284 45838
rect 25676 46452 25732 46462
rect 25676 46002 25732 46396
rect 25676 45950 25678 46002
rect 25730 45950 25732 46002
rect 24556 45726 24558 45778
rect 24610 45726 24612 45778
rect 24556 45714 24612 45726
rect 24892 45778 24948 45790
rect 24892 45726 24894 45778
rect 24946 45726 24948 45778
rect 24892 44434 24948 45726
rect 24892 44382 24894 44434
rect 24946 44382 24948 44434
rect 24780 44212 24836 44222
rect 24780 44118 24836 44156
rect 24892 43652 24948 44382
rect 24892 43586 24948 43596
rect 25564 45332 25620 45342
rect 25564 43538 25620 45276
rect 25564 43486 25566 43538
rect 25618 43486 25620 43538
rect 25564 43474 25620 43486
rect 25564 43204 25620 43214
rect 25228 41970 25284 41982
rect 25228 41918 25230 41970
rect 25282 41918 25284 41970
rect 24444 41244 25060 41300
rect 24108 41134 24110 41186
rect 24162 41134 24164 41186
rect 24108 41122 24164 41134
rect 24780 41076 24836 41086
rect 24780 40982 24836 41020
rect 23996 40516 24052 40526
rect 23660 40292 23716 40302
rect 23660 40290 23828 40292
rect 23660 40238 23662 40290
rect 23714 40238 23828 40290
rect 23660 40236 23828 40238
rect 23660 40226 23716 40236
rect 23660 38836 23716 38846
rect 23772 38836 23828 40236
rect 23996 40290 24052 40460
rect 24332 40404 24388 40414
rect 24332 40402 24948 40404
rect 24332 40350 24334 40402
rect 24386 40350 24948 40402
rect 24332 40348 24948 40350
rect 24332 40338 24388 40348
rect 23996 40238 23998 40290
rect 24050 40238 24052 40290
rect 23996 40226 24052 40238
rect 24780 39618 24836 39630
rect 24780 39566 24782 39618
rect 24834 39566 24836 39618
rect 24332 38836 24388 38846
rect 23772 38834 24388 38836
rect 23772 38782 24334 38834
rect 24386 38782 24388 38834
rect 23772 38780 24388 38782
rect 23660 38742 23716 38780
rect 24332 38770 24388 38780
rect 23548 38670 23550 38722
rect 23602 38670 23604 38722
rect 23548 38658 23604 38670
rect 24444 38724 24500 38734
rect 24220 38500 24276 38510
rect 23772 38276 23828 38286
rect 24220 38276 24276 38444
rect 23772 38274 24276 38276
rect 23772 38222 23774 38274
rect 23826 38222 24276 38274
rect 23772 38220 24276 38222
rect 23772 38210 23828 38220
rect 24220 38162 24276 38220
rect 24444 38274 24500 38668
rect 24780 38724 24836 39566
rect 24780 38658 24836 38668
rect 24444 38222 24446 38274
rect 24498 38222 24500 38274
rect 24444 38210 24500 38222
rect 24780 38276 24836 38286
rect 24780 38182 24836 38220
rect 24220 38110 24222 38162
rect 24274 38110 24276 38162
rect 24220 38098 24276 38110
rect 23436 35186 23492 35196
rect 23548 38050 23604 38062
rect 24892 38052 24948 40348
rect 23548 37998 23550 38050
rect 23602 37998 23604 38050
rect 23100 34412 23268 34468
rect 23100 31556 23156 34412
rect 23548 32788 23604 37998
rect 24668 37996 24892 38052
rect 24668 36594 24724 37996
rect 24892 37958 24948 37996
rect 24668 36542 24670 36594
rect 24722 36542 24724 36594
rect 24668 36530 24724 36542
rect 24444 35252 24500 35262
rect 24444 34132 24500 35196
rect 25004 35028 25060 41244
rect 25228 41076 25284 41918
rect 25452 41748 25508 41758
rect 25452 41654 25508 41692
rect 25228 41010 25284 41020
rect 25564 39730 25620 43148
rect 25676 42756 25732 45950
rect 26012 45332 26068 45342
rect 26012 45238 26068 45276
rect 26124 45330 26180 46508
rect 26124 45278 26126 45330
rect 26178 45278 26180 45330
rect 26124 45266 26180 45278
rect 26236 44882 26292 44894
rect 26236 44830 26238 44882
rect 26290 44830 26292 44882
rect 26124 43538 26180 43550
rect 26124 43486 26126 43538
rect 26178 43486 26180 43538
rect 26124 42980 26180 43486
rect 26124 42914 26180 42924
rect 26236 42978 26292 44830
rect 26348 43540 26404 48636
rect 26796 48356 26852 48366
rect 26572 48300 26796 48356
rect 26460 48244 26516 48254
rect 26460 48150 26516 48188
rect 26572 47570 26628 48300
rect 26796 48262 26852 48300
rect 26572 47518 26574 47570
rect 26626 47518 26628 47570
rect 26572 47506 26628 47518
rect 26460 44322 26516 44334
rect 26460 44270 26462 44322
rect 26514 44270 26516 44322
rect 26460 43762 26516 44270
rect 26460 43710 26462 43762
rect 26514 43710 26516 43762
rect 26460 43698 26516 43710
rect 26348 43484 26516 43540
rect 26236 42926 26238 42978
rect 26290 42926 26292 42978
rect 26236 42914 26292 42926
rect 26012 42866 26068 42878
rect 26012 42814 26014 42866
rect 26066 42814 26068 42866
rect 25676 42754 25844 42756
rect 25676 42702 25678 42754
rect 25730 42702 25844 42754
rect 25676 42700 25844 42702
rect 25676 42690 25732 42700
rect 25676 41860 25732 41870
rect 25676 41766 25732 41804
rect 25788 40964 25844 42700
rect 25788 40898 25844 40908
rect 25900 41746 25956 41758
rect 25900 41694 25902 41746
rect 25954 41694 25956 41746
rect 25900 41076 25956 41694
rect 25900 40628 25956 41020
rect 25900 40562 25956 40572
rect 25564 39678 25566 39730
rect 25618 39678 25620 39730
rect 25564 39666 25620 39678
rect 25788 39508 25844 39518
rect 25564 39506 25844 39508
rect 25564 39454 25790 39506
rect 25842 39454 25844 39506
rect 25564 39452 25844 39454
rect 25340 39172 25396 39182
rect 25340 38946 25396 39116
rect 25340 38894 25342 38946
rect 25394 38894 25396 38946
rect 25340 38882 25396 38894
rect 25228 38836 25284 38846
rect 25228 38742 25284 38780
rect 25564 38500 25620 39452
rect 25788 39442 25844 39452
rect 26012 38948 26068 42814
rect 26236 41860 26292 41870
rect 26236 41186 26292 41804
rect 26348 41748 26404 41758
rect 26348 41654 26404 41692
rect 26236 41134 26238 41186
rect 26290 41134 26292 41186
rect 26236 41122 26292 41134
rect 26236 40964 26292 40974
rect 26236 39058 26292 40908
rect 26460 39620 26516 43484
rect 26796 43538 26852 43550
rect 26796 43486 26798 43538
rect 26850 43486 26852 43538
rect 26796 43204 26852 43486
rect 26796 43138 26852 43148
rect 26796 42980 26852 42990
rect 26796 42532 26852 42924
rect 26684 42530 26852 42532
rect 26684 42478 26798 42530
rect 26850 42478 26852 42530
rect 26684 42476 26852 42478
rect 26460 39564 26628 39620
rect 26236 39006 26238 39058
rect 26290 39006 26292 39058
rect 26124 38948 26180 38958
rect 25564 38434 25620 38444
rect 25676 38946 26180 38948
rect 25676 38894 26126 38946
rect 26178 38894 26180 38946
rect 25676 38892 26180 38894
rect 25452 38276 25508 38286
rect 25676 38276 25732 38892
rect 26124 38882 26180 38892
rect 26236 38612 26292 39006
rect 26124 38556 26292 38612
rect 26460 38834 26516 38846
rect 26460 38782 26462 38834
rect 26514 38782 26516 38834
rect 26460 38612 26516 38782
rect 26124 38500 26180 38556
rect 26460 38546 26516 38556
rect 25452 38162 25508 38220
rect 25452 38110 25454 38162
rect 25506 38110 25508 38162
rect 25340 37378 25396 37390
rect 25340 37326 25342 37378
rect 25394 37326 25396 37378
rect 25228 36932 25284 36942
rect 25228 35588 25284 36876
rect 25228 35522 25284 35532
rect 25004 34962 25060 34972
rect 25340 35476 25396 37326
rect 25452 37266 25508 38110
rect 25452 37214 25454 37266
rect 25506 37214 25508 37266
rect 25452 37202 25508 37214
rect 25564 38274 25732 38276
rect 25564 38222 25678 38274
rect 25730 38222 25732 38274
rect 25564 38220 25732 38222
rect 24668 34356 24724 34366
rect 24444 34130 24612 34132
rect 24444 34078 24446 34130
rect 24498 34078 24612 34130
rect 24444 34076 24612 34078
rect 24444 34066 24500 34076
rect 24556 33572 24612 34076
rect 24668 33796 24724 34300
rect 25340 34130 25396 35420
rect 25452 35474 25508 35486
rect 25452 35422 25454 35474
rect 25506 35422 25508 35474
rect 25452 34356 25508 35422
rect 25564 35476 25620 38220
rect 25676 38210 25732 38220
rect 25900 38444 26180 38500
rect 25900 37266 25956 38444
rect 26572 38388 26628 39564
rect 26684 38668 26740 42476
rect 26796 42466 26852 42476
rect 26796 41076 26852 41086
rect 26796 40982 26852 41020
rect 26908 39058 26964 50316
rect 27020 49028 27076 49038
rect 27020 48934 27076 48972
rect 27132 48580 27188 50372
rect 27020 48524 27188 48580
rect 27020 39172 27076 48524
rect 27132 48354 27188 48366
rect 27132 48302 27134 48354
rect 27186 48302 27188 48354
rect 27132 48244 27188 48302
rect 27132 47236 27188 48188
rect 27244 48356 27300 48366
rect 27244 47570 27300 48300
rect 27244 47518 27246 47570
rect 27298 47518 27300 47570
rect 27244 47506 27300 47518
rect 27132 47170 27188 47180
rect 27356 46788 27412 51102
rect 27468 50428 27524 58270
rect 27580 56868 27636 56878
rect 27580 56084 27636 56812
rect 27804 56194 27860 58492
rect 28476 57540 28532 57550
rect 28028 57092 28084 57102
rect 28028 56998 28084 57036
rect 28252 56868 28308 56878
rect 28252 56774 28308 56812
rect 28364 56866 28420 56878
rect 28364 56814 28366 56866
rect 28418 56814 28420 56866
rect 27804 56142 27806 56194
rect 27858 56142 27860 56194
rect 27804 56130 27860 56142
rect 27916 56754 27972 56766
rect 27916 56702 27918 56754
rect 27970 56702 27972 56754
rect 27580 53954 27636 56028
rect 27580 53902 27582 53954
rect 27634 53902 27636 53954
rect 27580 53890 27636 53902
rect 27692 55410 27748 55422
rect 27692 55358 27694 55410
rect 27746 55358 27748 55410
rect 27580 52386 27636 52398
rect 27580 52334 27582 52386
rect 27634 52334 27636 52386
rect 27580 52276 27636 52334
rect 27692 52276 27748 55358
rect 27804 54628 27860 54638
rect 27916 54628 27972 56702
rect 28364 55412 28420 56814
rect 28364 55346 28420 55356
rect 27804 54626 27972 54628
rect 27804 54574 27806 54626
rect 27858 54574 27972 54626
rect 27804 54572 27972 54574
rect 27804 54562 27860 54572
rect 28476 53732 28532 57484
rect 35196 57260 35460 57270
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35196 57194 35460 57204
rect 29036 56756 29092 56766
rect 29036 55298 29092 56700
rect 29372 56196 29428 56206
rect 29260 55412 29316 55422
rect 29260 55318 29316 55356
rect 29036 55246 29038 55298
rect 29090 55246 29092 55298
rect 29036 55234 29092 55246
rect 29372 55298 29428 56140
rect 29932 56196 29988 56206
rect 29932 55970 29988 56140
rect 29932 55918 29934 55970
rect 29986 55918 29988 55970
rect 29932 55906 29988 55918
rect 35196 55692 35460 55702
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35196 55626 35460 55636
rect 29372 55246 29374 55298
rect 29426 55246 29428 55298
rect 29372 55234 29428 55246
rect 29596 55300 29652 55310
rect 29652 55244 29988 55300
rect 29596 55206 29652 55244
rect 29932 54402 29988 55244
rect 29932 54350 29934 54402
rect 29986 54350 29988 54402
rect 29932 54338 29988 54350
rect 35980 54514 36036 54526
rect 35980 54462 35982 54514
rect 36034 54462 36036 54514
rect 35196 54124 35460 54134
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35196 54058 35460 54068
rect 28476 52948 28532 53676
rect 28476 52882 28532 52892
rect 33068 52948 33124 52958
rect 33068 52854 33124 52892
rect 28700 52836 28756 52846
rect 28700 52742 28756 52780
rect 33852 52836 33908 52846
rect 33852 52834 34132 52836
rect 33852 52782 33854 52834
rect 33906 52782 34132 52834
rect 33852 52780 34132 52782
rect 33852 52770 33908 52780
rect 27580 52274 27748 52276
rect 27580 52222 27582 52274
rect 27634 52222 27748 52274
rect 27580 52220 27748 52222
rect 27580 52210 27636 52220
rect 27692 51940 27748 52220
rect 32956 52164 33012 52174
rect 27692 51884 27972 51940
rect 27804 51266 27860 51278
rect 27804 51214 27806 51266
rect 27858 51214 27860 51266
rect 27804 51154 27860 51214
rect 27804 51102 27806 51154
rect 27858 51102 27860 51154
rect 27804 51090 27860 51102
rect 27916 50428 27972 51884
rect 32956 50818 33012 52108
rect 33740 52164 33796 52174
rect 33740 52070 33796 52108
rect 34076 52050 34132 52780
rect 35980 52834 36036 54462
rect 37996 54290 38052 54302
rect 37996 54238 37998 54290
rect 38050 54238 38052 54290
rect 37996 53172 38052 54238
rect 37996 53106 38052 53116
rect 35980 52782 35982 52834
rect 36034 52782 36036 52834
rect 35980 52770 36036 52782
rect 35196 52556 35460 52566
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35196 52490 35460 52500
rect 34076 51998 34078 52050
rect 34130 51998 34132 52050
rect 34076 51986 34132 51998
rect 37772 51378 37828 51390
rect 37772 51326 37774 51378
rect 37826 51326 37828 51378
rect 36764 51154 36820 51166
rect 36764 51102 36766 51154
rect 36818 51102 36820 51154
rect 35196 50988 35460 50998
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35196 50922 35460 50932
rect 32956 50766 32958 50818
rect 33010 50766 33012 50818
rect 32956 50754 33012 50766
rect 33180 50764 33572 50820
rect 33180 50428 33236 50764
rect 33516 50706 33572 50764
rect 33516 50654 33518 50706
rect 33570 50654 33572 50706
rect 33516 50642 33572 50654
rect 33292 50596 33348 50606
rect 33292 50594 33460 50596
rect 33292 50542 33294 50594
rect 33346 50542 33460 50594
rect 33292 50540 33460 50542
rect 33292 50530 33348 50540
rect 27468 50372 27636 50428
rect 27468 48356 27524 48366
rect 27468 48262 27524 48300
rect 27132 46732 27412 46788
rect 27132 43652 27188 46732
rect 27356 46564 27412 46574
rect 27356 46470 27412 46508
rect 27580 45332 27636 50372
rect 27580 45266 27636 45276
rect 27804 50372 27972 50428
rect 33068 50372 33236 50428
rect 27804 44548 27860 50372
rect 31164 49810 31220 49822
rect 31164 49758 31166 49810
rect 31218 49758 31220 49810
rect 28364 49698 28420 49710
rect 28364 49646 28366 49698
rect 28418 49646 28420 49698
rect 27916 49028 27972 49038
rect 27916 46676 27972 48972
rect 28028 48132 28084 48142
rect 28028 48038 28084 48076
rect 28364 47124 28420 49646
rect 30492 49700 30548 49710
rect 30492 49606 30548 49644
rect 29148 49140 29204 49150
rect 29148 49046 29204 49084
rect 30268 49140 30324 49150
rect 29932 48132 29988 48142
rect 29932 47570 29988 48076
rect 29932 47518 29934 47570
rect 29986 47518 29988 47570
rect 28364 47058 28420 47068
rect 29260 47124 29316 47134
rect 28028 46676 28084 46686
rect 27916 46674 28084 46676
rect 27916 46622 28030 46674
rect 28082 46622 28084 46674
rect 27916 46620 28084 46622
rect 28028 46610 28084 46620
rect 28588 46116 28644 46126
rect 27804 44492 27972 44548
rect 27468 43652 27524 43662
rect 27804 43652 27860 43662
rect 27132 43650 27412 43652
rect 27132 43598 27134 43650
rect 27186 43598 27412 43650
rect 27132 43596 27412 43598
rect 27132 43586 27188 43596
rect 27020 39106 27076 39116
rect 26908 39006 26910 39058
rect 26962 39006 26964 39058
rect 26908 38948 26964 39006
rect 26908 38892 27300 38948
rect 27020 38724 27076 38734
rect 26684 38612 26852 38668
rect 26460 38332 26628 38388
rect 26012 38276 26068 38286
rect 26012 38182 26068 38220
rect 26236 38052 26292 38062
rect 26236 37958 26292 37996
rect 26460 37380 26516 38332
rect 26460 37286 26516 37324
rect 26572 38162 26628 38174
rect 26572 38110 26574 38162
rect 26626 38110 26628 38162
rect 25900 37214 25902 37266
rect 25954 37214 25956 37266
rect 25900 37202 25956 37214
rect 26572 36708 26628 38110
rect 26684 38052 26740 38062
rect 26684 37938 26740 37996
rect 26684 37886 26686 37938
rect 26738 37886 26740 37938
rect 26684 37266 26740 37886
rect 26684 37214 26686 37266
rect 26738 37214 26740 37266
rect 26684 37202 26740 37214
rect 26796 36932 26852 38612
rect 26908 38276 26964 38286
rect 26908 38182 26964 38220
rect 26796 36866 26852 36876
rect 26908 37044 26964 37054
rect 25676 36652 26628 36708
rect 25676 35698 25732 36652
rect 26796 36372 26852 36382
rect 25788 36370 26852 36372
rect 25788 36318 26798 36370
rect 26850 36318 26852 36370
rect 25788 36316 26852 36318
rect 25788 35922 25844 36316
rect 26796 36306 26852 36316
rect 25788 35870 25790 35922
rect 25842 35870 25844 35922
rect 25788 35858 25844 35870
rect 25676 35646 25678 35698
rect 25730 35646 25732 35698
rect 25676 35634 25732 35646
rect 26908 35698 26964 36988
rect 26908 35646 26910 35698
rect 26962 35646 26964 35698
rect 26908 35634 26964 35646
rect 25788 35476 25844 35486
rect 25564 35474 25844 35476
rect 25564 35422 25790 35474
rect 25842 35422 25844 35474
rect 25564 35420 25844 35422
rect 25788 35410 25844 35420
rect 25452 34290 25508 34300
rect 25564 35140 25620 35150
rect 25564 34132 25620 35084
rect 25340 34078 25342 34130
rect 25394 34078 25396 34130
rect 25340 34066 25396 34078
rect 25452 34130 25620 34132
rect 25452 34078 25566 34130
rect 25618 34078 25620 34130
rect 25452 34076 25620 34078
rect 24668 33730 24724 33740
rect 23996 33516 24948 33572
rect 23996 33460 24052 33516
rect 23548 32674 23604 32732
rect 23548 32622 23550 32674
rect 23602 32622 23604 32674
rect 23548 32610 23604 32622
rect 23772 33458 24052 33460
rect 23772 33406 23998 33458
rect 24050 33406 24052 33458
rect 23772 33404 24052 33406
rect 23772 32674 23828 33404
rect 23996 33394 24052 33404
rect 24892 33458 24948 33516
rect 24892 33406 24894 33458
rect 24946 33406 24948 33458
rect 24892 33394 24948 33406
rect 24220 32788 24276 32798
rect 24220 32694 24276 32732
rect 23772 32622 23774 32674
rect 23826 32622 23828 32674
rect 23772 32610 23828 32622
rect 23212 32564 23268 32574
rect 23212 32004 23268 32508
rect 24332 32564 24388 32574
rect 24332 32470 24388 32508
rect 23212 31938 23268 31948
rect 23324 32450 23380 32462
rect 23324 32398 23326 32450
rect 23378 32398 23380 32450
rect 23212 31780 23268 31790
rect 23324 31780 23380 32398
rect 25340 32452 25396 32462
rect 25452 32452 25508 34076
rect 25564 34066 25620 34076
rect 26236 34020 26292 34030
rect 26012 34018 26292 34020
rect 26012 33966 26238 34018
rect 26290 33966 26292 34018
rect 26012 33964 26292 33966
rect 26012 33570 26068 33964
rect 26236 33954 26292 33964
rect 26012 33518 26014 33570
rect 26066 33518 26068 33570
rect 26012 33506 26068 33518
rect 26348 33460 26404 33470
rect 26348 33348 26404 33404
rect 26796 33460 26852 33470
rect 26796 33366 26852 33404
rect 26236 33346 26404 33348
rect 26236 33294 26350 33346
rect 26402 33294 26404 33346
rect 26236 33292 26404 33294
rect 26124 33124 26180 33134
rect 26124 33030 26180 33068
rect 25340 32450 25508 32452
rect 25340 32398 25342 32450
rect 25394 32398 25508 32450
rect 25340 32396 25508 32398
rect 25340 32386 25396 32396
rect 24220 32338 24276 32350
rect 24220 32286 24222 32338
rect 24274 32286 24276 32338
rect 23212 31778 23380 31780
rect 23212 31726 23214 31778
rect 23266 31726 23380 31778
rect 23212 31724 23380 31726
rect 23436 31890 23492 31902
rect 23436 31838 23438 31890
rect 23490 31838 23492 31890
rect 23212 31714 23268 31724
rect 23436 31556 23492 31838
rect 23100 31500 23492 31556
rect 23212 30996 23268 31006
rect 22988 30994 23268 30996
rect 22988 30942 23214 30994
rect 23266 30942 23268 30994
rect 22988 30940 23268 30942
rect 23436 30996 23492 31500
rect 23996 30996 24052 31006
rect 23436 30994 24052 30996
rect 23436 30942 23998 30994
rect 24050 30942 24052 30994
rect 23436 30940 24052 30942
rect 21980 30772 22036 30782
rect 21980 30770 22148 30772
rect 21980 30718 21982 30770
rect 22034 30718 22148 30770
rect 21980 30716 22148 30718
rect 21980 30706 22036 30716
rect 20860 30322 21364 30324
rect 20860 30270 20862 30322
rect 20914 30270 21364 30322
rect 20860 30268 21364 30270
rect 20860 30258 20916 30268
rect 21308 30210 21364 30268
rect 22092 30322 22148 30716
rect 22092 30270 22094 30322
rect 22146 30270 22148 30322
rect 22092 30258 22148 30270
rect 23212 30324 23268 30940
rect 23996 30930 24052 30940
rect 24220 30882 24276 32286
rect 25452 32004 25508 32014
rect 25452 31218 25508 31948
rect 26236 32004 26292 33292
rect 26348 33282 26404 33292
rect 25452 31166 25454 31218
rect 25506 31166 25508 31218
rect 25452 31154 25508 31166
rect 25564 31666 25620 31678
rect 25564 31614 25566 31666
rect 25618 31614 25620 31666
rect 24668 30996 24724 31006
rect 24668 30902 24724 30940
rect 25228 30996 25284 31006
rect 25228 30902 25284 30940
rect 24220 30830 24222 30882
rect 24274 30830 24276 30882
rect 24220 30818 24276 30830
rect 25564 30882 25620 31614
rect 26124 31220 26180 31230
rect 26236 31220 26292 31948
rect 26348 32564 26404 32574
rect 26348 31778 26404 32508
rect 26348 31726 26350 31778
rect 26402 31726 26404 31778
rect 26348 31714 26404 31726
rect 26124 31218 26292 31220
rect 26124 31166 26126 31218
rect 26178 31166 26292 31218
rect 26124 31164 26292 31166
rect 26124 31154 26180 31164
rect 27020 30996 27076 38668
rect 27132 38612 27188 38622
rect 27132 37266 27188 38556
rect 27132 37214 27134 37266
rect 27186 37214 27188 37266
rect 27132 37202 27188 37214
rect 27244 38050 27300 38892
rect 27244 37998 27246 38050
rect 27298 37998 27300 38050
rect 27132 36708 27188 36718
rect 27132 35252 27188 36652
rect 27132 35186 27188 35196
rect 27244 33460 27300 37998
rect 27356 38052 27412 43596
rect 27468 43558 27524 43596
rect 27580 43650 27860 43652
rect 27580 43598 27806 43650
rect 27858 43598 27860 43650
rect 27580 43596 27860 43598
rect 27580 42980 27636 43596
rect 27804 43586 27860 43596
rect 27580 42914 27636 42924
rect 27804 41970 27860 41982
rect 27804 41918 27806 41970
rect 27858 41918 27860 41970
rect 27804 41300 27860 41918
rect 27804 41234 27860 41244
rect 27804 41076 27860 41086
rect 27804 40962 27860 41020
rect 27804 40910 27806 40962
rect 27858 40910 27860 40962
rect 27804 40898 27860 40910
rect 27916 38500 27972 44492
rect 28028 43652 28084 43662
rect 28028 43540 28084 43596
rect 28588 43650 28644 46060
rect 28588 43598 28590 43650
rect 28642 43598 28644 43650
rect 28588 43586 28644 43598
rect 29260 45778 29316 47068
rect 29932 46116 29988 47518
rect 30156 47458 30212 47470
rect 30156 47406 30158 47458
rect 30210 47406 30212 47458
rect 30156 46676 30212 47406
rect 30156 46610 30212 46620
rect 29932 46050 29988 46060
rect 29260 45726 29262 45778
rect 29314 45726 29316 45778
rect 28364 43540 28420 43550
rect 28028 43538 28420 43540
rect 28028 43486 28030 43538
rect 28082 43486 28366 43538
rect 28418 43486 28420 43538
rect 28028 43484 28420 43486
rect 28028 43474 28084 43484
rect 28364 43474 28420 43484
rect 28700 43540 28756 43550
rect 28700 43204 28756 43484
rect 28364 43148 28756 43204
rect 28140 42868 28196 42878
rect 28140 42194 28196 42812
rect 28364 42754 28420 43148
rect 29260 43092 29316 45726
rect 29596 45890 29652 45902
rect 30044 45892 30100 45902
rect 29596 45838 29598 45890
rect 29650 45838 29652 45890
rect 29596 45106 29652 45838
rect 29596 45054 29598 45106
rect 29650 45054 29652 45106
rect 29596 43764 29652 45054
rect 29596 43698 29652 43708
rect 29932 45890 30100 45892
rect 29932 45838 30046 45890
rect 30098 45838 30100 45890
rect 29932 45836 30100 45838
rect 29596 43538 29652 43550
rect 29596 43486 29598 43538
rect 29650 43486 29652 43538
rect 29260 43036 29428 43092
rect 28364 42702 28366 42754
rect 28418 42702 28420 42754
rect 28364 42644 28420 42702
rect 28700 42980 28756 42990
rect 28700 42754 28756 42924
rect 28700 42702 28702 42754
rect 28754 42702 28756 42754
rect 28700 42690 28756 42702
rect 29260 42756 29316 42766
rect 28364 42578 28420 42588
rect 28476 42530 28532 42542
rect 28476 42478 28478 42530
rect 28530 42478 28532 42530
rect 28140 42142 28142 42194
rect 28194 42142 28196 42194
rect 28140 42130 28196 42142
rect 28252 42196 28308 42206
rect 28252 41970 28308 42140
rect 28476 42084 28532 42478
rect 28924 42308 28980 42318
rect 28476 42018 28532 42028
rect 28700 42252 28924 42308
rect 28252 41918 28254 41970
rect 28306 41918 28308 41970
rect 28252 41906 28308 41918
rect 28364 41970 28420 41982
rect 28364 41918 28366 41970
rect 28418 41918 28420 41970
rect 28364 41524 28420 41918
rect 28364 41458 28420 41468
rect 28700 41186 28756 42252
rect 28924 42242 28980 42252
rect 28700 41134 28702 41186
rect 28754 41134 28756 41186
rect 28700 41122 28756 41134
rect 29148 42084 29204 42094
rect 28364 41076 28420 41086
rect 29148 41076 29204 42028
rect 29260 41970 29316 42700
rect 29260 41918 29262 41970
rect 29314 41918 29316 41970
rect 29260 41906 29316 41918
rect 29372 42420 29428 43036
rect 29596 42980 29652 43486
rect 29596 42914 29652 42924
rect 29820 43538 29876 43550
rect 29820 43486 29822 43538
rect 29874 43486 29876 43538
rect 29484 42754 29540 42766
rect 29484 42702 29486 42754
rect 29538 42702 29540 42754
rect 29484 42644 29540 42702
rect 29484 42578 29540 42588
rect 29708 42754 29764 42766
rect 29708 42702 29710 42754
rect 29762 42702 29764 42754
rect 29372 41972 29428 42364
rect 29596 42532 29652 42542
rect 29484 41972 29540 41982
rect 29372 41970 29540 41972
rect 29372 41918 29486 41970
rect 29538 41918 29540 41970
rect 29372 41916 29540 41918
rect 29484 41906 29540 41916
rect 29372 41748 29428 41758
rect 29372 41410 29428 41692
rect 29372 41358 29374 41410
rect 29426 41358 29428 41410
rect 29372 41346 29428 41358
rect 29484 41524 29540 41534
rect 29260 41076 29316 41086
rect 29148 41074 29316 41076
rect 29148 41022 29262 41074
rect 29314 41022 29316 41074
rect 29148 41020 29316 41022
rect 28364 40982 28420 41020
rect 28476 40962 28532 40974
rect 28476 40910 28478 40962
rect 28530 40910 28532 40962
rect 28476 40628 28532 40910
rect 29260 40740 29316 41020
rect 29260 40674 29316 40684
rect 28476 40562 28532 40572
rect 27916 38444 28084 38500
rect 27580 38332 27972 38388
rect 27580 38274 27636 38332
rect 27580 38222 27582 38274
rect 27634 38222 27636 38274
rect 27580 38210 27636 38222
rect 27692 38164 27748 38174
rect 27356 37996 27636 38052
rect 27468 37826 27524 37838
rect 27468 37774 27470 37826
rect 27522 37774 27524 37826
rect 27356 37380 27412 37390
rect 27356 37266 27412 37324
rect 27356 37214 27358 37266
rect 27410 37214 27412 37266
rect 27356 36260 27412 37214
rect 27468 36260 27524 37774
rect 27580 36708 27636 37996
rect 27580 36642 27636 36652
rect 27692 37044 27748 38108
rect 27916 37380 27972 38332
rect 28028 38276 28084 38444
rect 28028 38164 28084 38220
rect 28028 38162 28532 38164
rect 28028 38110 28030 38162
rect 28082 38110 28532 38162
rect 28028 38108 28532 38110
rect 28028 38098 28084 38108
rect 28476 37490 28532 38108
rect 29484 38162 29540 41468
rect 29596 41298 29652 42476
rect 29708 42084 29764 42702
rect 29820 42308 29876 43486
rect 29820 42242 29876 42252
rect 29932 42196 29988 45836
rect 30044 45826 30100 45836
rect 30156 45106 30212 45118
rect 30156 45054 30158 45106
rect 30210 45054 30212 45106
rect 30156 43764 30212 45054
rect 30268 43988 30324 49084
rect 31164 49028 31220 49758
rect 32396 49700 32452 49710
rect 32396 49140 32452 49644
rect 32172 49084 32396 49140
rect 31164 48962 31220 48972
rect 31948 49028 32004 49038
rect 31948 48934 32004 48972
rect 31276 48914 31332 48926
rect 31276 48862 31278 48914
rect 31330 48862 31332 48914
rect 31276 48466 31332 48862
rect 31276 48414 31278 48466
rect 31330 48414 31332 48466
rect 31276 48356 31332 48414
rect 31276 48290 31332 48300
rect 32060 48916 32116 48926
rect 31836 48244 31892 48254
rect 31836 48150 31892 48188
rect 31836 47908 31892 47918
rect 31836 47570 31892 47852
rect 31836 47518 31838 47570
rect 31890 47518 31892 47570
rect 30492 47348 30548 47358
rect 30828 47348 30884 47358
rect 30492 47346 30884 47348
rect 30492 47294 30494 47346
rect 30546 47294 30830 47346
rect 30882 47294 30884 47346
rect 30492 47292 30884 47294
rect 30492 47282 30548 47292
rect 30828 47282 30884 47292
rect 31500 47236 31556 47246
rect 30828 46786 30884 46798
rect 30828 46734 30830 46786
rect 30882 46734 30884 46786
rect 30380 46004 30436 46014
rect 30828 46004 30884 46734
rect 31388 46788 31444 46798
rect 31500 46788 31556 47180
rect 31388 46786 31556 46788
rect 31388 46734 31390 46786
rect 31442 46734 31556 46786
rect 31388 46732 31556 46734
rect 31388 46722 31444 46732
rect 30380 46002 31444 46004
rect 30380 45950 30382 46002
rect 30434 45950 31444 46002
rect 30380 45948 31444 45950
rect 30380 45938 30436 45948
rect 31388 45890 31444 45948
rect 31388 45838 31390 45890
rect 31442 45838 31444 45890
rect 31388 45826 31444 45838
rect 30828 45220 30884 45230
rect 30828 45126 30884 45164
rect 30604 44324 30660 44334
rect 30940 44324 30996 44334
rect 30604 44322 30996 44324
rect 30604 44270 30606 44322
rect 30658 44270 30942 44322
rect 30994 44270 30996 44322
rect 30604 44268 30996 44270
rect 30604 44258 30660 44268
rect 30268 43932 30772 43988
rect 30716 43764 30772 43932
rect 30156 43708 30436 43764
rect 30044 43540 30100 43550
rect 30044 43446 30100 43484
rect 30268 43538 30324 43550
rect 30268 43486 30270 43538
rect 30322 43486 30324 43538
rect 30156 43314 30212 43326
rect 30156 43262 30158 43314
rect 30210 43262 30212 43314
rect 30044 42642 30100 42654
rect 30044 42590 30046 42642
rect 30098 42590 30100 42642
rect 30044 42308 30100 42590
rect 30156 42308 30212 43262
rect 30268 42868 30324 43486
rect 30268 42802 30324 42812
rect 30380 42420 30436 43708
rect 30716 43708 30884 43764
rect 30716 43650 30772 43708
rect 30716 43598 30718 43650
rect 30770 43598 30772 43650
rect 30716 43586 30772 43598
rect 30828 43650 30884 43708
rect 30828 43598 30830 43650
rect 30882 43598 30884 43650
rect 30828 43586 30884 43598
rect 30604 43314 30660 43326
rect 30604 43262 30606 43314
rect 30658 43262 30660 43314
rect 30604 42756 30660 43262
rect 30940 42756 30996 44268
rect 30604 42662 30660 42700
rect 30828 42700 30996 42756
rect 31164 43650 31220 43662
rect 31164 43598 31166 43650
rect 31218 43598 31220 43650
rect 30380 42364 30660 42420
rect 30156 42252 30436 42308
rect 30044 42242 30100 42252
rect 29932 42130 29988 42140
rect 30268 42084 30324 42094
rect 29708 42018 29764 42028
rect 30156 42082 30324 42084
rect 30156 42030 30270 42082
rect 30322 42030 30324 42082
rect 30156 42028 30324 42030
rect 30156 41972 30212 42028
rect 30268 42018 30324 42028
rect 29820 41916 30212 41972
rect 29708 41860 29764 41870
rect 29820 41860 29876 41916
rect 29708 41858 29876 41860
rect 29708 41806 29710 41858
rect 29762 41806 29876 41858
rect 29708 41804 29876 41806
rect 29708 41794 29764 41804
rect 29596 41246 29598 41298
rect 29650 41246 29652 41298
rect 29596 41234 29652 41246
rect 30044 41636 30100 41646
rect 30044 41076 30100 41580
rect 30044 40402 30100 41020
rect 30156 40626 30212 41916
rect 30380 41860 30436 42252
rect 30380 41794 30436 41804
rect 30156 40574 30158 40626
rect 30210 40574 30212 40626
rect 30156 40562 30212 40574
rect 30380 40628 30436 40638
rect 30492 40628 30548 42364
rect 30604 42082 30660 42364
rect 30604 42030 30606 42082
rect 30658 42030 30660 42082
rect 30604 42018 30660 42030
rect 30828 41972 30884 42700
rect 31164 42642 31220 43598
rect 31388 43540 31444 43550
rect 31500 43540 31556 46732
rect 31724 46788 31780 46798
rect 31724 46694 31780 46732
rect 31612 46676 31668 46686
rect 31612 45220 31668 46620
rect 31836 46564 31892 47518
rect 32060 46898 32116 48860
rect 32172 48354 32228 49084
rect 32396 49046 32452 49084
rect 32956 48802 33012 48814
rect 32956 48750 32958 48802
rect 33010 48750 33012 48802
rect 32508 48468 32564 48478
rect 32508 48374 32564 48412
rect 32172 48302 32174 48354
rect 32226 48302 32228 48354
rect 32172 48290 32228 48302
rect 32284 48354 32340 48366
rect 32284 48302 32286 48354
rect 32338 48302 32340 48354
rect 32284 47012 32340 48302
rect 32060 46846 32062 46898
rect 32114 46846 32116 46898
rect 32060 46834 32116 46846
rect 32172 46956 32340 47012
rect 32396 48356 32452 48366
rect 31948 46788 32004 46798
rect 31948 46694 32004 46732
rect 32172 46564 32228 46956
rect 32284 46788 32340 46798
rect 32396 46788 32452 48300
rect 32620 48244 32676 48254
rect 32620 47572 32676 48188
rect 32956 47796 33012 48750
rect 32956 47730 33012 47740
rect 33068 47684 33124 50372
rect 33292 49140 33348 49150
rect 33292 49026 33348 49084
rect 33404 49138 33460 50540
rect 33404 49086 33406 49138
rect 33458 49086 33460 49138
rect 33404 49074 33460 49086
rect 34860 49810 34916 49822
rect 34860 49758 34862 49810
rect 34914 49758 34916 49810
rect 33292 48974 33294 49026
rect 33346 48974 33348 49026
rect 33292 48242 33348 48974
rect 34860 49028 34916 49758
rect 36764 49812 36820 51102
rect 36764 49746 36820 49756
rect 35644 49698 35700 49710
rect 35644 49646 35646 49698
rect 35698 49646 35700 49698
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35196 49354 35460 49364
rect 35644 49138 35700 49646
rect 37772 49698 37828 51326
rect 37772 49646 37774 49698
rect 37826 49646 37828 49698
rect 37772 49634 37828 49646
rect 35644 49086 35646 49138
rect 35698 49086 35700 49138
rect 35644 49074 35700 49086
rect 34860 48962 34916 48972
rect 35084 49028 35140 49038
rect 34412 48916 34468 48926
rect 35084 48916 35140 48972
rect 35420 49028 35476 49038
rect 35420 48934 35476 48972
rect 35980 49026 36036 49038
rect 35980 48974 35982 49026
rect 36034 48974 36036 49026
rect 34412 48822 34468 48860
rect 34972 48860 35140 48916
rect 35980 48916 36036 48974
rect 33516 48802 33572 48814
rect 33516 48750 33518 48802
rect 33570 48750 33572 48802
rect 33516 48356 33572 48750
rect 33740 48804 33796 48814
rect 33740 48710 33796 48748
rect 34524 48804 34580 48814
rect 33628 48356 33684 48366
rect 33572 48354 33684 48356
rect 33572 48302 33630 48354
rect 33682 48302 33684 48354
rect 33572 48300 33684 48302
rect 33516 48262 33572 48300
rect 33628 48290 33684 48300
rect 33292 48190 33294 48242
rect 33346 48190 33348 48242
rect 33292 48178 33348 48190
rect 33180 48130 33236 48142
rect 33180 48078 33182 48130
rect 33234 48078 33236 48130
rect 33180 47908 33236 48078
rect 33180 47842 33236 47852
rect 34076 47908 34132 47918
rect 33740 47684 33796 47694
rect 33068 47682 33796 47684
rect 33068 47630 33742 47682
rect 33794 47630 33796 47682
rect 33068 47628 33796 47630
rect 32620 47516 33124 47572
rect 32620 47458 32676 47516
rect 32620 47406 32622 47458
rect 32674 47406 32676 47458
rect 32620 47394 32676 47406
rect 32284 46786 32452 46788
rect 32284 46734 32286 46786
rect 32338 46734 32452 46786
rect 32284 46732 32452 46734
rect 32956 47346 33012 47358
rect 32956 47294 32958 47346
rect 33010 47294 33012 47346
rect 32956 46788 33012 47294
rect 32284 46722 32340 46732
rect 32956 46722 33012 46732
rect 33068 46786 33124 47516
rect 33068 46734 33070 46786
rect 33122 46734 33124 46786
rect 33068 46722 33124 46734
rect 33180 47460 33236 47470
rect 31836 46508 32004 46564
rect 31948 45220 32004 46508
rect 31612 45154 31668 45164
rect 31836 45164 32004 45220
rect 32060 46508 32228 46564
rect 32508 46676 32564 46686
rect 31836 44772 31892 45164
rect 31948 44996 32004 45006
rect 31948 44902 32004 44940
rect 31836 44716 32004 44772
rect 31724 43652 31780 43662
rect 31724 43650 31892 43652
rect 31724 43598 31726 43650
rect 31778 43598 31892 43650
rect 31724 43596 31892 43598
rect 31724 43586 31780 43596
rect 31444 43484 31556 43540
rect 31164 42590 31166 42642
rect 31218 42590 31220 42642
rect 30940 42532 30996 42542
rect 30940 42438 30996 42476
rect 30716 41412 30772 41422
rect 30604 41356 30716 41412
rect 30604 41298 30660 41356
rect 30716 41346 30772 41356
rect 30604 41246 30606 41298
rect 30658 41246 30660 41298
rect 30604 41234 30660 41246
rect 30380 40626 30492 40628
rect 30380 40574 30382 40626
rect 30434 40574 30492 40626
rect 30380 40572 30492 40574
rect 30380 40562 30436 40572
rect 30492 40534 30548 40572
rect 30716 41076 30772 41086
rect 30716 40626 30772 41020
rect 30716 40574 30718 40626
rect 30770 40574 30772 40626
rect 30716 40562 30772 40574
rect 30044 40350 30046 40402
rect 30098 40350 30100 40402
rect 30044 40338 30100 40350
rect 30604 40404 30660 40414
rect 30604 40310 30660 40348
rect 29596 39732 29652 39742
rect 29596 39638 29652 39676
rect 30828 39732 30884 41916
rect 31052 41970 31108 41982
rect 31052 41918 31054 41970
rect 31106 41918 31108 41970
rect 31052 41636 31108 41918
rect 31052 41570 31108 41580
rect 31052 41186 31108 41198
rect 31052 41134 31054 41186
rect 31106 41134 31108 41186
rect 31052 40964 31108 41134
rect 31164 41188 31220 42590
rect 31276 42644 31332 42654
rect 31276 42420 31332 42588
rect 31276 42354 31332 42364
rect 31276 42196 31332 42206
rect 31276 42082 31332 42140
rect 31276 42030 31278 42082
rect 31330 42030 31332 42082
rect 31276 42018 31332 42030
rect 31388 41972 31444 43484
rect 31724 42868 31780 42878
rect 31612 42644 31668 42654
rect 31612 42550 31668 42588
rect 31724 42308 31780 42812
rect 31612 42252 31780 42308
rect 31500 41972 31556 41982
rect 31388 41970 31556 41972
rect 31388 41918 31502 41970
rect 31554 41918 31556 41970
rect 31388 41916 31556 41918
rect 31500 41906 31556 41916
rect 31612 41524 31668 42252
rect 31836 42196 31892 43596
rect 31948 42980 32004 44716
rect 32060 43204 32116 46508
rect 32396 46452 32452 46462
rect 32060 43138 32116 43148
rect 32172 46396 32396 46452
rect 32172 45218 32228 46396
rect 32396 46386 32452 46396
rect 32172 45166 32174 45218
rect 32226 45166 32228 45218
rect 32172 43762 32228 45166
rect 32172 43710 32174 43762
rect 32226 43710 32228 43762
rect 31948 42924 32116 42980
rect 31948 42756 32004 42766
rect 31948 42196 32004 42700
rect 32060 42642 32116 42924
rect 32060 42590 32062 42642
rect 32114 42590 32116 42642
rect 32060 42308 32116 42590
rect 32172 42644 32228 43710
rect 32284 46116 32340 46126
rect 32284 45778 32340 46060
rect 32284 45726 32286 45778
rect 32338 45726 32340 45778
rect 32284 43650 32340 45726
rect 32396 45666 32452 45678
rect 32396 45614 32398 45666
rect 32450 45614 32452 45666
rect 32396 45108 32452 45614
rect 32396 45014 32452 45052
rect 32284 43598 32286 43650
rect 32338 43598 32340 43650
rect 32284 43586 32340 43598
rect 32396 43538 32452 43550
rect 32396 43486 32398 43538
rect 32450 43486 32452 43538
rect 32396 42868 32452 43486
rect 32172 42578 32228 42588
rect 32284 42812 32452 42868
rect 32284 42530 32340 42812
rect 32508 42756 32564 46620
rect 33180 46564 33236 47404
rect 33068 46508 33236 46564
rect 33292 46674 33348 46686
rect 33292 46622 33294 46674
rect 33346 46622 33348 46674
rect 33068 45330 33124 46508
rect 33292 46452 33348 46622
rect 33292 46386 33348 46396
rect 33068 45278 33070 45330
rect 33122 45278 33124 45330
rect 33068 45266 33124 45278
rect 33180 45778 33236 45790
rect 33180 45726 33182 45778
rect 33234 45726 33236 45778
rect 33180 45220 33236 45726
rect 33292 45666 33348 45678
rect 33292 45614 33294 45666
rect 33346 45614 33348 45666
rect 33292 45332 33348 45614
rect 33292 45266 33348 45276
rect 33404 45666 33460 45678
rect 33404 45614 33406 45666
rect 33458 45614 33460 45666
rect 33180 45154 33236 45164
rect 33292 45108 33348 45118
rect 33404 45108 33460 45614
rect 33348 45052 33460 45108
rect 33292 45014 33348 45052
rect 33180 44996 33236 45006
rect 33516 44996 33572 47628
rect 33740 47618 33796 47628
rect 34076 47458 34132 47852
rect 34076 47406 34078 47458
rect 34130 47406 34132 47458
rect 34076 47394 34132 47406
rect 34300 47796 34356 47806
rect 34300 47458 34356 47740
rect 34300 47406 34302 47458
rect 34354 47406 34356 47458
rect 34300 47394 34356 47406
rect 33740 46676 33796 46686
rect 33740 46582 33796 46620
rect 34524 46564 34580 48748
rect 34636 48802 34692 48814
rect 34636 48750 34638 48802
rect 34690 48750 34692 48802
rect 34636 47460 34692 48750
rect 34748 48802 34804 48814
rect 34748 48750 34750 48802
rect 34802 48750 34804 48802
rect 34748 47684 34804 48750
rect 34860 48804 34916 48814
rect 34860 48710 34916 48748
rect 34748 47618 34804 47628
rect 34860 48130 34916 48142
rect 34860 48078 34862 48130
rect 34914 48078 34916 48130
rect 34860 47460 34916 48078
rect 34636 47404 34916 47460
rect 34636 46564 34692 46574
rect 34524 46562 34692 46564
rect 34524 46510 34638 46562
rect 34690 46510 34692 46562
rect 34524 46508 34692 46510
rect 34412 45332 34468 45342
rect 34076 45220 34132 45230
rect 34076 45106 34132 45164
rect 34076 45054 34078 45106
rect 34130 45054 34132 45106
rect 34076 45042 34132 45054
rect 34300 45108 34356 45118
rect 34300 45014 34356 45052
rect 32620 42868 32676 42878
rect 32620 42866 33124 42868
rect 32620 42814 32622 42866
rect 32674 42814 33124 42866
rect 32620 42812 33124 42814
rect 32620 42802 32676 42812
rect 32284 42478 32286 42530
rect 32338 42478 32340 42530
rect 32284 42308 32340 42478
rect 32060 42252 32228 42308
rect 31948 42140 32116 42196
rect 31836 42130 31892 42140
rect 31500 41468 31668 41524
rect 31724 41970 31780 41982
rect 31724 41918 31726 41970
rect 31778 41918 31780 41970
rect 31388 41300 31444 41310
rect 31388 41206 31444 41244
rect 31276 41188 31332 41198
rect 31164 41186 31332 41188
rect 31164 41134 31278 41186
rect 31330 41134 31332 41186
rect 31164 41132 31332 41134
rect 31500 41188 31556 41468
rect 31724 41412 31780 41918
rect 31948 41970 32004 41982
rect 31948 41918 31950 41970
rect 32002 41918 32004 41970
rect 31724 41346 31780 41356
rect 31836 41524 31892 41534
rect 31724 41188 31780 41198
rect 31500 41186 31780 41188
rect 31500 41134 31726 41186
rect 31778 41134 31780 41186
rect 31500 41132 31780 41134
rect 31276 41122 31332 41132
rect 31724 41122 31780 41132
rect 31836 41074 31892 41468
rect 31836 41022 31838 41074
rect 31890 41022 31892 41074
rect 31052 40898 31108 40908
rect 31500 40964 31556 40974
rect 31388 40852 31444 40862
rect 30940 40628 30996 40638
rect 30940 40402 30996 40572
rect 30940 40350 30942 40402
rect 30994 40350 30996 40402
rect 30940 40338 30996 40350
rect 31388 40402 31444 40796
rect 31500 40628 31556 40908
rect 31836 40852 31892 41022
rect 31948 41076 32004 41918
rect 31948 41010 32004 41020
rect 32060 40964 32116 42140
rect 32060 40898 32116 40908
rect 31836 40786 31892 40796
rect 31948 40628 32004 40638
rect 31500 40626 32004 40628
rect 31500 40574 31950 40626
rect 32002 40574 32004 40626
rect 31500 40572 32004 40574
rect 31948 40562 32004 40572
rect 31388 40350 31390 40402
rect 31442 40350 31444 40402
rect 31388 40338 31444 40350
rect 32060 40404 32116 40414
rect 32060 40310 32116 40348
rect 30828 39618 30884 39676
rect 30828 39566 30830 39618
rect 30882 39566 30884 39618
rect 30828 39554 30884 39566
rect 29484 38110 29486 38162
rect 29538 38110 29540 38162
rect 29484 38098 29540 38110
rect 31612 38164 31668 38174
rect 32172 38164 32228 42252
rect 32284 42242 32340 42252
rect 32396 42700 32564 42756
rect 33068 42754 33124 42812
rect 33068 42702 33070 42754
rect 33122 42702 33124 42754
rect 32284 41972 32340 41982
rect 32396 41972 32452 42700
rect 33068 42690 33124 42702
rect 33180 42756 33236 44940
rect 33404 44940 33572 44996
rect 33180 42690 33236 42700
rect 33292 43540 33348 43550
rect 33292 42754 33348 43484
rect 33404 43538 33460 44940
rect 34412 43988 34468 45276
rect 34636 45218 34692 46508
rect 34748 46452 34804 46462
rect 34748 46002 34804 46396
rect 34748 45950 34750 46002
rect 34802 45950 34804 46002
rect 34748 45938 34804 45950
rect 34636 45166 34638 45218
rect 34690 45166 34692 45218
rect 34636 45154 34692 45166
rect 34748 44884 34804 44894
rect 34748 44790 34804 44828
rect 34860 44882 34916 47404
rect 34972 44996 35028 48860
rect 35980 48850 36036 48860
rect 35644 48804 35700 48814
rect 35644 48710 35700 48748
rect 35868 48802 35924 48814
rect 35868 48750 35870 48802
rect 35922 48750 35924 48802
rect 34972 44930 35028 44940
rect 35084 48692 35140 48702
rect 35084 46676 35140 48636
rect 35868 48468 35924 48750
rect 35868 48402 35924 48412
rect 38220 48242 38276 48254
rect 38220 48190 38222 48242
rect 38274 48190 38276 48242
rect 36876 48130 36932 48142
rect 36876 48078 36878 48130
rect 36930 48078 36932 48130
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 36092 47684 36148 47694
rect 36092 46786 36148 47628
rect 36876 47124 36932 48078
rect 36876 47058 36932 47068
rect 36092 46734 36094 46786
rect 36146 46734 36148 46786
rect 36092 46722 36148 46734
rect 35308 46676 35364 46686
rect 35084 46674 35364 46676
rect 35084 46622 35310 46674
rect 35362 46622 35364 46674
rect 35084 46620 35364 46622
rect 35084 45108 35140 46620
rect 35308 46610 35364 46620
rect 38220 46562 38276 48190
rect 38220 46510 38222 46562
rect 38274 46510 38276 46562
rect 38220 46498 38276 46510
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 36428 45890 36484 45902
rect 36428 45838 36430 45890
rect 36482 45838 36484 45890
rect 35308 45108 35364 45118
rect 35084 45106 35364 45108
rect 35084 45054 35310 45106
rect 35362 45054 35364 45106
rect 35084 45052 35364 45054
rect 34860 44830 34862 44882
rect 34914 44830 34916 44882
rect 34300 43932 34468 43988
rect 33404 43486 33406 43538
rect 33458 43486 33460 43538
rect 33404 43474 33460 43486
rect 33516 43650 33572 43662
rect 33516 43598 33518 43650
rect 33570 43598 33572 43650
rect 33292 42702 33294 42754
rect 33346 42702 33348 42754
rect 33292 42690 33348 42702
rect 33404 42756 33460 42766
rect 33404 42662 33460 42700
rect 32844 42642 32900 42654
rect 32844 42590 32846 42642
rect 32898 42590 32900 42642
rect 32508 42532 32564 42542
rect 32508 42530 32788 42532
rect 32508 42478 32510 42530
rect 32562 42478 32788 42530
rect 32508 42476 32788 42478
rect 32508 42466 32564 42476
rect 32284 41970 32452 41972
rect 32284 41918 32286 41970
rect 32338 41918 32452 41970
rect 32284 41916 32452 41918
rect 32284 41906 32340 41916
rect 32396 41748 32452 41916
rect 32396 41682 32452 41692
rect 32620 42308 32676 42318
rect 32620 41186 32676 42252
rect 32620 41134 32622 41186
rect 32674 41134 32676 41186
rect 32620 41122 32676 41134
rect 32732 42196 32788 42476
rect 32844 42420 32900 42590
rect 32844 42354 32900 42364
rect 32956 42644 33012 42654
rect 32956 42308 33012 42588
rect 33180 42532 33236 42542
rect 33180 42438 33236 42476
rect 33292 42420 33348 42430
rect 32956 42252 33236 42308
rect 32732 41074 32788 42140
rect 32956 41970 33012 41982
rect 32956 41918 32958 41970
rect 33010 41918 33012 41970
rect 32956 41860 33012 41918
rect 33180 41972 33236 42252
rect 33292 42196 33348 42364
rect 33516 42196 33572 43598
rect 33964 43540 34020 43550
rect 33292 42194 33572 42196
rect 33292 42142 33294 42194
rect 33346 42142 33572 42194
rect 33292 42140 33572 42142
rect 33740 43426 33796 43438
rect 33740 43374 33742 43426
rect 33794 43374 33796 43426
rect 33292 42130 33348 42140
rect 33292 41972 33348 41982
rect 33180 41970 33348 41972
rect 33180 41918 33294 41970
rect 33346 41918 33348 41970
rect 33180 41916 33348 41918
rect 33292 41906 33348 41916
rect 33516 41972 33572 41982
rect 32956 41794 33012 41804
rect 33180 41748 33236 41758
rect 33180 41186 33236 41692
rect 33180 41134 33182 41186
rect 33234 41134 33236 41186
rect 33180 41122 33236 41134
rect 32732 41022 32734 41074
rect 32786 41022 32788 41074
rect 32732 41010 32788 41022
rect 33516 41076 33572 41916
rect 33628 41970 33684 41982
rect 33628 41918 33630 41970
rect 33682 41918 33684 41970
rect 33628 41748 33684 41918
rect 33740 41860 33796 43374
rect 33964 41972 34020 43484
rect 33964 41906 34020 41916
rect 34076 42532 34132 42542
rect 33740 41794 33796 41804
rect 33628 41682 33684 41692
rect 33516 41074 33908 41076
rect 33516 41022 33518 41074
rect 33570 41022 33908 41074
rect 33516 41020 33908 41022
rect 33516 41010 33572 41020
rect 32956 40964 33012 40974
rect 32956 40870 33012 40908
rect 32508 40852 32564 40862
rect 32396 40740 32452 40750
rect 32396 40626 32452 40684
rect 32396 40574 32398 40626
rect 32450 40574 32452 40626
rect 32396 40562 32452 40574
rect 32508 40514 32564 40796
rect 32508 40462 32510 40514
rect 32562 40462 32564 40514
rect 32508 40450 32564 40462
rect 33852 40514 33908 41020
rect 33852 40462 33854 40514
rect 33906 40462 33908 40514
rect 33852 40450 33908 40462
rect 33180 40402 33236 40414
rect 33180 40350 33182 40402
rect 33234 40350 33236 40402
rect 33180 39732 33236 40350
rect 33180 39730 33460 39732
rect 33180 39678 33182 39730
rect 33234 39678 33460 39730
rect 33180 39676 33460 39678
rect 33180 39666 33236 39676
rect 33404 38834 33460 39676
rect 34076 38948 34132 42476
rect 34300 42196 34356 43932
rect 34412 43764 34468 43774
rect 34860 43764 34916 44830
rect 35084 44436 35140 45052
rect 35308 45042 35364 45052
rect 36092 44994 36148 45006
rect 36092 44942 36094 44994
rect 36146 44942 36148 44994
rect 36092 44884 36148 44942
rect 36428 44996 36484 45838
rect 36428 44930 36484 44940
rect 38220 44996 38276 45006
rect 38220 44902 38276 44940
rect 36092 44818 36148 44828
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 35084 44434 35364 44436
rect 35084 44382 35086 44434
rect 35138 44382 35364 44434
rect 35084 44380 35364 44382
rect 35084 44370 35140 44380
rect 34412 43762 34916 43764
rect 34412 43710 34414 43762
rect 34466 43710 34916 43762
rect 34412 43708 34916 43710
rect 34412 43698 34468 43708
rect 35308 43540 35364 44380
rect 35308 43538 35588 43540
rect 35308 43486 35310 43538
rect 35362 43486 35588 43538
rect 35308 43484 35588 43486
rect 35308 43474 35364 43484
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 34748 42756 34804 42766
rect 34412 42196 34468 42206
rect 34636 42196 34692 42206
rect 34300 42194 34468 42196
rect 34300 42142 34414 42194
rect 34466 42142 34468 42194
rect 34300 42140 34468 42142
rect 34412 42130 34468 42140
rect 34524 42140 34636 42196
rect 34188 41970 34244 41982
rect 34188 41918 34190 41970
rect 34242 41918 34244 41970
rect 34188 40964 34244 41918
rect 34524 41970 34580 42140
rect 34636 42130 34692 42140
rect 34524 41918 34526 41970
rect 34578 41918 34580 41970
rect 34524 41906 34580 41918
rect 34636 41972 34692 41982
rect 34636 41878 34692 41916
rect 34748 41970 34804 42700
rect 35420 42532 35476 42542
rect 35420 42438 35476 42476
rect 34748 41918 34750 41970
rect 34802 41918 34804 41970
rect 34748 41906 34804 41918
rect 35420 41972 35476 41982
rect 35532 41972 35588 43484
rect 36092 43426 36148 43438
rect 36092 43374 36094 43426
rect 36146 43374 36148 43426
rect 36092 42196 36148 43374
rect 38220 43426 38276 43438
rect 38220 43374 38222 43426
rect 38274 43374 38276 43426
rect 36428 42754 36484 42766
rect 36428 42702 36430 42754
rect 36482 42702 36484 42754
rect 36092 42130 36148 42140
rect 36316 42308 36372 42318
rect 35420 41970 35588 41972
rect 35420 41918 35422 41970
rect 35474 41918 35588 41970
rect 35420 41916 35588 41918
rect 35420 41906 35476 41916
rect 36092 41860 36148 41870
rect 36092 41766 36148 41804
rect 34972 41748 35028 41758
rect 34972 41410 35028 41692
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 34972 41358 34974 41410
rect 35026 41358 35028 41410
rect 34972 41346 35028 41358
rect 36316 41186 36372 42252
rect 36428 41860 36484 42702
rect 38220 42308 38276 43374
rect 38220 42242 38276 42252
rect 36428 41794 36484 41804
rect 38220 41860 38276 41870
rect 38220 41766 38276 41804
rect 36316 41134 36318 41186
rect 36370 41134 36372 41186
rect 36316 41122 36372 41134
rect 34188 40898 34244 40908
rect 35980 40404 36036 40414
rect 35980 40290 36036 40348
rect 35980 40238 35982 40290
rect 36034 40238 36036 40290
rect 35980 40226 36036 40238
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 34972 39060 35028 39070
rect 34188 38948 34244 38958
rect 34076 38946 34244 38948
rect 34076 38894 34190 38946
rect 34242 38894 34244 38946
rect 34076 38892 34244 38894
rect 34188 38882 34244 38892
rect 33404 38782 33406 38834
rect 33458 38782 33460 38834
rect 31612 38162 32228 38164
rect 31612 38110 31614 38162
rect 31666 38110 32228 38162
rect 31612 38108 32228 38110
rect 32396 38612 32452 38622
rect 32396 38164 32452 38556
rect 33404 38612 33460 38782
rect 33404 38546 33460 38556
rect 34972 38274 35028 39004
rect 36316 38722 36372 38734
rect 36316 38670 36318 38722
rect 36370 38670 36372 38722
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 34972 38222 34974 38274
rect 35026 38222 35028 38274
rect 34972 38210 35028 38222
rect 31612 38098 31668 38108
rect 32396 38050 32452 38108
rect 32396 37998 32398 38050
rect 32450 37998 32452 38050
rect 32396 37986 32452 37998
rect 36316 38050 36372 38670
rect 36316 37998 36318 38050
rect 36370 37998 36372 38050
rect 36316 37986 36372 37998
rect 28476 37438 28478 37490
rect 28530 37438 28532 37490
rect 28476 37426 28532 37438
rect 28028 37380 28084 37390
rect 27916 37378 28084 37380
rect 27916 37326 28030 37378
rect 28082 37326 28084 37378
rect 27916 37324 28084 37326
rect 28028 37314 28084 37324
rect 27580 36484 27636 36494
rect 27692 36484 27748 36988
rect 28924 37154 28980 37166
rect 28924 37102 28926 37154
rect 28978 37102 28980 37154
rect 27580 36482 28196 36484
rect 27580 36430 27582 36482
rect 27634 36430 28196 36482
rect 27580 36428 28196 36430
rect 27580 36418 27636 36428
rect 28028 36260 28084 36270
rect 27468 36204 27748 36260
rect 27356 36194 27412 36204
rect 27692 35810 27748 36204
rect 28028 36166 28084 36204
rect 27692 35758 27694 35810
rect 27746 35758 27748 35810
rect 27692 35746 27748 35758
rect 27244 33394 27300 33404
rect 27468 33124 27524 33134
rect 27468 32674 27524 33068
rect 27468 32622 27470 32674
rect 27522 32622 27524 32674
rect 27468 32610 27524 32622
rect 28140 32564 28196 36428
rect 28924 36260 28980 37102
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 38220 36372 38276 36382
rect 38220 36278 38276 36316
rect 28924 36194 28980 36204
rect 29820 36260 29876 36270
rect 29820 35586 29876 36204
rect 29820 35534 29822 35586
rect 29874 35534 29876 35586
rect 29820 35522 29876 35534
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 28140 32470 28196 32508
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 27020 30930 27076 30940
rect 38220 31106 38276 31118
rect 38220 31054 38222 31106
rect 38274 31054 38276 31106
rect 25564 30830 25566 30882
rect 25618 30830 25620 30882
rect 25564 30818 25620 30830
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 23212 30258 23268 30268
rect 24220 30324 24276 30334
rect 24220 30230 24276 30268
rect 38220 30324 38276 31054
rect 38220 30258 38276 30268
rect 21308 30158 21310 30210
rect 21362 30158 21364 30210
rect 21308 30146 21364 30158
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 38220 23266 38276 23278
rect 38220 23214 38222 23266
rect 38274 23214 38276 23266
rect 38220 22932 38276 23214
rect 38220 22866 38276 22876
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 2940 3332 2996 3342
rect 2716 3330 2996 3332
rect 2716 3278 2942 3330
rect 2994 3278 2996 3330
rect 2716 3276 2996 3278
rect 2716 800 2772 3276
rect 2940 3266 2996 3276
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 2688 0 2800 800
<< via2 >>
rect 4476 96458 4532 96460
rect 4476 96406 4478 96458
rect 4478 96406 4530 96458
rect 4530 96406 4532 96458
rect 4476 96404 4532 96406
rect 4580 96458 4636 96460
rect 4580 96406 4582 96458
rect 4582 96406 4634 96458
rect 4634 96406 4636 96458
rect 4580 96404 4636 96406
rect 4684 96458 4740 96460
rect 4684 96406 4686 96458
rect 4686 96406 4738 96458
rect 4738 96406 4740 96458
rect 4684 96404 4740 96406
rect 35196 96458 35252 96460
rect 35196 96406 35198 96458
rect 35198 96406 35250 96458
rect 35250 96406 35252 96458
rect 35196 96404 35252 96406
rect 35300 96458 35356 96460
rect 35300 96406 35302 96458
rect 35302 96406 35354 96458
rect 35354 96406 35356 96458
rect 35300 96404 35356 96406
rect 35404 96458 35460 96460
rect 35404 96406 35406 96458
rect 35406 96406 35458 96458
rect 35458 96406 35460 96458
rect 35404 96404 35460 96406
rect 19836 95674 19892 95676
rect 19836 95622 19838 95674
rect 19838 95622 19890 95674
rect 19890 95622 19892 95674
rect 19836 95620 19892 95622
rect 19940 95674 19996 95676
rect 19940 95622 19942 95674
rect 19942 95622 19994 95674
rect 19994 95622 19996 95674
rect 19940 95620 19996 95622
rect 20044 95674 20100 95676
rect 20044 95622 20046 95674
rect 20046 95622 20098 95674
rect 20098 95622 20100 95674
rect 20044 95620 20100 95622
rect 4476 94890 4532 94892
rect 4476 94838 4478 94890
rect 4478 94838 4530 94890
rect 4530 94838 4532 94890
rect 4476 94836 4532 94838
rect 4580 94890 4636 94892
rect 4580 94838 4582 94890
rect 4582 94838 4634 94890
rect 4634 94838 4636 94890
rect 4580 94836 4636 94838
rect 4684 94890 4740 94892
rect 4684 94838 4686 94890
rect 4686 94838 4738 94890
rect 4738 94838 4740 94890
rect 4684 94836 4740 94838
rect 35196 94890 35252 94892
rect 35196 94838 35198 94890
rect 35198 94838 35250 94890
rect 35250 94838 35252 94890
rect 35196 94836 35252 94838
rect 35300 94890 35356 94892
rect 35300 94838 35302 94890
rect 35302 94838 35354 94890
rect 35354 94838 35356 94890
rect 35300 94836 35356 94838
rect 35404 94890 35460 94892
rect 35404 94838 35406 94890
rect 35406 94838 35458 94890
rect 35458 94838 35460 94890
rect 35404 94836 35460 94838
rect 19836 94106 19892 94108
rect 19836 94054 19838 94106
rect 19838 94054 19890 94106
rect 19890 94054 19892 94106
rect 19836 94052 19892 94054
rect 19940 94106 19996 94108
rect 19940 94054 19942 94106
rect 19942 94054 19994 94106
rect 19994 94054 19996 94106
rect 19940 94052 19996 94054
rect 20044 94106 20100 94108
rect 20044 94054 20046 94106
rect 20046 94054 20098 94106
rect 20098 94054 20100 94106
rect 20044 94052 20100 94054
rect 4476 93322 4532 93324
rect 4476 93270 4478 93322
rect 4478 93270 4530 93322
rect 4530 93270 4532 93322
rect 4476 93268 4532 93270
rect 4580 93322 4636 93324
rect 4580 93270 4582 93322
rect 4582 93270 4634 93322
rect 4634 93270 4636 93322
rect 4580 93268 4636 93270
rect 4684 93322 4740 93324
rect 4684 93270 4686 93322
rect 4686 93270 4738 93322
rect 4738 93270 4740 93322
rect 4684 93268 4740 93270
rect 35196 93322 35252 93324
rect 35196 93270 35198 93322
rect 35198 93270 35250 93322
rect 35250 93270 35252 93322
rect 35196 93268 35252 93270
rect 35300 93322 35356 93324
rect 35300 93270 35302 93322
rect 35302 93270 35354 93322
rect 35354 93270 35356 93322
rect 35300 93268 35356 93270
rect 35404 93322 35460 93324
rect 35404 93270 35406 93322
rect 35406 93270 35458 93322
rect 35458 93270 35460 93322
rect 35404 93268 35460 93270
rect 19836 92538 19892 92540
rect 19836 92486 19838 92538
rect 19838 92486 19890 92538
rect 19890 92486 19892 92538
rect 19836 92484 19892 92486
rect 19940 92538 19996 92540
rect 19940 92486 19942 92538
rect 19942 92486 19994 92538
rect 19994 92486 19996 92538
rect 19940 92484 19996 92486
rect 20044 92538 20100 92540
rect 20044 92486 20046 92538
rect 20046 92486 20098 92538
rect 20098 92486 20100 92538
rect 20044 92484 20100 92486
rect 4476 91754 4532 91756
rect 4476 91702 4478 91754
rect 4478 91702 4530 91754
rect 4530 91702 4532 91754
rect 4476 91700 4532 91702
rect 4580 91754 4636 91756
rect 4580 91702 4582 91754
rect 4582 91702 4634 91754
rect 4634 91702 4636 91754
rect 4580 91700 4636 91702
rect 4684 91754 4740 91756
rect 4684 91702 4686 91754
rect 4686 91702 4738 91754
rect 4738 91702 4740 91754
rect 4684 91700 4740 91702
rect 35196 91754 35252 91756
rect 35196 91702 35198 91754
rect 35198 91702 35250 91754
rect 35250 91702 35252 91754
rect 35196 91700 35252 91702
rect 35300 91754 35356 91756
rect 35300 91702 35302 91754
rect 35302 91702 35354 91754
rect 35354 91702 35356 91754
rect 35300 91700 35356 91702
rect 35404 91754 35460 91756
rect 35404 91702 35406 91754
rect 35406 91702 35458 91754
rect 35458 91702 35460 91754
rect 35404 91700 35460 91702
rect 19836 90970 19892 90972
rect 19836 90918 19838 90970
rect 19838 90918 19890 90970
rect 19890 90918 19892 90970
rect 19836 90916 19892 90918
rect 19940 90970 19996 90972
rect 19940 90918 19942 90970
rect 19942 90918 19994 90970
rect 19994 90918 19996 90970
rect 19940 90916 19996 90918
rect 20044 90970 20100 90972
rect 20044 90918 20046 90970
rect 20046 90918 20098 90970
rect 20098 90918 20100 90970
rect 20044 90916 20100 90918
rect 4476 90186 4532 90188
rect 4476 90134 4478 90186
rect 4478 90134 4530 90186
rect 4530 90134 4532 90186
rect 4476 90132 4532 90134
rect 4580 90186 4636 90188
rect 4580 90134 4582 90186
rect 4582 90134 4634 90186
rect 4634 90134 4636 90186
rect 4580 90132 4636 90134
rect 4684 90186 4740 90188
rect 4684 90134 4686 90186
rect 4686 90134 4738 90186
rect 4738 90134 4740 90186
rect 4684 90132 4740 90134
rect 35196 90186 35252 90188
rect 35196 90134 35198 90186
rect 35198 90134 35250 90186
rect 35250 90134 35252 90186
rect 35196 90132 35252 90134
rect 35300 90186 35356 90188
rect 35300 90134 35302 90186
rect 35302 90134 35354 90186
rect 35354 90134 35356 90186
rect 35300 90132 35356 90134
rect 35404 90186 35460 90188
rect 35404 90134 35406 90186
rect 35406 90134 35458 90186
rect 35458 90134 35460 90186
rect 35404 90132 35460 90134
rect 19836 89402 19892 89404
rect 19836 89350 19838 89402
rect 19838 89350 19890 89402
rect 19890 89350 19892 89402
rect 19836 89348 19892 89350
rect 19940 89402 19996 89404
rect 19940 89350 19942 89402
rect 19942 89350 19994 89402
rect 19994 89350 19996 89402
rect 19940 89348 19996 89350
rect 20044 89402 20100 89404
rect 20044 89350 20046 89402
rect 20046 89350 20098 89402
rect 20098 89350 20100 89402
rect 20044 89348 20100 89350
rect 4476 88618 4532 88620
rect 4476 88566 4478 88618
rect 4478 88566 4530 88618
rect 4530 88566 4532 88618
rect 4476 88564 4532 88566
rect 4580 88618 4636 88620
rect 4580 88566 4582 88618
rect 4582 88566 4634 88618
rect 4634 88566 4636 88618
rect 4580 88564 4636 88566
rect 4684 88618 4740 88620
rect 4684 88566 4686 88618
rect 4686 88566 4738 88618
rect 4738 88566 4740 88618
rect 4684 88564 4740 88566
rect 35196 88618 35252 88620
rect 35196 88566 35198 88618
rect 35198 88566 35250 88618
rect 35250 88566 35252 88618
rect 35196 88564 35252 88566
rect 35300 88618 35356 88620
rect 35300 88566 35302 88618
rect 35302 88566 35354 88618
rect 35354 88566 35356 88618
rect 35300 88564 35356 88566
rect 35404 88618 35460 88620
rect 35404 88566 35406 88618
rect 35406 88566 35458 88618
rect 35458 88566 35460 88618
rect 35404 88564 35460 88566
rect 19836 87834 19892 87836
rect 19836 87782 19838 87834
rect 19838 87782 19890 87834
rect 19890 87782 19892 87834
rect 19836 87780 19892 87782
rect 19940 87834 19996 87836
rect 19940 87782 19942 87834
rect 19942 87782 19994 87834
rect 19994 87782 19996 87834
rect 19940 87780 19996 87782
rect 20044 87834 20100 87836
rect 20044 87782 20046 87834
rect 20046 87782 20098 87834
rect 20098 87782 20100 87834
rect 20044 87780 20100 87782
rect 4476 87050 4532 87052
rect 4476 86998 4478 87050
rect 4478 86998 4530 87050
rect 4530 86998 4532 87050
rect 4476 86996 4532 86998
rect 4580 87050 4636 87052
rect 4580 86998 4582 87050
rect 4582 86998 4634 87050
rect 4634 86998 4636 87050
rect 4580 86996 4636 86998
rect 4684 87050 4740 87052
rect 4684 86998 4686 87050
rect 4686 86998 4738 87050
rect 4738 86998 4740 87050
rect 4684 86996 4740 86998
rect 35196 87050 35252 87052
rect 35196 86998 35198 87050
rect 35198 86998 35250 87050
rect 35250 86998 35252 87050
rect 35196 86996 35252 86998
rect 35300 87050 35356 87052
rect 35300 86998 35302 87050
rect 35302 86998 35354 87050
rect 35354 86998 35356 87050
rect 35300 86996 35356 86998
rect 35404 87050 35460 87052
rect 35404 86998 35406 87050
rect 35406 86998 35458 87050
rect 35458 86998 35460 87050
rect 35404 86996 35460 86998
rect 19836 86266 19892 86268
rect 19836 86214 19838 86266
rect 19838 86214 19890 86266
rect 19890 86214 19892 86266
rect 19836 86212 19892 86214
rect 19940 86266 19996 86268
rect 19940 86214 19942 86266
rect 19942 86214 19994 86266
rect 19994 86214 19996 86266
rect 19940 86212 19996 86214
rect 20044 86266 20100 86268
rect 20044 86214 20046 86266
rect 20046 86214 20098 86266
rect 20098 86214 20100 86266
rect 20044 86212 20100 86214
rect 4476 85482 4532 85484
rect 4476 85430 4478 85482
rect 4478 85430 4530 85482
rect 4530 85430 4532 85482
rect 4476 85428 4532 85430
rect 4580 85482 4636 85484
rect 4580 85430 4582 85482
rect 4582 85430 4634 85482
rect 4634 85430 4636 85482
rect 4580 85428 4636 85430
rect 4684 85482 4740 85484
rect 4684 85430 4686 85482
rect 4686 85430 4738 85482
rect 4738 85430 4740 85482
rect 4684 85428 4740 85430
rect 35196 85482 35252 85484
rect 35196 85430 35198 85482
rect 35198 85430 35250 85482
rect 35250 85430 35252 85482
rect 35196 85428 35252 85430
rect 35300 85482 35356 85484
rect 35300 85430 35302 85482
rect 35302 85430 35354 85482
rect 35354 85430 35356 85482
rect 35300 85428 35356 85430
rect 35404 85482 35460 85484
rect 35404 85430 35406 85482
rect 35406 85430 35458 85482
rect 35458 85430 35460 85482
rect 35404 85428 35460 85430
rect 19836 84698 19892 84700
rect 19836 84646 19838 84698
rect 19838 84646 19890 84698
rect 19890 84646 19892 84698
rect 19836 84644 19892 84646
rect 19940 84698 19996 84700
rect 19940 84646 19942 84698
rect 19942 84646 19994 84698
rect 19994 84646 19996 84698
rect 19940 84644 19996 84646
rect 20044 84698 20100 84700
rect 20044 84646 20046 84698
rect 20046 84646 20098 84698
rect 20098 84646 20100 84698
rect 20044 84644 20100 84646
rect 4476 83914 4532 83916
rect 4476 83862 4478 83914
rect 4478 83862 4530 83914
rect 4530 83862 4532 83914
rect 4476 83860 4532 83862
rect 4580 83914 4636 83916
rect 4580 83862 4582 83914
rect 4582 83862 4634 83914
rect 4634 83862 4636 83914
rect 4580 83860 4636 83862
rect 4684 83914 4740 83916
rect 4684 83862 4686 83914
rect 4686 83862 4738 83914
rect 4738 83862 4740 83914
rect 4684 83860 4740 83862
rect 35196 83914 35252 83916
rect 35196 83862 35198 83914
rect 35198 83862 35250 83914
rect 35250 83862 35252 83914
rect 35196 83860 35252 83862
rect 35300 83914 35356 83916
rect 35300 83862 35302 83914
rect 35302 83862 35354 83914
rect 35354 83862 35356 83914
rect 35300 83860 35356 83862
rect 35404 83914 35460 83916
rect 35404 83862 35406 83914
rect 35406 83862 35458 83914
rect 35458 83862 35460 83914
rect 35404 83860 35460 83862
rect 19836 83130 19892 83132
rect 19836 83078 19838 83130
rect 19838 83078 19890 83130
rect 19890 83078 19892 83130
rect 19836 83076 19892 83078
rect 19940 83130 19996 83132
rect 19940 83078 19942 83130
rect 19942 83078 19994 83130
rect 19994 83078 19996 83130
rect 19940 83076 19996 83078
rect 20044 83130 20100 83132
rect 20044 83078 20046 83130
rect 20046 83078 20098 83130
rect 20098 83078 20100 83130
rect 20044 83076 20100 83078
rect 4476 82346 4532 82348
rect 4476 82294 4478 82346
rect 4478 82294 4530 82346
rect 4530 82294 4532 82346
rect 4476 82292 4532 82294
rect 4580 82346 4636 82348
rect 4580 82294 4582 82346
rect 4582 82294 4634 82346
rect 4634 82294 4636 82346
rect 4580 82292 4636 82294
rect 4684 82346 4740 82348
rect 4684 82294 4686 82346
rect 4686 82294 4738 82346
rect 4738 82294 4740 82346
rect 4684 82292 4740 82294
rect 35196 82346 35252 82348
rect 35196 82294 35198 82346
rect 35198 82294 35250 82346
rect 35250 82294 35252 82346
rect 35196 82292 35252 82294
rect 35300 82346 35356 82348
rect 35300 82294 35302 82346
rect 35302 82294 35354 82346
rect 35354 82294 35356 82346
rect 35300 82292 35356 82294
rect 35404 82346 35460 82348
rect 35404 82294 35406 82346
rect 35406 82294 35458 82346
rect 35458 82294 35460 82346
rect 35404 82292 35460 82294
rect 19836 81562 19892 81564
rect 19836 81510 19838 81562
rect 19838 81510 19890 81562
rect 19890 81510 19892 81562
rect 19836 81508 19892 81510
rect 19940 81562 19996 81564
rect 19940 81510 19942 81562
rect 19942 81510 19994 81562
rect 19994 81510 19996 81562
rect 19940 81508 19996 81510
rect 20044 81562 20100 81564
rect 20044 81510 20046 81562
rect 20046 81510 20098 81562
rect 20098 81510 20100 81562
rect 20044 81508 20100 81510
rect 4476 80778 4532 80780
rect 4476 80726 4478 80778
rect 4478 80726 4530 80778
rect 4530 80726 4532 80778
rect 4476 80724 4532 80726
rect 4580 80778 4636 80780
rect 4580 80726 4582 80778
rect 4582 80726 4634 80778
rect 4634 80726 4636 80778
rect 4580 80724 4636 80726
rect 4684 80778 4740 80780
rect 4684 80726 4686 80778
rect 4686 80726 4738 80778
rect 4738 80726 4740 80778
rect 4684 80724 4740 80726
rect 35196 80778 35252 80780
rect 35196 80726 35198 80778
rect 35198 80726 35250 80778
rect 35250 80726 35252 80778
rect 35196 80724 35252 80726
rect 35300 80778 35356 80780
rect 35300 80726 35302 80778
rect 35302 80726 35354 80778
rect 35354 80726 35356 80778
rect 35300 80724 35356 80726
rect 35404 80778 35460 80780
rect 35404 80726 35406 80778
rect 35406 80726 35458 80778
rect 35458 80726 35460 80778
rect 35404 80724 35460 80726
rect 19836 79994 19892 79996
rect 19836 79942 19838 79994
rect 19838 79942 19890 79994
rect 19890 79942 19892 79994
rect 19836 79940 19892 79942
rect 19940 79994 19996 79996
rect 19940 79942 19942 79994
rect 19942 79942 19994 79994
rect 19994 79942 19996 79994
rect 19940 79940 19996 79942
rect 20044 79994 20100 79996
rect 20044 79942 20046 79994
rect 20046 79942 20098 79994
rect 20098 79942 20100 79994
rect 20044 79940 20100 79942
rect 4476 79210 4532 79212
rect 4476 79158 4478 79210
rect 4478 79158 4530 79210
rect 4530 79158 4532 79210
rect 4476 79156 4532 79158
rect 4580 79210 4636 79212
rect 4580 79158 4582 79210
rect 4582 79158 4634 79210
rect 4634 79158 4636 79210
rect 4580 79156 4636 79158
rect 4684 79210 4740 79212
rect 4684 79158 4686 79210
rect 4686 79158 4738 79210
rect 4738 79158 4740 79210
rect 4684 79156 4740 79158
rect 35196 79210 35252 79212
rect 35196 79158 35198 79210
rect 35198 79158 35250 79210
rect 35250 79158 35252 79210
rect 35196 79156 35252 79158
rect 35300 79210 35356 79212
rect 35300 79158 35302 79210
rect 35302 79158 35354 79210
rect 35354 79158 35356 79210
rect 35300 79156 35356 79158
rect 35404 79210 35460 79212
rect 35404 79158 35406 79210
rect 35406 79158 35458 79210
rect 35458 79158 35460 79210
rect 35404 79156 35460 79158
rect 19836 78426 19892 78428
rect 19836 78374 19838 78426
rect 19838 78374 19890 78426
rect 19890 78374 19892 78426
rect 19836 78372 19892 78374
rect 19940 78426 19996 78428
rect 19940 78374 19942 78426
rect 19942 78374 19994 78426
rect 19994 78374 19996 78426
rect 19940 78372 19996 78374
rect 20044 78426 20100 78428
rect 20044 78374 20046 78426
rect 20046 78374 20098 78426
rect 20098 78374 20100 78426
rect 20044 78372 20100 78374
rect 4476 77642 4532 77644
rect 4476 77590 4478 77642
rect 4478 77590 4530 77642
rect 4530 77590 4532 77642
rect 4476 77588 4532 77590
rect 4580 77642 4636 77644
rect 4580 77590 4582 77642
rect 4582 77590 4634 77642
rect 4634 77590 4636 77642
rect 4580 77588 4636 77590
rect 4684 77642 4740 77644
rect 4684 77590 4686 77642
rect 4686 77590 4738 77642
rect 4738 77590 4740 77642
rect 4684 77588 4740 77590
rect 35196 77642 35252 77644
rect 35196 77590 35198 77642
rect 35198 77590 35250 77642
rect 35250 77590 35252 77642
rect 35196 77588 35252 77590
rect 35300 77642 35356 77644
rect 35300 77590 35302 77642
rect 35302 77590 35354 77642
rect 35354 77590 35356 77642
rect 35300 77588 35356 77590
rect 35404 77642 35460 77644
rect 35404 77590 35406 77642
rect 35406 77590 35458 77642
rect 35458 77590 35460 77642
rect 35404 77588 35460 77590
rect 19836 76858 19892 76860
rect 19836 76806 19838 76858
rect 19838 76806 19890 76858
rect 19890 76806 19892 76858
rect 19836 76804 19892 76806
rect 19940 76858 19996 76860
rect 19940 76806 19942 76858
rect 19942 76806 19994 76858
rect 19994 76806 19996 76858
rect 19940 76804 19996 76806
rect 20044 76858 20100 76860
rect 20044 76806 20046 76858
rect 20046 76806 20098 76858
rect 20098 76806 20100 76858
rect 20044 76804 20100 76806
rect 4476 76074 4532 76076
rect 4476 76022 4478 76074
rect 4478 76022 4530 76074
rect 4530 76022 4532 76074
rect 4476 76020 4532 76022
rect 4580 76074 4636 76076
rect 4580 76022 4582 76074
rect 4582 76022 4634 76074
rect 4634 76022 4636 76074
rect 4580 76020 4636 76022
rect 4684 76074 4740 76076
rect 4684 76022 4686 76074
rect 4686 76022 4738 76074
rect 4738 76022 4740 76074
rect 4684 76020 4740 76022
rect 35196 76074 35252 76076
rect 35196 76022 35198 76074
rect 35198 76022 35250 76074
rect 35250 76022 35252 76074
rect 35196 76020 35252 76022
rect 35300 76074 35356 76076
rect 35300 76022 35302 76074
rect 35302 76022 35354 76074
rect 35354 76022 35356 76074
rect 35300 76020 35356 76022
rect 35404 76074 35460 76076
rect 35404 76022 35406 76074
rect 35406 76022 35458 76074
rect 35458 76022 35460 76074
rect 35404 76020 35460 76022
rect 19836 75290 19892 75292
rect 19836 75238 19838 75290
rect 19838 75238 19890 75290
rect 19890 75238 19892 75290
rect 19836 75236 19892 75238
rect 19940 75290 19996 75292
rect 19940 75238 19942 75290
rect 19942 75238 19994 75290
rect 19994 75238 19996 75290
rect 19940 75236 19996 75238
rect 20044 75290 20100 75292
rect 20044 75238 20046 75290
rect 20046 75238 20098 75290
rect 20098 75238 20100 75290
rect 20044 75236 20100 75238
rect 4476 74506 4532 74508
rect 4476 74454 4478 74506
rect 4478 74454 4530 74506
rect 4530 74454 4532 74506
rect 4476 74452 4532 74454
rect 4580 74506 4636 74508
rect 4580 74454 4582 74506
rect 4582 74454 4634 74506
rect 4634 74454 4636 74506
rect 4580 74452 4636 74454
rect 4684 74506 4740 74508
rect 4684 74454 4686 74506
rect 4686 74454 4738 74506
rect 4738 74454 4740 74506
rect 4684 74452 4740 74454
rect 35196 74506 35252 74508
rect 35196 74454 35198 74506
rect 35198 74454 35250 74506
rect 35250 74454 35252 74506
rect 35196 74452 35252 74454
rect 35300 74506 35356 74508
rect 35300 74454 35302 74506
rect 35302 74454 35354 74506
rect 35354 74454 35356 74506
rect 35300 74452 35356 74454
rect 35404 74506 35460 74508
rect 35404 74454 35406 74506
rect 35406 74454 35458 74506
rect 35458 74454 35460 74506
rect 35404 74452 35460 74454
rect 19836 73722 19892 73724
rect 19836 73670 19838 73722
rect 19838 73670 19890 73722
rect 19890 73670 19892 73722
rect 19836 73668 19892 73670
rect 19940 73722 19996 73724
rect 19940 73670 19942 73722
rect 19942 73670 19994 73722
rect 19994 73670 19996 73722
rect 19940 73668 19996 73670
rect 20044 73722 20100 73724
rect 20044 73670 20046 73722
rect 20046 73670 20098 73722
rect 20098 73670 20100 73722
rect 20044 73668 20100 73670
rect 4476 72938 4532 72940
rect 4476 72886 4478 72938
rect 4478 72886 4530 72938
rect 4530 72886 4532 72938
rect 4476 72884 4532 72886
rect 4580 72938 4636 72940
rect 4580 72886 4582 72938
rect 4582 72886 4634 72938
rect 4634 72886 4636 72938
rect 4580 72884 4636 72886
rect 4684 72938 4740 72940
rect 4684 72886 4686 72938
rect 4686 72886 4738 72938
rect 4738 72886 4740 72938
rect 4684 72884 4740 72886
rect 35196 72938 35252 72940
rect 35196 72886 35198 72938
rect 35198 72886 35250 72938
rect 35250 72886 35252 72938
rect 35196 72884 35252 72886
rect 35300 72938 35356 72940
rect 35300 72886 35302 72938
rect 35302 72886 35354 72938
rect 35354 72886 35356 72938
rect 35300 72884 35356 72886
rect 35404 72938 35460 72940
rect 35404 72886 35406 72938
rect 35406 72886 35458 72938
rect 35458 72886 35460 72938
rect 35404 72884 35460 72886
rect 19836 72154 19892 72156
rect 19836 72102 19838 72154
rect 19838 72102 19890 72154
rect 19890 72102 19892 72154
rect 19836 72100 19892 72102
rect 19940 72154 19996 72156
rect 19940 72102 19942 72154
rect 19942 72102 19994 72154
rect 19994 72102 19996 72154
rect 19940 72100 19996 72102
rect 20044 72154 20100 72156
rect 20044 72102 20046 72154
rect 20046 72102 20098 72154
rect 20098 72102 20100 72154
rect 20044 72100 20100 72102
rect 4476 71370 4532 71372
rect 4476 71318 4478 71370
rect 4478 71318 4530 71370
rect 4530 71318 4532 71370
rect 4476 71316 4532 71318
rect 4580 71370 4636 71372
rect 4580 71318 4582 71370
rect 4582 71318 4634 71370
rect 4634 71318 4636 71370
rect 4580 71316 4636 71318
rect 4684 71370 4740 71372
rect 4684 71318 4686 71370
rect 4686 71318 4738 71370
rect 4738 71318 4740 71370
rect 4684 71316 4740 71318
rect 35196 71370 35252 71372
rect 35196 71318 35198 71370
rect 35198 71318 35250 71370
rect 35250 71318 35252 71370
rect 35196 71316 35252 71318
rect 35300 71370 35356 71372
rect 35300 71318 35302 71370
rect 35302 71318 35354 71370
rect 35354 71318 35356 71370
rect 35300 71316 35356 71318
rect 35404 71370 35460 71372
rect 35404 71318 35406 71370
rect 35406 71318 35458 71370
rect 35458 71318 35460 71370
rect 35404 71316 35460 71318
rect 19836 70586 19892 70588
rect 19836 70534 19838 70586
rect 19838 70534 19890 70586
rect 19890 70534 19892 70586
rect 19836 70532 19892 70534
rect 19940 70586 19996 70588
rect 19940 70534 19942 70586
rect 19942 70534 19994 70586
rect 19994 70534 19996 70586
rect 19940 70532 19996 70534
rect 20044 70586 20100 70588
rect 20044 70534 20046 70586
rect 20046 70534 20098 70586
rect 20098 70534 20100 70586
rect 20044 70532 20100 70534
rect 4476 69802 4532 69804
rect 4476 69750 4478 69802
rect 4478 69750 4530 69802
rect 4530 69750 4532 69802
rect 4476 69748 4532 69750
rect 4580 69802 4636 69804
rect 4580 69750 4582 69802
rect 4582 69750 4634 69802
rect 4634 69750 4636 69802
rect 4580 69748 4636 69750
rect 4684 69802 4740 69804
rect 4684 69750 4686 69802
rect 4686 69750 4738 69802
rect 4738 69750 4740 69802
rect 4684 69748 4740 69750
rect 13020 69356 13076 69412
rect 2044 68738 2100 68740
rect 2044 68686 2046 68738
rect 2046 68686 2098 68738
rect 2098 68686 2100 68738
rect 2044 68684 2100 68686
rect 9660 68738 9716 68740
rect 9660 68686 9662 68738
rect 9662 68686 9714 68738
rect 9714 68686 9716 68738
rect 9660 68684 9716 68686
rect 8316 68572 8372 68628
rect 1708 68460 1764 68516
rect 2492 68514 2548 68516
rect 2492 68462 2494 68514
rect 2494 68462 2546 68514
rect 2546 68462 2548 68514
rect 2492 68460 2548 68462
rect 4476 68234 4532 68236
rect 4476 68182 4478 68234
rect 4478 68182 4530 68234
rect 4530 68182 4532 68234
rect 4476 68180 4532 68182
rect 4580 68234 4636 68236
rect 4580 68182 4582 68234
rect 4582 68182 4634 68234
rect 4634 68182 4636 68234
rect 4580 68180 4636 68182
rect 4684 68234 4740 68236
rect 4684 68182 4686 68234
rect 4686 68182 4738 68234
rect 4738 68182 4740 68234
rect 4684 68180 4740 68182
rect 1708 67900 1764 67956
rect 7644 67954 7700 67956
rect 7644 67902 7646 67954
rect 7646 67902 7698 67954
rect 7698 67902 7700 67954
rect 7644 67900 7700 67902
rect 2044 67340 2100 67396
rect 1708 67228 1764 67284
rect 2492 67228 2548 67284
rect 8204 67340 8260 67396
rect 2044 67170 2100 67172
rect 2044 67118 2046 67170
rect 2046 67118 2098 67170
rect 2098 67118 2100 67170
rect 2044 67116 2100 67118
rect 9772 68572 9828 68628
rect 9772 68402 9828 68404
rect 9772 68350 9774 68402
rect 9774 68350 9826 68402
rect 9826 68350 9828 68402
rect 9772 68348 9828 68350
rect 8764 67900 8820 67956
rect 1708 66556 1764 66612
rect 2492 66556 2548 66612
rect 4476 66666 4532 66668
rect 4476 66614 4478 66666
rect 4478 66614 4530 66666
rect 4530 66614 4532 66666
rect 4476 66612 4532 66614
rect 4580 66666 4636 66668
rect 4580 66614 4582 66666
rect 4582 66614 4634 66666
rect 4634 66614 4636 66666
rect 4580 66612 4636 66614
rect 4684 66666 4740 66668
rect 4684 66614 4686 66666
rect 4686 66614 4738 66666
rect 4738 66614 4740 66666
rect 4684 66612 4740 66614
rect 10108 67676 10164 67732
rect 8652 67004 8708 67060
rect 4476 65098 4532 65100
rect 4476 65046 4478 65098
rect 4478 65046 4530 65098
rect 4530 65046 4532 65098
rect 4476 65044 4532 65046
rect 4580 65098 4636 65100
rect 4580 65046 4582 65098
rect 4582 65046 4634 65098
rect 4634 65046 4636 65098
rect 4580 65044 4636 65046
rect 4684 65098 4740 65100
rect 4684 65046 4686 65098
rect 4686 65046 4738 65098
rect 4738 65046 4740 65098
rect 4684 65044 4740 65046
rect 2380 64594 2436 64596
rect 2380 64542 2382 64594
rect 2382 64542 2434 64594
rect 2434 64542 2436 64594
rect 2380 64540 2436 64542
rect 2716 64594 2772 64596
rect 2716 64542 2718 64594
rect 2718 64542 2770 64594
rect 2770 64542 2772 64594
rect 2716 64540 2772 64542
rect 8652 64594 8708 64596
rect 8652 64542 8654 64594
rect 8654 64542 8706 64594
rect 8706 64542 8708 64594
rect 8652 64540 8708 64542
rect 9884 67116 9940 67172
rect 9436 67058 9492 67060
rect 9436 67006 9438 67058
rect 9438 67006 9490 67058
rect 9490 67006 9492 67058
rect 9436 67004 9492 67006
rect 8876 64764 8932 64820
rect 1820 64428 1876 64484
rect 1820 63868 1876 63924
rect 2044 63756 2100 63812
rect 3164 64482 3220 64484
rect 3164 64430 3166 64482
rect 3166 64430 3218 64482
rect 3218 64430 3220 64482
rect 3164 64428 3220 64430
rect 2156 63308 2212 63364
rect 1708 63196 1764 63252
rect 9436 65548 9492 65604
rect 11788 68348 11844 68404
rect 11452 67730 11508 67732
rect 11452 67678 11454 67730
rect 11454 67678 11506 67730
rect 11506 67678 11508 67730
rect 11452 67676 11508 67678
rect 12348 67730 12404 67732
rect 12348 67678 12350 67730
rect 12350 67678 12402 67730
rect 12402 67678 12404 67730
rect 12348 67676 12404 67678
rect 12908 67730 12964 67732
rect 12908 67678 12910 67730
rect 12910 67678 12962 67730
rect 12962 67678 12964 67730
rect 12908 67676 12964 67678
rect 12796 67618 12852 67620
rect 12796 67566 12798 67618
rect 12798 67566 12850 67618
rect 12850 67566 12852 67618
rect 12796 67564 12852 67566
rect 11228 66444 11284 66500
rect 12572 66444 12628 66500
rect 15260 69410 15316 69412
rect 15260 69358 15262 69410
rect 15262 69358 15314 69410
rect 15314 69358 15316 69410
rect 15260 69356 15316 69358
rect 13244 68514 13300 68516
rect 13244 68462 13246 68514
rect 13246 68462 13298 68514
rect 13298 68462 13300 68514
rect 13244 68460 13300 68462
rect 13580 67618 13636 67620
rect 13580 67566 13582 67618
rect 13582 67566 13634 67618
rect 13634 67566 13636 67618
rect 13580 67564 13636 67566
rect 10892 65548 10948 65604
rect 8988 63980 9044 64036
rect 4476 63530 4532 63532
rect 4476 63478 4478 63530
rect 4478 63478 4530 63530
rect 4530 63478 4532 63530
rect 4476 63476 4532 63478
rect 4580 63530 4636 63532
rect 4580 63478 4582 63530
rect 4582 63478 4634 63530
rect 4634 63478 4636 63530
rect 4580 63476 4636 63478
rect 4684 63530 4740 63532
rect 4684 63478 4686 63530
rect 4686 63478 4738 63530
rect 4738 63478 4740 63530
rect 4684 63476 4740 63478
rect 2492 63196 2548 63252
rect 2044 63026 2100 63028
rect 2044 62974 2046 63026
rect 2046 62974 2098 63026
rect 2098 62974 2100 63026
rect 2044 62972 2100 62974
rect 8876 63026 8932 63028
rect 8876 62974 8878 63026
rect 8878 62974 8930 63026
rect 8930 62974 8932 63026
rect 8876 62972 8932 62974
rect 1708 62524 1764 62580
rect 2492 62524 2548 62580
rect 8092 62578 8148 62580
rect 8092 62526 8094 62578
rect 8094 62526 8146 62578
rect 8146 62526 8148 62578
rect 8092 62524 8148 62526
rect 8988 62524 9044 62580
rect 4476 61962 4532 61964
rect 4476 61910 4478 61962
rect 4478 61910 4530 61962
rect 4530 61910 4532 61962
rect 4476 61908 4532 61910
rect 4580 61962 4636 61964
rect 4580 61910 4582 61962
rect 4582 61910 4634 61962
rect 4634 61910 4636 61962
rect 4580 61908 4636 61910
rect 4684 61962 4740 61964
rect 4684 61910 4686 61962
rect 4686 61910 4738 61962
rect 4738 61910 4740 61962
rect 4684 61908 4740 61910
rect 4476 60394 4532 60396
rect 4476 60342 4478 60394
rect 4478 60342 4530 60394
rect 4530 60342 4532 60394
rect 4476 60340 4532 60342
rect 4580 60394 4636 60396
rect 4580 60342 4582 60394
rect 4582 60342 4634 60394
rect 4634 60342 4636 60394
rect 4580 60340 4636 60342
rect 4684 60394 4740 60396
rect 4684 60342 4686 60394
rect 4686 60342 4738 60394
rect 4738 60342 4740 60394
rect 4684 60340 4740 60342
rect 6076 60396 6132 60452
rect 1708 59890 1764 59892
rect 1708 59838 1710 59890
rect 1710 59838 1762 59890
rect 1762 59838 1764 59890
rect 1708 59836 1764 59838
rect 2492 59890 2548 59892
rect 2492 59838 2494 59890
rect 2494 59838 2546 59890
rect 2546 59838 2548 59890
rect 2492 59836 2548 59838
rect 2044 59778 2100 59780
rect 2044 59726 2046 59778
rect 2046 59726 2098 59778
rect 2098 59726 2100 59778
rect 2044 59724 2100 59726
rect 1708 59164 1764 59220
rect 4476 58826 4532 58828
rect 4476 58774 4478 58826
rect 4478 58774 4530 58826
rect 4530 58774 4532 58826
rect 4476 58772 4532 58774
rect 4580 58826 4636 58828
rect 4580 58774 4582 58826
rect 4582 58774 4634 58826
rect 4634 58774 4636 58826
rect 4580 58772 4636 58774
rect 4684 58826 4740 58828
rect 4684 58774 4686 58826
rect 4686 58774 4738 58826
rect 4738 58774 4740 58826
rect 4684 58772 4740 58774
rect 8204 59218 8260 59220
rect 8204 59166 8206 59218
rect 8206 59166 8258 59218
rect 8258 59166 8260 59218
rect 8204 59164 8260 59166
rect 2044 58210 2100 58212
rect 2044 58158 2046 58210
rect 2046 58158 2098 58210
rect 2098 58158 2100 58210
rect 2044 58156 2100 58158
rect 1708 57820 1764 57876
rect 2492 57820 2548 57876
rect 7756 58156 7812 58212
rect 2044 57762 2100 57764
rect 2044 57710 2046 57762
rect 2046 57710 2098 57762
rect 2098 57710 2100 57762
rect 2044 57708 2100 57710
rect 1708 57148 1764 57204
rect 2492 57148 2548 57204
rect 4476 57258 4532 57260
rect 4476 57206 4478 57258
rect 4478 57206 4530 57258
rect 4530 57206 4532 57258
rect 4476 57204 4532 57206
rect 4580 57258 4636 57260
rect 4580 57206 4582 57258
rect 4582 57206 4634 57258
rect 4634 57206 4636 57258
rect 4580 57204 4636 57206
rect 4684 57258 4740 57260
rect 4684 57206 4686 57258
rect 4686 57206 4738 57258
rect 4738 57206 4740 57258
rect 4684 57204 4740 57206
rect 8876 62242 8932 62244
rect 8876 62190 8878 62242
rect 8878 62190 8930 62242
rect 8930 62190 8932 62242
rect 8876 62188 8932 62190
rect 8764 61740 8820 61796
rect 9212 59724 9268 59780
rect 1708 56476 1764 56532
rect 2044 56306 2100 56308
rect 2044 56254 2046 56306
rect 2046 56254 2098 56306
rect 2098 56254 2100 56306
rect 2044 56252 2100 56254
rect 2492 56476 2548 56532
rect 7420 56252 7476 56308
rect 2156 56140 2212 56196
rect 1708 55804 1764 55860
rect 2492 55804 2548 55860
rect 4476 55690 4532 55692
rect 4476 55638 4478 55690
rect 4478 55638 4530 55690
rect 4530 55638 4532 55690
rect 4476 55636 4532 55638
rect 4580 55690 4636 55692
rect 4580 55638 4582 55690
rect 4582 55638 4634 55690
rect 4634 55638 4636 55690
rect 4580 55636 4636 55638
rect 4684 55690 4740 55692
rect 4684 55638 4686 55690
rect 4686 55638 4738 55690
rect 4738 55638 4740 55690
rect 4684 55636 4740 55638
rect 2044 55244 2100 55300
rect 6636 55970 6692 55972
rect 6636 55918 6638 55970
rect 6638 55918 6690 55970
rect 6690 55918 6692 55970
rect 6636 55916 6692 55918
rect 7644 55692 7700 55748
rect 6300 55468 6356 55524
rect 1708 55186 1764 55188
rect 1708 55134 1710 55186
rect 1710 55134 1762 55186
rect 1762 55134 1764 55186
rect 1708 55132 1764 55134
rect 2492 55186 2548 55188
rect 2492 55134 2494 55186
rect 2494 55134 2546 55186
rect 2546 55134 2548 55186
rect 2492 55132 2548 55134
rect 4476 54122 4532 54124
rect 4476 54070 4478 54122
rect 4478 54070 4530 54122
rect 4530 54070 4532 54122
rect 4476 54068 4532 54070
rect 4580 54122 4636 54124
rect 4580 54070 4582 54122
rect 4582 54070 4634 54122
rect 4634 54070 4636 54122
rect 4580 54068 4636 54070
rect 4684 54122 4740 54124
rect 4684 54070 4686 54122
rect 4686 54070 4738 54122
rect 4738 54070 4740 54122
rect 4684 54068 4740 54070
rect 1708 53116 1764 53172
rect 2044 52108 2100 52164
rect 2492 53116 2548 53172
rect 4476 52554 4532 52556
rect 4476 52502 4478 52554
rect 4478 52502 4530 52554
rect 4530 52502 4532 52554
rect 4476 52500 4532 52502
rect 4580 52554 4636 52556
rect 4580 52502 4582 52554
rect 4582 52502 4634 52554
rect 4634 52502 4636 52554
rect 4580 52500 4636 52502
rect 4684 52554 4740 52556
rect 4684 52502 4686 52554
rect 4686 52502 4738 52554
rect 4738 52502 4740 52554
rect 4684 52500 4740 52502
rect 2156 51996 2212 52052
rect 1708 51772 1764 51828
rect 2492 51772 2548 51828
rect 2044 51490 2100 51492
rect 2044 51438 2046 51490
rect 2046 51438 2098 51490
rect 2098 51438 2100 51490
rect 2044 51436 2100 51438
rect 6972 55186 7028 55188
rect 6972 55134 6974 55186
rect 6974 55134 7026 55186
rect 7026 55134 7028 55186
rect 6972 55132 7028 55134
rect 8092 55132 8148 55188
rect 8204 56028 8260 56084
rect 8316 55356 8372 55412
rect 8540 56140 8596 56196
rect 8652 58156 8708 58212
rect 8652 55244 8708 55300
rect 7868 53676 7924 53732
rect 1708 51100 1764 51156
rect 2492 51100 2548 51156
rect 4476 50986 4532 50988
rect 4476 50934 4478 50986
rect 4478 50934 4530 50986
rect 4530 50934 4532 50986
rect 4476 50932 4532 50934
rect 4580 50986 4636 50988
rect 4580 50934 4582 50986
rect 4582 50934 4634 50986
rect 4634 50934 4636 50986
rect 4580 50932 4636 50934
rect 4684 50986 4740 50988
rect 4684 50934 4686 50986
rect 4686 50934 4738 50986
rect 4738 50934 4740 50986
rect 4684 50932 4740 50934
rect 2716 50540 2772 50596
rect 1708 50482 1764 50484
rect 1708 50430 1710 50482
rect 1710 50430 1762 50482
rect 1762 50430 1764 50482
rect 1708 50428 1764 50430
rect 2044 50370 2100 50372
rect 2044 50318 2046 50370
rect 2046 50318 2098 50370
rect 2098 50318 2100 50370
rect 2044 50316 2100 50318
rect 2044 49922 2100 49924
rect 2044 49870 2046 49922
rect 2046 49870 2098 49922
rect 2098 49870 2100 49922
rect 2044 49868 2100 49870
rect 2492 50428 2548 50484
rect 2380 49756 2436 49812
rect 3164 49756 3220 49812
rect 7756 50482 7812 50484
rect 7756 50430 7758 50482
rect 7758 50430 7810 50482
rect 7810 50430 7812 50482
rect 7756 50428 7812 50430
rect 8652 54460 8708 54516
rect 9100 55804 9156 55860
rect 11340 64764 11396 64820
rect 10108 64316 10164 64372
rect 9996 63868 10052 63924
rect 9436 60396 9492 60452
rect 10220 63980 10276 64036
rect 10892 63922 10948 63924
rect 10892 63870 10894 63922
rect 10894 63870 10946 63922
rect 10946 63870 10948 63922
rect 10892 63868 10948 63870
rect 11452 62524 11508 62580
rect 10220 62412 10276 62468
rect 11004 62412 11060 62468
rect 10332 62242 10388 62244
rect 10332 62190 10334 62242
rect 10334 62190 10386 62242
rect 10386 62190 10388 62242
rect 10332 62188 10388 62190
rect 10108 61740 10164 61796
rect 9548 59388 9604 59444
rect 9660 61292 9716 61348
rect 10444 61458 10500 61460
rect 10444 61406 10446 61458
rect 10446 61406 10498 61458
rect 10498 61406 10500 61458
rect 10444 61404 10500 61406
rect 10332 61346 10388 61348
rect 10332 61294 10334 61346
rect 10334 61294 10386 61346
rect 10386 61294 10388 61346
rect 10332 61292 10388 61294
rect 9436 59218 9492 59220
rect 9436 59166 9438 59218
rect 9438 59166 9490 59218
rect 9490 59166 9492 59218
rect 9436 59164 9492 59166
rect 9772 59724 9828 59780
rect 10332 59388 10388 59444
rect 9772 58210 9828 58212
rect 9772 58158 9774 58210
rect 9774 58158 9826 58210
rect 9826 58158 9828 58210
rect 9772 58156 9828 58158
rect 10108 58156 10164 58212
rect 9436 56082 9492 56084
rect 9436 56030 9438 56082
rect 9438 56030 9490 56082
rect 9490 56030 9492 56082
rect 9436 56028 9492 56030
rect 9660 55970 9716 55972
rect 9660 55918 9662 55970
rect 9662 55918 9714 55970
rect 9714 55918 9716 55970
rect 9660 55916 9716 55918
rect 10108 56194 10164 56196
rect 10108 56142 10110 56194
rect 10110 56142 10162 56194
rect 10162 56142 10164 56194
rect 10108 56140 10164 56142
rect 9996 56028 10052 56084
rect 8764 53564 8820 53620
rect 8876 54684 8932 54740
rect 9324 55356 9380 55412
rect 9212 55244 9268 55300
rect 9772 55804 9828 55860
rect 9660 55298 9716 55300
rect 9660 55246 9662 55298
rect 9662 55246 9714 55298
rect 9714 55246 9716 55298
rect 9660 55244 9716 55246
rect 9772 54738 9828 54740
rect 9772 54686 9774 54738
rect 9774 54686 9826 54738
rect 9826 54686 9828 54738
rect 9772 54684 9828 54686
rect 8540 51996 8596 52052
rect 8540 51324 8596 51380
rect 7196 49868 7252 49924
rect 1708 49644 1764 49700
rect 2940 49698 2996 49700
rect 2940 49646 2942 49698
rect 2942 49646 2994 49698
rect 2994 49646 2996 49698
rect 2940 49644 2996 49646
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 1708 49084 1764 49140
rect 2044 48914 2100 48916
rect 2044 48862 2046 48914
rect 2046 48862 2098 48914
rect 2098 48862 2100 48914
rect 2044 48860 2100 48862
rect 1708 48412 1764 48468
rect 2492 48412 2548 48468
rect 8764 50204 8820 50260
rect 8204 49756 8260 49812
rect 9100 54460 9156 54516
rect 8988 51772 9044 51828
rect 6636 48914 6692 48916
rect 6636 48862 6638 48914
rect 6638 48862 6690 48914
rect 6690 48862 6692 48914
rect 6636 48860 6692 48862
rect 5964 48412 6020 48468
rect 6636 48466 6692 48468
rect 6636 48414 6638 48466
rect 6638 48414 6690 48466
rect 6690 48414 6692 48466
rect 6636 48412 6692 48414
rect 2044 48354 2100 48356
rect 2044 48302 2046 48354
rect 2046 48302 2098 48354
rect 2098 48302 2100 48354
rect 2044 48300 2100 48302
rect 1708 47740 1764 47796
rect 7084 48748 7140 48804
rect 7980 48300 8036 48356
rect 2492 47740 2548 47796
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 2044 45218 2100 45220
rect 2044 45166 2046 45218
rect 2046 45166 2098 45218
rect 2098 45166 2100 45218
rect 2044 45164 2100 45166
rect 1708 44940 1764 44996
rect 2492 44994 2548 44996
rect 2492 44942 2494 44994
rect 2494 44942 2546 44994
rect 2546 44942 2548 44994
rect 2492 44940 2548 44942
rect 5964 44828 6020 44884
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 1708 44380 1764 44436
rect 2044 44098 2100 44100
rect 2044 44046 2046 44098
rect 2046 44046 2098 44098
rect 2098 44046 2100 44098
rect 2044 44044 2100 44046
rect 1708 43708 1764 43764
rect 2492 43708 2548 43764
rect 5292 43538 5348 43540
rect 5292 43486 5294 43538
rect 5294 43486 5346 43538
rect 5346 43486 5348 43538
rect 5292 43484 5348 43486
rect 6636 45164 6692 45220
rect 6860 44882 6916 44884
rect 6860 44830 6862 44882
rect 6862 44830 6914 44882
rect 6914 44830 6916 44882
rect 6860 44828 6916 44830
rect 6972 44716 7028 44772
rect 8428 48802 8484 48804
rect 8428 48750 8430 48802
rect 8430 48750 8482 48802
rect 8482 48750 8484 48802
rect 8428 48748 8484 48750
rect 7308 46508 7364 46564
rect 8540 46562 8596 46564
rect 8540 46510 8542 46562
rect 8542 46510 8594 46562
rect 8594 46510 8596 46562
rect 8540 46508 8596 46510
rect 8092 44716 8148 44772
rect 9100 49756 9156 49812
rect 8876 47292 8932 47348
rect 8876 46956 8932 47012
rect 8764 46786 8820 46788
rect 8764 46734 8766 46786
rect 8766 46734 8818 46786
rect 8818 46734 8820 46786
rect 8764 46732 8820 46734
rect 8988 46674 9044 46676
rect 8988 46622 8990 46674
rect 8990 46622 9042 46674
rect 9042 46622 9044 46674
rect 8988 46620 9044 46622
rect 9212 45276 9268 45332
rect 8764 45164 8820 45220
rect 7644 44098 7700 44100
rect 7644 44046 7646 44098
rect 7646 44046 7698 44098
rect 7698 44046 7700 44098
rect 7644 44044 7700 44046
rect 8204 43762 8260 43764
rect 8204 43710 8206 43762
rect 8206 43710 8258 43762
rect 8258 43710 8260 43762
rect 8204 43708 8260 43710
rect 6524 43484 6580 43540
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 6524 42700 6580 42756
rect 7084 42754 7140 42756
rect 7084 42702 7086 42754
rect 7086 42702 7138 42754
rect 7138 42702 7140 42754
rect 7084 42700 7140 42702
rect 8316 42476 8372 42532
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 1820 41020 1876 41076
rect 2492 41074 2548 41076
rect 2492 41022 2494 41074
rect 2494 41022 2546 41074
rect 2546 41022 2548 41074
rect 2492 41020 2548 41022
rect 2044 40962 2100 40964
rect 2044 40910 2046 40962
rect 2046 40910 2098 40962
rect 2098 40910 2100 40962
rect 2044 40908 2100 40910
rect 1820 40348 1876 40404
rect 1708 40236 1764 40292
rect 1708 39676 1764 39732
rect 2492 40236 2548 40292
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 2044 39564 2100 39620
rect 9548 53676 9604 53732
rect 9436 51772 9492 51828
rect 9772 51884 9828 51940
rect 9996 51660 10052 51716
rect 10556 55020 10612 55076
rect 10220 51884 10276 51940
rect 9772 51378 9828 51380
rect 9772 51326 9774 51378
rect 9774 51326 9826 51378
rect 9826 51326 9828 51378
rect 9772 51324 9828 51326
rect 9660 50540 9716 50596
rect 9548 50482 9604 50484
rect 9548 50430 9550 50482
rect 9550 50430 9602 50482
rect 9602 50430 9604 50482
rect 9548 50428 9604 50430
rect 9772 50482 9828 50484
rect 9772 50430 9774 50482
rect 9774 50430 9826 50482
rect 9826 50430 9828 50482
rect 9772 50428 9828 50430
rect 10668 50428 10724 50484
rect 10332 50204 10388 50260
rect 9772 49644 9828 49700
rect 9660 46956 9716 47012
rect 9436 46786 9492 46788
rect 9436 46734 9438 46786
rect 9438 46734 9490 46786
rect 9490 46734 9492 46786
rect 9436 46732 9492 46734
rect 9660 45724 9716 45780
rect 9436 44156 9492 44212
rect 10220 49810 10276 49812
rect 10220 49758 10222 49810
rect 10222 49758 10274 49810
rect 10274 49758 10276 49810
rect 10220 49756 10276 49758
rect 10556 48412 10612 48468
rect 10220 47292 10276 47348
rect 9884 45330 9940 45332
rect 9884 45278 9886 45330
rect 9886 45278 9938 45330
rect 9938 45278 9940 45330
rect 9884 45276 9940 45278
rect 12460 61292 12516 61348
rect 11788 60396 11844 60452
rect 12236 60396 12292 60452
rect 11116 59442 11172 59444
rect 11116 59390 11118 59442
rect 11118 59390 11170 59442
rect 11170 59390 11172 59442
rect 11116 59388 11172 59390
rect 11452 58604 11508 58660
rect 14140 67842 14196 67844
rect 14140 67790 14142 67842
rect 14142 67790 14194 67842
rect 14194 67790 14196 67842
rect 14140 67788 14196 67790
rect 13916 66780 13972 66836
rect 13356 64652 13412 64708
rect 12684 62748 12740 62804
rect 13244 62412 13300 62468
rect 13916 63868 13972 63924
rect 13692 63810 13748 63812
rect 13692 63758 13694 63810
rect 13694 63758 13746 63810
rect 13746 63758 13748 63810
rect 13692 63756 13748 63758
rect 14140 64706 14196 64708
rect 14140 64654 14142 64706
rect 14142 64654 14194 64706
rect 14194 64654 14196 64706
rect 14140 64652 14196 64654
rect 15820 68460 15876 68516
rect 15484 67842 15540 67844
rect 15484 67790 15486 67842
rect 15486 67790 15538 67842
rect 15538 67790 15540 67842
rect 15484 67788 15540 67790
rect 15820 67788 15876 67844
rect 14476 67676 14532 67732
rect 16604 67676 16660 67732
rect 16716 67900 16772 67956
rect 14588 63868 14644 63924
rect 13916 62412 13972 62468
rect 13804 62076 13860 62132
rect 13804 61458 13860 61460
rect 13804 61406 13806 61458
rect 13806 61406 13858 61458
rect 13858 61406 13860 61458
rect 13804 61404 13860 61406
rect 13580 61292 13636 61348
rect 13244 60396 13300 60452
rect 13468 59890 13524 59892
rect 13468 59838 13470 59890
rect 13470 59838 13522 59890
rect 13522 59838 13524 59890
rect 13468 59836 13524 59838
rect 13356 59724 13412 59780
rect 12908 58156 12964 58212
rect 13020 57762 13076 57764
rect 13020 57710 13022 57762
rect 13022 57710 13074 57762
rect 13074 57710 13076 57762
rect 13020 57708 13076 57710
rect 13692 59778 13748 59780
rect 13692 59726 13694 59778
rect 13694 59726 13746 59778
rect 13746 59726 13748 59778
rect 13692 59724 13748 59726
rect 14364 63308 14420 63364
rect 15708 62972 15764 63028
rect 14924 62748 14980 62804
rect 14700 62578 14756 62580
rect 14700 62526 14702 62578
rect 14702 62526 14754 62578
rect 14754 62526 14756 62578
rect 14700 62524 14756 62526
rect 13692 58658 13748 58660
rect 13692 58606 13694 58658
rect 13694 58606 13746 58658
rect 13746 58606 13748 58658
rect 13692 58604 13748 58606
rect 13468 58210 13524 58212
rect 13468 58158 13470 58210
rect 13470 58158 13522 58210
rect 13522 58158 13524 58210
rect 13468 58156 13524 58158
rect 11564 55410 11620 55412
rect 11564 55358 11566 55410
rect 11566 55358 11618 55410
rect 11618 55358 11620 55410
rect 11564 55356 11620 55358
rect 11004 55074 11060 55076
rect 11004 55022 11006 55074
rect 11006 55022 11058 55074
rect 11058 55022 11060 55074
rect 11004 55020 11060 55022
rect 11900 55020 11956 55076
rect 12012 55468 12068 55524
rect 12908 56812 12964 56868
rect 12236 55356 12292 55412
rect 12684 56588 12740 56644
rect 11452 52162 11508 52164
rect 11452 52110 11454 52162
rect 11454 52110 11506 52162
rect 11506 52110 11508 52162
rect 11452 52108 11508 52110
rect 11788 52108 11844 52164
rect 11676 51938 11732 51940
rect 11676 51886 11678 51938
rect 11678 51886 11730 51938
rect 11730 51886 11732 51938
rect 11676 51884 11732 51886
rect 11452 51436 11508 51492
rect 11452 50428 11508 50484
rect 11228 50316 11284 50372
rect 10220 45218 10276 45220
rect 10220 45166 10222 45218
rect 10222 45166 10274 45218
rect 10274 45166 10276 45218
rect 10220 45164 10276 45166
rect 10780 46844 10836 46900
rect 10780 46620 10836 46676
rect 10780 45724 10836 45780
rect 10892 45106 10948 45108
rect 10892 45054 10894 45106
rect 10894 45054 10946 45106
rect 10946 45054 10948 45106
rect 10892 45052 10948 45054
rect 9212 41244 9268 41300
rect 9660 40908 9716 40964
rect 9884 42866 9940 42868
rect 9884 42814 9886 42866
rect 9886 42814 9938 42866
rect 9938 42814 9940 42866
rect 9884 42812 9940 42814
rect 9772 40626 9828 40628
rect 9772 40574 9774 40626
rect 9774 40574 9826 40626
rect 9826 40574 9828 40626
rect 9772 40572 9828 40574
rect 10108 42700 10164 42756
rect 10556 42812 10612 42868
rect 10556 42530 10612 42532
rect 10556 42478 10558 42530
rect 10558 42478 10610 42530
rect 10610 42478 10612 42530
rect 10556 42476 10612 42478
rect 12124 52162 12180 52164
rect 12124 52110 12126 52162
rect 12126 52110 12178 52162
rect 12178 52110 12180 52162
rect 12124 52108 12180 52110
rect 12460 54796 12516 54852
rect 13468 56642 13524 56644
rect 13468 56590 13470 56642
rect 13470 56590 13522 56642
rect 13522 56590 13524 56642
rect 13468 56588 13524 56590
rect 14364 62354 14420 62356
rect 14364 62302 14366 62354
rect 14366 62302 14418 62354
rect 14418 62302 14420 62354
rect 14364 62300 14420 62302
rect 16044 62748 16100 62804
rect 15596 62354 15652 62356
rect 15596 62302 15598 62354
rect 15598 62302 15650 62354
rect 15650 62302 15652 62354
rect 15596 62300 15652 62302
rect 14812 61292 14868 61348
rect 14476 59890 14532 59892
rect 14476 59838 14478 59890
rect 14478 59838 14530 59890
rect 14530 59838 14532 59890
rect 14476 59836 14532 59838
rect 15036 59836 15092 59892
rect 14252 58434 14308 58436
rect 14252 58382 14254 58434
rect 14254 58382 14306 58434
rect 14306 58382 14308 58434
rect 14252 58380 14308 58382
rect 17612 69356 17668 69412
rect 17724 68514 17780 68516
rect 17724 68462 17726 68514
rect 17726 68462 17778 68514
rect 17778 68462 17780 68514
rect 17724 68460 17780 68462
rect 17612 68348 17668 68404
rect 17388 67900 17444 67956
rect 17836 67900 17892 67956
rect 17724 67842 17780 67844
rect 17724 67790 17726 67842
rect 17726 67790 17778 67842
rect 17778 67790 17780 67842
rect 17724 67788 17780 67790
rect 17948 67564 18004 67620
rect 16716 66834 16772 66836
rect 16716 66782 16718 66834
rect 16718 66782 16770 66834
rect 16770 66782 16772 66834
rect 16716 66780 16772 66782
rect 18172 69356 18228 69412
rect 18172 67730 18228 67732
rect 18172 67678 18174 67730
rect 18174 67678 18226 67730
rect 18226 67678 18228 67730
rect 18172 67676 18228 67678
rect 19516 69580 19572 69636
rect 18956 68626 19012 68628
rect 18956 68574 18958 68626
rect 18958 68574 19010 68626
rect 19010 68574 19012 68626
rect 18956 68572 19012 68574
rect 18508 67564 18564 67620
rect 18396 66892 18452 66948
rect 17836 63196 17892 63252
rect 16492 62972 16548 63028
rect 17276 63026 17332 63028
rect 17276 62974 17278 63026
rect 17278 62974 17330 63026
rect 17330 62974 17332 63026
rect 17276 62972 17332 62974
rect 17388 62860 17444 62916
rect 16828 62578 16884 62580
rect 16828 62526 16830 62578
rect 16830 62526 16882 62578
rect 16882 62526 16884 62578
rect 16828 62524 16884 62526
rect 17836 62636 17892 62692
rect 18284 63756 18340 63812
rect 19852 69580 19908 69636
rect 20076 69468 20132 69524
rect 20636 69634 20692 69636
rect 20636 69582 20638 69634
rect 20638 69582 20690 69634
rect 20690 69582 20692 69634
rect 20636 69580 20692 69582
rect 20412 69522 20468 69524
rect 20412 69470 20414 69522
rect 20414 69470 20466 69522
rect 20466 69470 20468 69522
rect 20412 69468 20468 69470
rect 19836 69018 19892 69020
rect 19836 68966 19838 69018
rect 19838 68966 19890 69018
rect 19890 68966 19892 69018
rect 19836 68964 19892 68966
rect 19940 69018 19996 69020
rect 19940 68966 19942 69018
rect 19942 68966 19994 69018
rect 19994 68966 19996 69018
rect 19940 68964 19996 68966
rect 20044 69018 20100 69020
rect 20044 68966 20046 69018
rect 20046 68966 20098 69018
rect 20098 68966 20100 69018
rect 20044 68964 20100 68966
rect 19628 68796 19684 68852
rect 20412 68796 20468 68852
rect 19628 68460 19684 68516
rect 20076 68348 20132 68404
rect 19836 67450 19892 67452
rect 19836 67398 19838 67450
rect 19838 67398 19890 67450
rect 19890 67398 19892 67450
rect 19836 67396 19892 67398
rect 19940 67450 19996 67452
rect 19940 67398 19942 67450
rect 19942 67398 19994 67450
rect 19994 67398 19996 67450
rect 19940 67396 19996 67398
rect 20044 67450 20100 67452
rect 20044 67398 20046 67450
rect 20046 67398 20098 67450
rect 20098 67398 20100 67450
rect 20044 67396 20100 67398
rect 20524 68460 20580 68516
rect 21084 68514 21140 68516
rect 21084 68462 21086 68514
rect 21086 68462 21138 68514
rect 21138 68462 21140 68514
rect 21084 68460 21140 68462
rect 24444 69916 24500 69972
rect 22316 69522 22372 69524
rect 22316 69470 22318 69522
rect 22318 69470 22370 69522
rect 22370 69470 22372 69522
rect 22316 69468 22372 69470
rect 23548 69468 23604 69524
rect 25228 69970 25284 69972
rect 25228 69918 25230 69970
rect 25230 69918 25282 69970
rect 25282 69918 25284 69970
rect 25228 69916 25284 69918
rect 25564 70082 25620 70084
rect 25564 70030 25566 70082
rect 25566 70030 25618 70082
rect 25618 70030 25620 70082
rect 25564 70028 25620 70030
rect 26124 70082 26180 70084
rect 26124 70030 26126 70082
rect 26126 70030 26178 70082
rect 26178 70030 26180 70082
rect 26124 70028 26180 70030
rect 27692 70028 27748 70084
rect 24668 68738 24724 68740
rect 24668 68686 24670 68738
rect 24670 68686 24722 68738
rect 24722 68686 24724 68738
rect 24668 68684 24724 68686
rect 24332 68460 24388 68516
rect 23996 68124 24052 68180
rect 24556 67954 24612 67956
rect 24556 67902 24558 67954
rect 24558 67902 24610 67954
rect 24610 67902 24612 67954
rect 24556 67900 24612 67902
rect 24668 68460 24724 68516
rect 19516 66780 19572 66836
rect 19836 65882 19892 65884
rect 19836 65830 19838 65882
rect 19838 65830 19890 65882
rect 19890 65830 19892 65882
rect 19836 65828 19892 65830
rect 19940 65882 19996 65884
rect 19940 65830 19942 65882
rect 19942 65830 19994 65882
rect 19994 65830 19996 65882
rect 19940 65828 19996 65830
rect 20044 65882 20100 65884
rect 20044 65830 20046 65882
rect 20046 65830 20098 65882
rect 20098 65830 20100 65882
rect 20044 65828 20100 65830
rect 19836 64314 19892 64316
rect 19836 64262 19838 64314
rect 19838 64262 19890 64314
rect 19890 64262 19892 64314
rect 19836 64260 19892 64262
rect 19940 64314 19996 64316
rect 19940 64262 19942 64314
rect 19942 64262 19994 64314
rect 19994 64262 19996 64314
rect 19940 64260 19996 64262
rect 20044 64314 20100 64316
rect 20044 64262 20046 64314
rect 20046 64262 20098 64314
rect 20098 64262 20100 64314
rect 20044 64260 20100 64262
rect 18060 63362 18116 63364
rect 18060 63310 18062 63362
rect 18062 63310 18114 63362
rect 18114 63310 18116 63362
rect 18060 63308 18116 63310
rect 18956 63308 19012 63364
rect 19404 63138 19460 63140
rect 19404 63086 19406 63138
rect 19406 63086 19458 63138
rect 19458 63086 19460 63138
rect 19404 63084 19460 63086
rect 18396 62972 18452 63028
rect 17612 62188 17668 62244
rect 17724 62300 17780 62356
rect 17612 61404 17668 61460
rect 16828 59218 16884 59220
rect 16828 59166 16830 59218
rect 16830 59166 16882 59218
rect 16882 59166 16884 59218
rect 16828 59164 16884 59166
rect 14028 56866 14084 56868
rect 14028 56814 14030 56866
rect 14030 56814 14082 56866
rect 14082 56814 14084 56866
rect 14028 56812 14084 56814
rect 15036 57372 15092 57428
rect 14252 56754 14308 56756
rect 14252 56702 14254 56754
rect 14254 56702 14306 56754
rect 14306 56702 14308 56754
rect 14252 56700 14308 56702
rect 13692 54796 13748 54852
rect 16716 57596 16772 57652
rect 16604 56924 16660 56980
rect 15484 56642 15540 56644
rect 15484 56590 15486 56642
rect 15486 56590 15538 56642
rect 15538 56590 15540 56642
rect 15484 56588 15540 56590
rect 14924 54572 14980 54628
rect 15484 54572 15540 54628
rect 17388 59890 17444 59892
rect 17388 59838 17390 59890
rect 17390 59838 17442 59890
rect 17442 59838 17444 59890
rect 17388 59836 17444 59838
rect 17948 62524 18004 62580
rect 18172 61516 18228 61572
rect 18844 62860 18900 62916
rect 18732 62412 18788 62468
rect 19516 62466 19572 62468
rect 19516 62414 19518 62466
rect 19518 62414 19570 62466
rect 19570 62414 19572 62466
rect 19516 62412 19572 62414
rect 18956 62354 19012 62356
rect 18956 62302 18958 62354
rect 18958 62302 19010 62354
rect 19010 62302 19012 62354
rect 18956 62300 19012 62302
rect 18956 61852 19012 61908
rect 19964 63308 20020 63364
rect 20188 63196 20244 63252
rect 19836 62746 19892 62748
rect 19836 62694 19838 62746
rect 19838 62694 19890 62746
rect 19890 62694 19892 62746
rect 19836 62692 19892 62694
rect 19940 62746 19996 62748
rect 19940 62694 19942 62746
rect 19942 62694 19994 62746
rect 19994 62694 19996 62746
rect 19940 62692 19996 62694
rect 20044 62746 20100 62748
rect 20044 62694 20046 62746
rect 20046 62694 20098 62746
rect 20098 62694 20100 62746
rect 20044 62692 20100 62694
rect 19628 62300 19684 62356
rect 19628 62130 19684 62132
rect 19628 62078 19630 62130
rect 19630 62078 19682 62130
rect 19682 62078 19684 62130
rect 19628 62076 19684 62078
rect 19292 61852 19348 61908
rect 19964 61852 20020 61908
rect 19740 61794 19796 61796
rect 19740 61742 19742 61794
rect 19742 61742 19794 61794
rect 19794 61742 19796 61794
rect 19740 61740 19796 61742
rect 18732 61458 18788 61460
rect 18732 61406 18734 61458
rect 18734 61406 18786 61458
rect 18786 61406 18788 61458
rect 18732 61404 18788 61406
rect 18172 59948 18228 60004
rect 18732 60786 18788 60788
rect 18732 60734 18734 60786
rect 18734 60734 18786 60786
rect 18786 60734 18788 60786
rect 18732 60732 18788 60734
rect 17612 59218 17668 59220
rect 17612 59166 17614 59218
rect 17614 59166 17666 59218
rect 17666 59166 17668 59218
rect 17612 59164 17668 59166
rect 17500 58156 17556 58212
rect 19404 61292 19460 61348
rect 20188 61852 20244 61908
rect 20188 61570 20244 61572
rect 20188 61518 20190 61570
rect 20190 61518 20242 61570
rect 20242 61518 20244 61570
rect 20188 61516 20244 61518
rect 19628 61180 19684 61236
rect 19404 60732 19460 60788
rect 19292 60002 19348 60004
rect 19292 59950 19294 60002
rect 19294 59950 19346 60002
rect 19346 59950 19348 60002
rect 19292 59948 19348 59950
rect 19516 60844 19572 60900
rect 19836 61178 19892 61180
rect 19836 61126 19838 61178
rect 19838 61126 19890 61178
rect 19890 61126 19892 61178
rect 19836 61124 19892 61126
rect 19940 61178 19996 61180
rect 19940 61126 19942 61178
rect 19942 61126 19994 61178
rect 19994 61126 19996 61178
rect 19940 61124 19996 61126
rect 20044 61178 20100 61180
rect 20044 61126 20046 61178
rect 20046 61126 20098 61178
rect 20098 61126 20100 61178
rect 20044 61124 20100 61126
rect 20076 60674 20132 60676
rect 20076 60622 20078 60674
rect 20078 60622 20130 60674
rect 20130 60622 20132 60674
rect 20076 60620 20132 60622
rect 19964 60508 20020 60564
rect 20412 62076 20468 62132
rect 20748 61458 20804 61460
rect 20748 61406 20750 61458
rect 20750 61406 20802 61458
rect 20802 61406 20804 61458
rect 20748 61404 20804 61406
rect 25116 68124 25172 68180
rect 25228 68796 25284 68852
rect 26124 68796 26180 68852
rect 25788 68738 25844 68740
rect 25788 68686 25790 68738
rect 25790 68686 25842 68738
rect 25842 68686 25844 68738
rect 25788 68684 25844 68686
rect 25452 68460 25508 68516
rect 23884 67730 23940 67732
rect 23884 67678 23886 67730
rect 23886 67678 23938 67730
rect 23938 67678 23940 67730
rect 23884 67676 23940 67678
rect 24668 67676 24724 67732
rect 25452 67900 25508 67956
rect 23548 67004 23604 67060
rect 25788 68124 25844 68180
rect 25228 67058 25284 67060
rect 25228 67006 25230 67058
rect 25230 67006 25282 67058
rect 25282 67006 25284 67058
rect 25228 67004 25284 67006
rect 25676 67004 25732 67060
rect 22988 65436 23044 65492
rect 23884 65490 23940 65492
rect 23884 65438 23886 65490
rect 23886 65438 23938 65490
rect 23938 65438 23940 65490
rect 23884 65436 23940 65438
rect 24668 65490 24724 65492
rect 24668 65438 24670 65490
rect 24670 65438 24722 65490
rect 24722 65438 24724 65490
rect 24668 65436 24724 65438
rect 25340 65436 25396 65492
rect 24444 64428 24500 64484
rect 25340 64428 25396 64484
rect 24332 63922 24388 63924
rect 24332 63870 24334 63922
rect 24334 63870 24386 63922
rect 24386 63870 24388 63922
rect 24332 63868 24388 63870
rect 21420 63810 21476 63812
rect 21420 63758 21422 63810
rect 21422 63758 21474 63810
rect 21474 63758 21476 63810
rect 21420 63756 21476 63758
rect 21420 63084 21476 63140
rect 21532 63196 21588 63252
rect 22764 63138 22820 63140
rect 22764 63086 22766 63138
rect 22766 63086 22818 63138
rect 22818 63086 22820 63138
rect 22764 63084 22820 63086
rect 22092 62412 22148 62468
rect 24332 63084 24388 63140
rect 23324 62412 23380 62468
rect 23884 62860 23940 62916
rect 25788 66892 25844 66948
rect 25452 63980 25508 64036
rect 24892 63138 24948 63140
rect 24892 63086 24894 63138
rect 24894 63086 24946 63138
rect 24946 63086 24948 63138
rect 24892 63084 24948 63086
rect 24668 62860 24724 62916
rect 24556 62466 24612 62468
rect 24556 62414 24558 62466
rect 24558 62414 24610 62466
rect 24610 62414 24612 62466
rect 24556 62412 24612 62414
rect 24220 62354 24276 62356
rect 24220 62302 24222 62354
rect 24222 62302 24274 62354
rect 24274 62302 24276 62354
rect 24220 62300 24276 62302
rect 23324 61458 23380 61460
rect 23324 61406 23326 61458
rect 23326 61406 23378 61458
rect 23378 61406 23380 61458
rect 23324 61404 23380 61406
rect 23212 61346 23268 61348
rect 23212 61294 23214 61346
rect 23214 61294 23266 61346
rect 23266 61294 23268 61346
rect 23212 61292 23268 61294
rect 24444 61346 24500 61348
rect 24444 61294 24446 61346
rect 24446 61294 24498 61346
rect 24498 61294 24500 61346
rect 24444 61292 24500 61294
rect 18508 59218 18564 59220
rect 18508 59166 18510 59218
rect 18510 59166 18562 59218
rect 18562 59166 18564 59218
rect 18508 59164 18564 59166
rect 17836 58434 17892 58436
rect 17836 58382 17838 58434
rect 17838 58382 17890 58434
rect 17890 58382 17892 58434
rect 17836 58380 17892 58382
rect 17276 56924 17332 56980
rect 17164 56642 17220 56644
rect 17164 56590 17166 56642
rect 17166 56590 17218 56642
rect 17218 56590 17220 56642
rect 17164 56588 17220 56590
rect 17724 57650 17780 57652
rect 17724 57598 17726 57650
rect 17726 57598 17778 57650
rect 17778 57598 17780 57650
rect 17724 57596 17780 57598
rect 17612 57372 17668 57428
rect 16604 55804 16660 55860
rect 15260 53228 15316 53284
rect 15148 53004 15204 53060
rect 17164 55186 17220 55188
rect 17164 55134 17166 55186
rect 17166 55134 17218 55186
rect 17218 55134 17220 55186
rect 17164 55132 17220 55134
rect 12236 51884 12292 51940
rect 11676 50540 11732 50596
rect 12124 50594 12180 50596
rect 12124 50542 12126 50594
rect 12126 50542 12178 50594
rect 12178 50542 12180 50594
rect 12124 50540 12180 50542
rect 12908 52050 12964 52052
rect 12908 51998 12910 52050
rect 12910 51998 12962 52050
rect 12962 51998 12964 52050
rect 12908 51996 12964 51998
rect 15036 52946 15092 52948
rect 15036 52894 15038 52946
rect 15038 52894 15090 52946
rect 15090 52894 15092 52946
rect 15036 52892 15092 52894
rect 15596 52668 15652 52724
rect 15596 51996 15652 52052
rect 14812 51436 14868 51492
rect 16044 53116 16100 53172
rect 16380 53618 16436 53620
rect 16380 53566 16382 53618
rect 16382 53566 16434 53618
rect 16434 53566 16436 53618
rect 16380 53564 16436 53566
rect 16940 53564 16996 53620
rect 16380 52892 16436 52948
rect 16492 53452 16548 53508
rect 18956 58210 19012 58212
rect 18956 58158 18958 58210
rect 18958 58158 19010 58210
rect 19010 58158 19012 58210
rect 18956 58156 19012 58158
rect 18620 57372 18676 57428
rect 18396 57036 18452 57092
rect 18060 56978 18116 56980
rect 18060 56926 18062 56978
rect 18062 56926 18114 56978
rect 18114 56926 18116 56978
rect 18060 56924 18116 56926
rect 18732 56140 18788 56196
rect 17500 56082 17556 56084
rect 17500 56030 17502 56082
rect 17502 56030 17554 56082
rect 17554 56030 17556 56082
rect 17500 56028 17556 56030
rect 17388 55244 17444 55300
rect 17836 55804 17892 55860
rect 17724 55356 17780 55412
rect 18396 55804 18452 55860
rect 17724 54572 17780 54628
rect 18172 53676 18228 53732
rect 18284 54460 18340 54516
rect 16268 52834 16324 52836
rect 16268 52782 16270 52834
rect 16270 52782 16322 52834
rect 16322 52782 16324 52834
rect 16268 52780 16324 52782
rect 18172 53452 18228 53508
rect 16604 53004 16660 53060
rect 17388 52946 17444 52948
rect 17388 52894 17390 52946
rect 17390 52894 17442 52946
rect 17442 52894 17444 52946
rect 17388 52892 17444 52894
rect 16716 52108 16772 52164
rect 16492 51884 16548 51940
rect 16716 51884 16772 51940
rect 14588 51266 14644 51268
rect 14588 51214 14590 51266
rect 14590 51214 14642 51266
rect 14642 51214 14644 51266
rect 14588 51212 14644 51214
rect 15708 51212 15764 51268
rect 12684 50428 12740 50484
rect 12908 50482 12964 50484
rect 12908 50430 12910 50482
rect 12910 50430 12962 50482
rect 12962 50430 12964 50482
rect 12908 50428 12964 50430
rect 15148 50482 15204 50484
rect 15148 50430 15150 50482
rect 15150 50430 15202 50482
rect 15202 50430 15204 50482
rect 15148 50428 15204 50430
rect 14812 50204 14868 50260
rect 15708 50428 15764 50484
rect 15260 50204 15316 50260
rect 14812 49308 14868 49364
rect 15708 49980 15764 50036
rect 18172 52780 18228 52836
rect 17948 51884 18004 51940
rect 16604 51490 16660 51492
rect 16604 51438 16606 51490
rect 16606 51438 16658 51490
rect 16658 51438 16660 51490
rect 16604 51436 16660 51438
rect 17836 51772 17892 51828
rect 16268 50540 16324 50596
rect 16380 50482 16436 50484
rect 16380 50430 16382 50482
rect 16382 50430 16434 50482
rect 16434 50430 16436 50482
rect 16380 50428 16436 50430
rect 11900 48242 11956 48244
rect 11900 48190 11902 48242
rect 11902 48190 11954 48242
rect 11954 48190 11956 48242
rect 11900 48188 11956 48190
rect 11340 47292 11396 47348
rect 11340 46898 11396 46900
rect 11340 46846 11342 46898
rect 11342 46846 11394 46898
rect 11394 46846 11396 46898
rect 11340 46844 11396 46846
rect 14924 46002 14980 46004
rect 14924 45950 14926 46002
rect 14926 45950 14978 46002
rect 14978 45950 14980 46002
rect 14924 45948 14980 45950
rect 14252 45836 14308 45892
rect 15036 45836 15092 45892
rect 12908 45612 12964 45668
rect 13916 45666 13972 45668
rect 13916 45614 13918 45666
rect 13918 45614 13970 45666
rect 13970 45614 13972 45666
rect 13916 45612 13972 45614
rect 12572 45052 12628 45108
rect 12908 44268 12964 44324
rect 13580 44322 13636 44324
rect 13580 44270 13582 44322
rect 13582 44270 13634 44322
rect 13634 44270 13636 44322
rect 13580 44268 13636 44270
rect 14588 45612 14644 45668
rect 14812 45330 14868 45332
rect 14812 45278 14814 45330
rect 14814 45278 14866 45330
rect 14866 45278 14868 45330
rect 14812 45276 14868 45278
rect 14476 45106 14532 45108
rect 14476 45054 14478 45106
rect 14478 45054 14530 45106
rect 14530 45054 14532 45106
rect 14476 45052 14532 45054
rect 14028 44268 14084 44324
rect 13916 44156 13972 44212
rect 14028 43708 14084 43764
rect 15484 48188 15540 48244
rect 16268 48188 16324 48244
rect 15484 47292 15540 47348
rect 16604 47964 16660 48020
rect 15372 45890 15428 45892
rect 15372 45838 15374 45890
rect 15374 45838 15426 45890
rect 15426 45838 15428 45890
rect 15372 45836 15428 45838
rect 15484 45164 15540 45220
rect 15372 44044 15428 44100
rect 10444 41244 10500 41300
rect 11228 41186 11284 41188
rect 11228 41134 11230 41186
rect 11230 41134 11282 41186
rect 11282 41134 11284 41186
rect 11228 41132 11284 41134
rect 10108 41020 10164 41076
rect 9772 40178 9828 40180
rect 9772 40126 9774 40178
rect 9774 40126 9826 40178
rect 9826 40126 9828 40178
rect 9772 40124 9828 40126
rect 6972 39452 7028 39508
rect 2044 39394 2100 39396
rect 2044 39342 2046 39394
rect 2046 39342 2098 39394
rect 2098 39342 2100 39394
rect 2044 39340 2100 39342
rect 1708 39004 1764 39060
rect 2492 39004 2548 39060
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 8204 39506 8260 39508
rect 8204 39454 8206 39506
rect 8206 39454 8258 39506
rect 8258 39454 8260 39506
rect 8204 39452 8260 39454
rect 8092 39340 8148 39396
rect 7532 39004 7588 39060
rect 7644 38946 7700 38948
rect 7644 38894 7646 38946
rect 7646 38894 7698 38946
rect 7698 38894 7700 38946
rect 7644 38892 7700 38894
rect 9548 39564 9604 39620
rect 8204 39116 8260 39172
rect 8428 38834 8484 38836
rect 8428 38782 8430 38834
rect 8430 38782 8482 38834
rect 8482 38782 8484 38834
rect 8428 38780 8484 38782
rect 9436 39004 9492 39060
rect 9660 39116 9716 39172
rect 10332 40626 10388 40628
rect 10332 40574 10334 40626
rect 10334 40574 10386 40626
rect 10386 40574 10388 40626
rect 10332 40572 10388 40574
rect 9772 39004 9828 39060
rect 11228 40124 11284 40180
rect 10332 39116 10388 39172
rect 10892 39004 10948 39060
rect 9884 38946 9940 38948
rect 9884 38894 9886 38946
rect 9886 38894 9938 38946
rect 9938 38894 9940 38946
rect 9884 38892 9940 38894
rect 8764 38780 8820 38836
rect 7868 37436 7924 37492
rect 8764 37436 8820 37492
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 8092 36204 8148 36260
rect 11900 41186 11956 41188
rect 11900 41134 11902 41186
rect 11902 41134 11954 41186
rect 11954 41134 11956 41186
rect 11900 41132 11956 41134
rect 11564 40460 11620 40516
rect 12908 40460 12964 40516
rect 13468 40460 13524 40516
rect 12572 39004 12628 39060
rect 12684 38946 12740 38948
rect 12684 38894 12686 38946
rect 12686 38894 12738 38946
rect 12738 38894 12740 38946
rect 12684 38892 12740 38894
rect 13692 39452 13748 39508
rect 14140 43372 14196 43428
rect 15708 44322 15764 44324
rect 15708 44270 15710 44322
rect 15710 44270 15762 44322
rect 15762 44270 15764 44322
rect 15708 44268 15764 44270
rect 15708 43708 15764 43764
rect 16156 44210 16212 44212
rect 16156 44158 16158 44210
rect 16158 44158 16210 44210
rect 16210 44158 16212 44210
rect 16156 44156 16212 44158
rect 16156 43538 16212 43540
rect 16156 43486 16158 43538
rect 16158 43486 16210 43538
rect 16210 43486 16212 43538
rect 16156 43484 16212 43486
rect 16940 46002 16996 46004
rect 16940 45950 16942 46002
rect 16942 45950 16994 46002
rect 16994 45950 16996 46002
rect 16940 45948 16996 45950
rect 16604 45106 16660 45108
rect 16604 45054 16606 45106
rect 16606 45054 16658 45106
rect 16658 45054 16660 45106
rect 16604 45052 16660 45054
rect 15596 43372 15652 43428
rect 15932 43426 15988 43428
rect 15932 43374 15934 43426
rect 15934 43374 15986 43426
rect 15986 43374 15988 43426
rect 15932 43372 15988 43374
rect 14700 42642 14756 42644
rect 14700 42590 14702 42642
rect 14702 42590 14754 42642
rect 14754 42590 14756 42642
rect 14700 42588 14756 42590
rect 14252 42140 14308 42196
rect 14140 41074 14196 41076
rect 14140 41022 14142 41074
rect 14142 41022 14194 41074
rect 14194 41022 14196 41074
rect 14140 41020 14196 41022
rect 16380 42588 16436 42644
rect 15708 40124 15764 40180
rect 14028 39228 14084 39284
rect 13244 39004 13300 39060
rect 14028 38946 14084 38948
rect 14028 38894 14030 38946
rect 14030 38894 14082 38946
rect 14082 38894 14084 38946
rect 14028 38892 14084 38894
rect 14700 38892 14756 38948
rect 13132 37996 13188 38052
rect 10332 36204 10388 36260
rect 11340 36258 11396 36260
rect 11340 36206 11342 36258
rect 11342 36206 11394 36258
rect 11394 36206 11396 36258
rect 11340 36204 11396 36206
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 12236 35084 12292 35140
rect 13468 35138 13524 35140
rect 13468 35086 13470 35138
rect 13470 35086 13522 35138
rect 13522 35086 13524 35138
rect 13468 35084 13524 35086
rect 14028 38050 14084 38052
rect 14028 37998 14030 38050
rect 14030 37998 14082 38050
rect 14082 37998 14084 38050
rect 14028 37996 14084 37998
rect 16604 42140 16660 42196
rect 17052 44492 17108 44548
rect 16716 41804 16772 41860
rect 16604 41692 16660 41748
rect 17724 50540 17780 50596
rect 18844 54626 18900 54628
rect 18844 54574 18846 54626
rect 18846 54574 18898 54626
rect 18898 54574 18900 54626
rect 18844 54572 18900 54574
rect 18956 54460 19012 54516
rect 19068 55244 19124 55300
rect 18396 53452 18452 53508
rect 19292 55132 19348 55188
rect 19836 59610 19892 59612
rect 19836 59558 19838 59610
rect 19838 59558 19890 59610
rect 19890 59558 19892 59610
rect 19836 59556 19892 59558
rect 19940 59610 19996 59612
rect 19940 59558 19942 59610
rect 19942 59558 19994 59610
rect 19994 59558 19996 59610
rect 19940 59556 19996 59558
rect 20044 59610 20100 59612
rect 20044 59558 20046 59610
rect 20046 59558 20098 59610
rect 20098 59558 20100 59610
rect 20044 59556 20100 59558
rect 21084 60956 21140 61012
rect 22204 61010 22260 61012
rect 22204 60958 22206 61010
rect 22206 60958 22258 61010
rect 22258 60958 22260 61010
rect 22204 60956 22260 60958
rect 21308 60562 21364 60564
rect 21308 60510 21310 60562
rect 21310 60510 21362 60562
rect 21362 60510 21364 60562
rect 21308 60508 21364 60510
rect 19836 58042 19892 58044
rect 19836 57990 19838 58042
rect 19838 57990 19890 58042
rect 19890 57990 19892 58042
rect 19836 57988 19892 57990
rect 19940 58042 19996 58044
rect 19940 57990 19942 58042
rect 19942 57990 19994 58042
rect 19994 57990 19996 58042
rect 19940 57988 19996 57990
rect 20044 58042 20100 58044
rect 20044 57990 20046 58042
rect 20046 57990 20098 58042
rect 20098 57990 20100 58042
rect 20044 57988 20100 57990
rect 19836 56474 19892 56476
rect 19836 56422 19838 56474
rect 19838 56422 19890 56474
rect 19890 56422 19892 56474
rect 19836 56420 19892 56422
rect 19940 56474 19996 56476
rect 19940 56422 19942 56474
rect 19942 56422 19994 56474
rect 19994 56422 19996 56474
rect 19940 56420 19996 56422
rect 20044 56474 20100 56476
rect 20044 56422 20046 56474
rect 20046 56422 20098 56474
rect 20098 56422 20100 56474
rect 20044 56420 20100 56422
rect 19836 54906 19892 54908
rect 19836 54854 19838 54906
rect 19838 54854 19890 54906
rect 19890 54854 19892 54906
rect 19836 54852 19892 54854
rect 19940 54906 19996 54908
rect 19940 54854 19942 54906
rect 19942 54854 19994 54906
rect 19994 54854 19996 54906
rect 19940 54852 19996 54854
rect 20044 54906 20100 54908
rect 20044 54854 20046 54906
rect 20046 54854 20098 54906
rect 20098 54854 20100 54906
rect 20044 54852 20100 54854
rect 19180 53730 19236 53732
rect 19180 53678 19182 53730
rect 19182 53678 19234 53730
rect 19234 53678 19236 53730
rect 19180 53676 19236 53678
rect 19292 53564 19348 53620
rect 18956 53228 19012 53284
rect 18732 53116 18788 53172
rect 18620 52050 18676 52052
rect 18620 51998 18622 52050
rect 18622 51998 18674 52050
rect 18674 51998 18676 52050
rect 18620 51996 18676 51998
rect 18508 51884 18564 51940
rect 18508 50428 18564 50484
rect 17500 48188 17556 48244
rect 17836 49980 17892 50036
rect 18396 49980 18452 50036
rect 18172 49308 18228 49364
rect 18060 48972 18116 49028
rect 18396 48466 18452 48468
rect 18396 48414 18398 48466
rect 18398 48414 18450 48466
rect 18450 48414 18452 48466
rect 18396 48412 18452 48414
rect 19516 53506 19572 53508
rect 19516 53454 19518 53506
rect 19518 53454 19570 53506
rect 19570 53454 19572 53506
rect 19516 53452 19572 53454
rect 20076 54514 20132 54516
rect 20076 54462 20078 54514
rect 20078 54462 20130 54514
rect 20130 54462 20132 54514
rect 20076 54460 20132 54462
rect 19740 53676 19796 53732
rect 19836 53338 19892 53340
rect 19836 53286 19838 53338
rect 19838 53286 19890 53338
rect 19890 53286 19892 53338
rect 19836 53284 19892 53286
rect 19940 53338 19996 53340
rect 19940 53286 19942 53338
rect 19942 53286 19994 53338
rect 19994 53286 19996 53338
rect 19940 53284 19996 53286
rect 20044 53338 20100 53340
rect 20044 53286 20046 53338
rect 20046 53286 20098 53338
rect 20098 53286 20100 53338
rect 20044 53284 20100 53286
rect 20748 53452 20804 53508
rect 20972 52892 21028 52948
rect 20076 52668 20132 52724
rect 20748 52108 20804 52164
rect 19836 51770 19892 51772
rect 19836 51718 19838 51770
rect 19838 51718 19890 51770
rect 19890 51718 19892 51770
rect 19836 51716 19892 51718
rect 19940 51770 19996 51772
rect 19940 51718 19942 51770
rect 19942 51718 19994 51770
rect 19994 51718 19996 51770
rect 19940 51716 19996 51718
rect 20044 51770 20100 51772
rect 20044 51718 20046 51770
rect 20046 51718 20098 51770
rect 20098 51718 20100 51770
rect 20044 51716 20100 51718
rect 20748 51772 20804 51828
rect 19740 50764 19796 50820
rect 21084 51436 21140 51492
rect 21084 50764 21140 50820
rect 18956 50428 19012 50484
rect 20636 50482 20692 50484
rect 20636 50430 20638 50482
rect 20638 50430 20690 50482
rect 20690 50430 20692 50482
rect 20636 50428 20692 50430
rect 19836 50202 19892 50204
rect 19836 50150 19838 50202
rect 19838 50150 19890 50202
rect 19890 50150 19892 50202
rect 19836 50148 19892 50150
rect 19940 50202 19996 50204
rect 19940 50150 19942 50202
rect 19942 50150 19994 50202
rect 19994 50150 19996 50202
rect 19940 50148 19996 50150
rect 20044 50202 20100 50204
rect 20044 50150 20046 50202
rect 20046 50150 20098 50202
rect 20098 50150 20100 50202
rect 20044 50148 20100 50150
rect 19068 48412 19124 48468
rect 18508 48130 18564 48132
rect 18508 48078 18510 48130
rect 18510 48078 18562 48130
rect 18562 48078 18564 48130
rect 18508 48076 18564 48078
rect 18732 48242 18788 48244
rect 18732 48190 18734 48242
rect 18734 48190 18786 48242
rect 18786 48190 18788 48242
rect 18732 48188 18788 48190
rect 17500 45948 17556 46004
rect 17948 47346 18004 47348
rect 17948 47294 17950 47346
rect 17950 47294 18002 47346
rect 18002 47294 18004 47346
rect 17948 47292 18004 47294
rect 18172 47234 18228 47236
rect 18172 47182 18174 47234
rect 18174 47182 18226 47234
rect 18226 47182 18228 47234
rect 18172 47180 18228 47182
rect 17948 45276 18004 45332
rect 17724 45052 17780 45108
rect 17276 44098 17332 44100
rect 17276 44046 17278 44098
rect 17278 44046 17330 44098
rect 17330 44046 17332 44098
rect 17276 44044 17332 44046
rect 17724 44044 17780 44100
rect 18060 45052 18116 45108
rect 18620 45330 18676 45332
rect 18620 45278 18622 45330
rect 18622 45278 18674 45330
rect 18674 45278 18676 45330
rect 18620 45276 18676 45278
rect 18396 45218 18452 45220
rect 18396 45166 18398 45218
rect 18398 45166 18450 45218
rect 18450 45166 18452 45218
rect 18396 45164 18452 45166
rect 18844 45052 18900 45108
rect 18508 44492 18564 44548
rect 18284 44044 18340 44100
rect 18396 44268 18452 44324
rect 18284 43538 18340 43540
rect 18284 43486 18286 43538
rect 18286 43486 18338 43538
rect 18338 43486 18340 43538
rect 18284 43484 18340 43486
rect 18732 44044 18788 44100
rect 18620 43426 18676 43428
rect 18620 43374 18622 43426
rect 18622 43374 18674 43426
rect 18674 43374 18676 43426
rect 18620 43372 18676 43374
rect 18172 42140 18228 42196
rect 17500 41692 17556 41748
rect 17164 40460 17220 40516
rect 16044 39452 16100 39508
rect 14924 38162 14980 38164
rect 14924 38110 14926 38162
rect 14926 38110 14978 38162
rect 14978 38110 14980 38162
rect 14924 38108 14980 38110
rect 17388 39506 17444 39508
rect 17388 39454 17390 39506
rect 17390 39454 17442 39506
rect 17442 39454 17444 39506
rect 17388 39452 17444 39454
rect 17388 39228 17444 39284
rect 16268 38780 16324 38836
rect 17836 38946 17892 38948
rect 17836 38894 17838 38946
rect 17838 38894 17890 38946
rect 17890 38894 17892 38946
rect 17836 38892 17892 38894
rect 14364 35586 14420 35588
rect 14364 35534 14366 35586
rect 14366 35534 14418 35586
rect 14418 35534 14420 35586
rect 14364 35532 14420 35534
rect 13580 34802 13636 34804
rect 13580 34750 13582 34802
rect 13582 34750 13634 34802
rect 13634 34750 13636 34802
rect 13580 34748 13636 34750
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 1708 33122 1764 33124
rect 1708 33070 1710 33122
rect 1710 33070 1762 33122
rect 1762 33070 1764 33122
rect 1708 33068 1764 33070
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 14364 34914 14420 34916
rect 14364 34862 14366 34914
rect 14366 34862 14418 34914
rect 14418 34862 14420 34914
rect 14364 34860 14420 34862
rect 14252 34802 14308 34804
rect 14252 34750 14254 34802
rect 14254 34750 14306 34802
rect 14306 34750 14308 34802
rect 14252 34748 14308 34750
rect 12572 33516 12628 33572
rect 14140 34690 14196 34692
rect 14140 34638 14142 34690
rect 14142 34638 14194 34690
rect 14194 34638 14196 34690
rect 14140 34636 14196 34638
rect 13692 33458 13748 33460
rect 13692 33406 13694 33458
rect 13694 33406 13746 33458
rect 13746 33406 13748 33458
rect 13692 33404 13748 33406
rect 13916 33570 13972 33572
rect 13916 33518 13918 33570
rect 13918 33518 13970 33570
rect 13970 33518 13972 33570
rect 13916 33516 13972 33518
rect 14028 33458 14084 33460
rect 14028 33406 14030 33458
rect 14030 33406 14082 33458
rect 14082 33406 14084 33458
rect 14028 33404 14084 33406
rect 15260 35810 15316 35812
rect 15260 35758 15262 35810
rect 15262 35758 15314 35810
rect 15314 35758 15316 35810
rect 15260 35756 15316 35758
rect 16156 35756 16212 35812
rect 15820 35586 15876 35588
rect 15820 35534 15822 35586
rect 15822 35534 15874 35586
rect 15874 35534 15876 35586
rect 15820 35532 15876 35534
rect 15260 34914 15316 34916
rect 15260 34862 15262 34914
rect 15262 34862 15314 34914
rect 15314 34862 15316 34914
rect 15260 34860 15316 34862
rect 15036 34636 15092 34692
rect 15260 34636 15316 34692
rect 14700 34018 14756 34020
rect 14700 33966 14702 34018
rect 14702 33966 14754 34018
rect 14754 33966 14756 34018
rect 14700 33964 14756 33966
rect 14476 33852 14532 33908
rect 14140 33292 14196 33348
rect 14252 33180 14308 33236
rect 14812 33346 14868 33348
rect 14812 33294 14814 33346
rect 14814 33294 14866 33346
rect 14866 33294 14868 33346
rect 14812 33292 14868 33294
rect 14924 33234 14980 33236
rect 14924 33182 14926 33234
rect 14926 33182 14978 33234
rect 14978 33182 14980 33234
rect 14924 33180 14980 33182
rect 12124 31612 12180 31668
rect 11452 30994 11508 30996
rect 11452 30942 11454 30994
rect 11454 30942 11506 30994
rect 11506 30942 11508 30994
rect 11452 30940 11508 30942
rect 14924 31948 14980 32004
rect 14476 31778 14532 31780
rect 14476 31726 14478 31778
rect 14478 31726 14530 31778
rect 14530 31726 14532 31778
rect 14476 31724 14532 31726
rect 14364 31666 14420 31668
rect 14364 31614 14366 31666
rect 14366 31614 14418 31666
rect 14418 31614 14420 31666
rect 14364 31612 14420 31614
rect 15372 34188 15428 34244
rect 15372 33964 15428 34020
rect 16380 34636 16436 34692
rect 16828 34860 16884 34916
rect 16044 34130 16100 34132
rect 16044 34078 16046 34130
rect 16046 34078 16098 34130
rect 16098 34078 16100 34130
rect 16044 34076 16100 34078
rect 16380 34242 16436 34244
rect 16380 34190 16382 34242
rect 16382 34190 16434 34242
rect 16434 34190 16436 34242
rect 16380 34188 16436 34190
rect 17948 38444 18004 38500
rect 18732 41970 18788 41972
rect 18732 41918 18734 41970
rect 18734 41918 18786 41970
rect 18786 41918 18788 41970
rect 18732 41916 18788 41918
rect 18732 41692 18788 41748
rect 18956 43260 19012 43316
rect 19180 48076 19236 48132
rect 19180 46674 19236 46676
rect 19180 46622 19182 46674
rect 19182 46622 19234 46674
rect 19234 46622 19236 46674
rect 19180 46620 19236 46622
rect 21420 57036 21476 57092
rect 21532 56812 21588 56868
rect 21420 53676 21476 53732
rect 21868 56866 21924 56868
rect 21868 56814 21870 56866
rect 21870 56814 21922 56866
rect 21922 56814 21924 56866
rect 21868 56812 21924 56814
rect 24780 60396 24836 60452
rect 24780 60002 24836 60004
rect 24780 59950 24782 60002
rect 24782 59950 24834 60002
rect 24834 59950 24836 60002
rect 24780 59948 24836 59950
rect 25676 64482 25732 64484
rect 25676 64430 25678 64482
rect 25678 64430 25730 64482
rect 25730 64430 25732 64482
rect 25676 64428 25732 64430
rect 26236 67058 26292 67060
rect 26236 67006 26238 67058
rect 26238 67006 26290 67058
rect 26290 67006 26292 67058
rect 26236 67004 26292 67006
rect 26684 68460 26740 68516
rect 26460 66780 26516 66836
rect 26236 64034 26292 64036
rect 26236 63982 26238 64034
rect 26238 63982 26290 64034
rect 26290 63982 26292 64034
rect 26236 63980 26292 63982
rect 25900 63868 25956 63924
rect 26012 63138 26068 63140
rect 26012 63086 26014 63138
rect 26014 63086 26066 63138
rect 26066 63086 26068 63138
rect 26012 63084 26068 63086
rect 25564 62860 25620 62916
rect 25452 62300 25508 62356
rect 25228 61404 25284 61460
rect 25340 60396 25396 60452
rect 23660 58156 23716 58212
rect 23212 56924 23268 56980
rect 22652 56866 22708 56868
rect 22652 56814 22654 56866
rect 22654 56814 22706 56866
rect 22706 56814 22708 56866
rect 22652 56812 22708 56814
rect 21756 56082 21812 56084
rect 21756 56030 21758 56082
rect 21758 56030 21810 56082
rect 21810 56030 21812 56082
rect 21756 56028 21812 56030
rect 21756 53676 21812 53732
rect 21532 53004 21588 53060
rect 21980 55410 22036 55412
rect 21980 55358 21982 55410
rect 21982 55358 22034 55410
rect 22034 55358 22036 55410
rect 21980 55356 22036 55358
rect 22092 55298 22148 55300
rect 22092 55246 22094 55298
rect 22094 55246 22146 55298
rect 22146 55246 22148 55298
rect 22092 55244 22148 55246
rect 21980 52892 22036 52948
rect 22092 53452 22148 53508
rect 21868 52162 21924 52164
rect 21868 52110 21870 52162
rect 21870 52110 21922 52162
rect 21922 52110 21924 52162
rect 21868 52108 21924 52110
rect 21756 51100 21812 51156
rect 20412 49026 20468 49028
rect 20412 48974 20414 49026
rect 20414 48974 20466 49026
rect 20466 48974 20468 49026
rect 20412 48972 20468 48974
rect 20860 48860 20916 48916
rect 19836 48634 19892 48636
rect 19836 48582 19838 48634
rect 19838 48582 19890 48634
rect 19890 48582 19892 48634
rect 19836 48580 19892 48582
rect 19940 48634 19996 48636
rect 19940 48582 19942 48634
rect 19942 48582 19994 48634
rect 19994 48582 19996 48634
rect 19940 48580 19996 48582
rect 20044 48634 20100 48636
rect 20044 48582 20046 48634
rect 20046 48582 20098 48634
rect 20098 48582 20100 48634
rect 20044 48580 20100 48582
rect 19516 47292 19572 47348
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 20300 48412 20356 48468
rect 21196 48748 21252 48804
rect 20524 48018 20580 48020
rect 20524 47966 20526 48018
rect 20526 47966 20578 48018
rect 20578 47966 20580 48018
rect 20524 47964 20580 47966
rect 20748 47682 20804 47684
rect 20748 47630 20750 47682
rect 20750 47630 20802 47682
rect 20802 47630 20804 47682
rect 20748 47628 20804 47630
rect 20412 47346 20468 47348
rect 20412 47294 20414 47346
rect 20414 47294 20466 47346
rect 20466 47294 20468 47346
rect 20412 47292 20468 47294
rect 20300 47180 20356 47236
rect 19180 44210 19236 44212
rect 19180 44158 19182 44210
rect 19182 44158 19234 44210
rect 19234 44158 19236 44210
rect 19180 44156 19236 44158
rect 19180 41692 19236 41748
rect 19404 44044 19460 44100
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 19964 45276 20020 45332
rect 19852 45106 19908 45108
rect 19852 45054 19854 45106
rect 19854 45054 19906 45106
rect 19906 45054 19908 45106
rect 19852 45052 19908 45054
rect 20188 44882 20244 44884
rect 20188 44830 20190 44882
rect 20190 44830 20242 44882
rect 20242 44830 20244 44882
rect 20188 44828 20244 44830
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 19852 43708 19908 43764
rect 20860 44828 20916 44884
rect 20748 44546 20804 44548
rect 20748 44494 20750 44546
rect 20750 44494 20802 44546
rect 20802 44494 20804 44546
rect 20748 44492 20804 44494
rect 20300 43596 20356 43652
rect 19628 43260 19684 43316
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 19852 42140 19908 42196
rect 19292 41020 19348 41076
rect 19068 40684 19124 40740
rect 19180 40908 19236 40964
rect 18620 40236 18676 40292
rect 18396 39058 18452 39060
rect 18396 39006 18398 39058
rect 18398 39006 18450 39058
rect 18450 39006 18452 39058
rect 18396 39004 18452 39006
rect 18284 38834 18340 38836
rect 18284 38782 18286 38834
rect 18286 38782 18338 38834
rect 18338 38782 18340 38834
rect 18284 38780 18340 38782
rect 18844 38834 18900 38836
rect 18844 38782 18846 38834
rect 18846 38782 18898 38834
rect 18898 38782 18900 38834
rect 18844 38780 18900 38782
rect 19964 41804 20020 41860
rect 19516 40908 19572 40964
rect 19836 40794 19892 40796
rect 19628 40684 19684 40740
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 19628 39900 19684 39956
rect 19516 39788 19572 39844
rect 20188 40626 20244 40628
rect 20188 40574 20190 40626
rect 20190 40574 20242 40626
rect 20242 40574 20244 40626
rect 20188 40572 20244 40574
rect 19852 39788 19908 39844
rect 21644 49810 21700 49812
rect 21644 49758 21646 49810
rect 21646 49758 21698 49810
rect 21698 49758 21700 49810
rect 21644 49756 21700 49758
rect 21420 48860 21476 48916
rect 21756 48802 21812 48804
rect 21756 48750 21758 48802
rect 21758 48750 21810 48802
rect 21810 48750 21812 48802
rect 21756 48748 21812 48750
rect 21532 48242 21588 48244
rect 21532 48190 21534 48242
rect 21534 48190 21586 48242
rect 21586 48190 21588 48242
rect 21532 48188 21588 48190
rect 21868 47068 21924 47124
rect 22764 56028 22820 56084
rect 22204 52834 22260 52836
rect 22204 52782 22206 52834
rect 22206 52782 22258 52834
rect 22258 52782 22260 52834
rect 22204 52780 22260 52782
rect 22316 51996 22372 52052
rect 23100 53564 23156 53620
rect 22428 51378 22484 51380
rect 22428 51326 22430 51378
rect 22430 51326 22482 51378
rect 22482 51326 22484 51378
rect 22428 51324 22484 51326
rect 22428 51100 22484 51156
rect 22652 49922 22708 49924
rect 22652 49870 22654 49922
rect 22654 49870 22706 49922
rect 22706 49870 22708 49922
rect 22652 49868 22708 49870
rect 23100 51490 23156 51492
rect 23100 51438 23102 51490
rect 23102 51438 23154 51490
rect 23154 51438 23156 51490
rect 23100 51436 23156 51438
rect 22764 49756 22820 49812
rect 22316 48242 22372 48244
rect 22316 48190 22318 48242
rect 22318 48190 22370 48242
rect 22370 48190 22372 48242
rect 22316 48188 22372 48190
rect 22876 48860 22932 48916
rect 23660 56476 23716 56532
rect 23884 53676 23940 53732
rect 23772 53004 23828 53060
rect 22764 48412 22820 48468
rect 22764 47628 22820 47684
rect 22204 46956 22260 47012
rect 21644 46114 21700 46116
rect 21644 46062 21646 46114
rect 21646 46062 21698 46114
rect 21698 46062 21700 46114
rect 21644 46060 21700 46062
rect 21644 45836 21700 45892
rect 21420 44492 21476 44548
rect 21420 43650 21476 43652
rect 21420 43598 21422 43650
rect 21422 43598 21474 43650
rect 21474 43598 21476 43650
rect 21420 43596 21476 43598
rect 20636 41916 20692 41972
rect 20636 41692 20692 41748
rect 20076 39788 20132 39844
rect 20636 39788 20692 39844
rect 19068 38946 19124 38948
rect 19068 38894 19070 38946
rect 19070 38894 19122 38946
rect 19122 38894 19124 38946
rect 19068 38892 19124 38894
rect 19180 39228 19236 39284
rect 19180 38444 19236 38500
rect 19404 39452 19460 39508
rect 20300 39618 20356 39620
rect 20300 39566 20302 39618
rect 20302 39566 20354 39618
rect 20354 39566 20356 39618
rect 20300 39564 20356 39566
rect 19852 39452 19908 39508
rect 19740 39394 19796 39396
rect 19740 39342 19742 39394
rect 19742 39342 19794 39394
rect 19794 39342 19796 39394
rect 19740 39340 19796 39342
rect 19836 39226 19892 39228
rect 19628 39116 19684 39172
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 19628 38834 19684 38836
rect 19628 38782 19630 38834
rect 19630 38782 19682 38834
rect 19682 38782 19684 38834
rect 19628 38780 19684 38782
rect 20636 39506 20692 39508
rect 20636 39454 20638 39506
rect 20638 39454 20690 39506
rect 20690 39454 20692 39506
rect 20636 39452 20692 39454
rect 20636 39004 20692 39060
rect 20412 38834 20468 38836
rect 20412 38782 20414 38834
rect 20414 38782 20466 38834
rect 20466 38782 20468 38834
rect 20412 38780 20468 38782
rect 20076 38108 20132 38164
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 20972 40290 21028 40292
rect 20972 40238 20974 40290
rect 20974 40238 21026 40290
rect 21026 40238 21028 40290
rect 20972 40236 21028 40238
rect 22092 46674 22148 46676
rect 22092 46622 22094 46674
rect 22094 46622 22146 46674
rect 22146 46622 22148 46674
rect 22092 46620 22148 46622
rect 21980 45836 22036 45892
rect 22092 45724 22148 45780
rect 22092 45164 22148 45220
rect 21756 44268 21812 44324
rect 21868 43596 21924 43652
rect 21644 42812 21700 42868
rect 21756 41804 21812 41860
rect 22428 46450 22484 46452
rect 22428 46398 22430 46450
rect 22430 46398 22482 46450
rect 22482 46398 22484 46450
rect 22428 46396 22484 46398
rect 22428 46060 22484 46116
rect 22204 43538 22260 43540
rect 22204 43486 22206 43538
rect 22206 43486 22258 43538
rect 22258 43486 22260 43538
rect 22204 43484 22260 43486
rect 22092 41916 22148 41972
rect 22092 41692 22148 41748
rect 21644 41356 21700 41412
rect 21756 41074 21812 41076
rect 21756 41022 21758 41074
rect 21758 41022 21810 41074
rect 21810 41022 21812 41074
rect 21756 41020 21812 41022
rect 21532 40348 21588 40404
rect 21420 40124 21476 40180
rect 21308 39900 21364 39956
rect 21532 39564 21588 39620
rect 21868 40908 21924 40964
rect 21868 40572 21924 40628
rect 21756 40290 21812 40292
rect 21756 40238 21758 40290
rect 21758 40238 21810 40290
rect 21810 40238 21812 40290
rect 21756 40236 21812 40238
rect 21980 40178 22036 40180
rect 21980 40126 21982 40178
rect 21982 40126 22034 40178
rect 22034 40126 22036 40178
rect 21980 40124 22036 40126
rect 23660 48748 23716 48804
rect 23100 47964 23156 48020
rect 22988 45164 23044 45220
rect 23436 44156 23492 44212
rect 22876 43484 22932 43540
rect 22428 43036 22484 43092
rect 22988 43036 23044 43092
rect 22988 42812 23044 42868
rect 22428 41356 22484 41412
rect 22540 41692 22596 41748
rect 22876 42082 22932 42084
rect 22876 42030 22878 42082
rect 22878 42030 22930 42082
rect 22930 42030 22932 42082
rect 22876 42028 22932 42030
rect 22988 41692 23044 41748
rect 22764 41468 22820 41524
rect 22428 40626 22484 40628
rect 22428 40574 22430 40626
rect 22430 40574 22482 40626
rect 22482 40574 22484 40626
rect 22428 40572 22484 40574
rect 23100 40348 23156 40404
rect 22764 40124 22820 40180
rect 22428 39452 22484 39508
rect 20748 38108 20804 38164
rect 22092 38722 22148 38724
rect 22092 38670 22094 38722
rect 22094 38670 22146 38722
rect 22146 38670 22148 38722
rect 22092 38668 22148 38670
rect 22092 38162 22148 38164
rect 22092 38110 22094 38162
rect 22094 38110 22146 38162
rect 22146 38110 22148 38162
rect 22092 38108 22148 38110
rect 21308 37436 21364 37492
rect 19964 37100 20020 37156
rect 17388 34860 17444 34916
rect 16940 34636 16996 34692
rect 16828 34076 16884 34132
rect 16268 33964 16324 34020
rect 16604 34018 16660 34020
rect 16604 33966 16606 34018
rect 16606 33966 16658 34018
rect 16658 33966 16660 34018
rect 16604 33964 16660 33966
rect 15596 33906 15652 33908
rect 15596 33854 15598 33906
rect 15598 33854 15650 33906
rect 15650 33854 15652 33906
rect 15596 33852 15652 33854
rect 17164 33628 17220 33684
rect 15484 33404 15540 33460
rect 15260 31948 15316 32004
rect 17724 33964 17780 34020
rect 19180 33964 19236 34020
rect 19068 33628 19124 33684
rect 17836 33516 17892 33572
rect 18732 33570 18788 33572
rect 18732 33518 18734 33570
rect 18734 33518 18786 33570
rect 18786 33518 18788 33570
rect 18732 33516 18788 33518
rect 16828 33346 16884 33348
rect 16828 33294 16830 33346
rect 16830 33294 16882 33346
rect 16882 33294 16884 33346
rect 16828 33292 16884 33294
rect 18956 33346 19012 33348
rect 18956 33294 18958 33346
rect 18958 33294 19010 33346
rect 19010 33294 19012 33346
rect 18956 33292 19012 33294
rect 15484 31778 15540 31780
rect 15484 31726 15486 31778
rect 15486 31726 15538 31778
rect 15538 31726 15540 31778
rect 15484 31724 15540 31726
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 22988 39618 23044 39620
rect 22988 39566 22990 39618
rect 22990 39566 23042 39618
rect 23042 39566 23044 39618
rect 22988 39564 23044 39566
rect 22764 39452 22820 39508
rect 23548 43148 23604 43204
rect 24108 53004 24164 53060
rect 24220 52892 24276 52948
rect 24444 57650 24500 57652
rect 24444 57598 24446 57650
rect 24446 57598 24498 57650
rect 24498 57598 24500 57650
rect 24444 57596 24500 57598
rect 25676 61404 25732 61460
rect 26236 62972 26292 63028
rect 25900 62412 25956 62468
rect 26796 67058 26852 67060
rect 26796 67006 26798 67058
rect 26798 67006 26850 67058
rect 26850 67006 26852 67058
rect 26796 67004 26852 67006
rect 27580 66892 27636 66948
rect 27356 66834 27412 66836
rect 27356 66782 27358 66834
rect 27358 66782 27410 66834
rect 27410 66782 27412 66834
rect 27356 66780 27412 66782
rect 25676 59948 25732 60004
rect 25900 59106 25956 59108
rect 25900 59054 25902 59106
rect 25902 59054 25954 59106
rect 25954 59054 25956 59106
rect 25900 59052 25956 59054
rect 26572 60620 26628 60676
rect 26460 59052 26516 59108
rect 25564 58546 25620 58548
rect 25564 58494 25566 58546
rect 25566 58494 25618 58546
rect 25618 58494 25620 58546
rect 25564 58492 25620 58494
rect 25676 58434 25732 58436
rect 25676 58382 25678 58434
rect 25678 58382 25730 58434
rect 25730 58382 25732 58434
rect 25676 58380 25732 58382
rect 25564 58210 25620 58212
rect 25564 58158 25566 58210
rect 25566 58158 25618 58210
rect 25618 58158 25620 58210
rect 25564 58156 25620 58158
rect 25116 57372 25172 57428
rect 24780 56754 24836 56756
rect 24780 56702 24782 56754
rect 24782 56702 24834 56754
rect 24834 56702 24836 56754
rect 24780 56700 24836 56702
rect 24444 56476 24500 56532
rect 25116 56476 25172 56532
rect 24556 56194 24612 56196
rect 24556 56142 24558 56194
rect 24558 56142 24610 56194
rect 24610 56142 24612 56194
rect 24556 56140 24612 56142
rect 24444 55244 24500 55300
rect 26236 57036 26292 57092
rect 26348 58716 26404 58772
rect 26348 57372 26404 57428
rect 25676 56924 25732 56980
rect 25676 56642 25732 56644
rect 25676 56590 25678 56642
rect 25678 56590 25730 56642
rect 25730 56590 25732 56642
rect 25676 56588 25732 56590
rect 25788 56476 25844 56532
rect 25900 56082 25956 56084
rect 25900 56030 25902 56082
rect 25902 56030 25954 56082
rect 25954 56030 25956 56082
rect 25900 56028 25956 56030
rect 25788 55858 25844 55860
rect 25788 55806 25790 55858
rect 25790 55806 25842 55858
rect 25842 55806 25844 55858
rect 25788 55804 25844 55806
rect 24444 53452 24500 53508
rect 24444 52050 24500 52052
rect 24444 51998 24446 52050
rect 24446 51998 24498 52050
rect 24498 51998 24500 52050
rect 24444 51996 24500 51998
rect 23996 48412 24052 48468
rect 25340 53564 25396 53620
rect 25228 51772 25284 51828
rect 24668 51378 24724 51380
rect 24668 51326 24670 51378
rect 24670 51326 24722 51378
rect 24722 51326 24724 51378
rect 24668 51324 24724 51326
rect 24556 49868 24612 49924
rect 25900 53676 25956 53732
rect 25676 51490 25732 51492
rect 25676 51438 25678 51490
rect 25678 51438 25730 51490
rect 25730 51438 25732 51490
rect 25676 51436 25732 51438
rect 25228 50428 25284 50484
rect 24220 48748 24276 48804
rect 25004 48412 25060 48468
rect 24108 47516 24164 47572
rect 23996 46956 24052 47012
rect 24108 45778 24164 45780
rect 24108 45726 24110 45778
rect 24110 45726 24162 45778
rect 24162 45726 24164 45778
rect 24108 45724 24164 45726
rect 23660 42812 23716 42868
rect 23548 42028 23604 42084
rect 23436 40962 23492 40964
rect 23436 40910 23438 40962
rect 23438 40910 23490 40962
rect 23490 40910 23492 40962
rect 23436 40908 23492 40910
rect 23324 40514 23380 40516
rect 23324 40462 23326 40514
rect 23326 40462 23378 40514
rect 23378 40462 23380 40514
rect 23324 40460 23380 40462
rect 23212 39116 23268 39172
rect 22652 38050 22708 38052
rect 22652 37998 22654 38050
rect 22654 37998 22706 38050
rect 22706 37998 22708 38050
rect 22652 37996 22708 37998
rect 21868 35868 21924 35924
rect 22540 35922 22596 35924
rect 22540 35870 22542 35922
rect 22542 35870 22594 35922
rect 22594 35870 22596 35922
rect 22540 35868 22596 35870
rect 19292 33404 19348 33460
rect 19628 34690 19684 34692
rect 19628 34638 19630 34690
rect 19630 34638 19682 34690
rect 19682 34638 19684 34690
rect 19628 34636 19684 34638
rect 18620 32450 18676 32452
rect 18620 32398 18622 32450
rect 18622 32398 18674 32450
rect 18674 32398 18676 32450
rect 18620 32396 18676 32398
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 21084 34354 21140 34356
rect 21084 34302 21086 34354
rect 21086 34302 21138 34354
rect 21138 34302 21140 34354
rect 21084 34300 21140 34302
rect 21756 34300 21812 34356
rect 20076 34188 20132 34244
rect 20636 34130 20692 34132
rect 20636 34078 20638 34130
rect 20638 34078 20690 34130
rect 20690 34078 20692 34130
rect 20636 34076 20692 34078
rect 21420 34018 21476 34020
rect 21420 33966 21422 34018
rect 21422 33966 21474 34018
rect 21474 33966 21476 34018
rect 21420 33964 21476 33966
rect 19740 33628 19796 33684
rect 20636 33852 20692 33908
rect 21420 33740 21476 33796
rect 20076 33404 20132 33460
rect 20524 33628 20580 33684
rect 20300 33346 20356 33348
rect 20300 33294 20302 33346
rect 20302 33294 20354 33346
rect 20354 33294 20356 33346
rect 20300 33292 20356 33294
rect 22204 35474 22260 35476
rect 22204 35422 22206 35474
rect 22206 35422 22258 35474
rect 22258 35422 22260 35474
rect 22204 35420 22260 35422
rect 22204 35196 22260 35252
rect 22764 35084 22820 35140
rect 22876 35196 22932 35252
rect 22652 35026 22708 35028
rect 22652 34974 22654 35026
rect 22654 34974 22706 35026
rect 22706 34974 22708 35026
rect 22652 34972 22708 34974
rect 21644 34130 21700 34132
rect 21644 34078 21646 34130
rect 21646 34078 21698 34130
rect 21698 34078 21700 34130
rect 21644 34076 21700 34078
rect 22092 33964 22148 34020
rect 21532 33628 21588 33684
rect 22428 33852 22484 33908
rect 20076 33068 20132 33124
rect 20300 33068 20356 33124
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19628 32396 19684 32452
rect 18620 31836 18676 31892
rect 14700 30994 14756 30996
rect 14700 30942 14702 30994
rect 14702 30942 14754 30994
rect 14754 30942 14756 30994
rect 14700 30940 14756 30942
rect 17500 30994 17556 30996
rect 17500 30942 17502 30994
rect 17502 30942 17554 30994
rect 17554 30942 17556 30994
rect 17500 30940 17556 30942
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 18620 30940 18676 30996
rect 22764 32732 22820 32788
rect 20748 31836 20804 31892
rect 22540 31948 22596 32004
rect 21756 31836 21812 31892
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 23100 35196 23156 35252
rect 23324 39452 23380 39508
rect 24332 43708 24388 43764
rect 24108 41692 24164 41748
rect 24668 48242 24724 48244
rect 24668 48190 24670 48242
rect 24670 48190 24722 48242
rect 24722 48190 24724 48242
rect 24668 48188 24724 48190
rect 24556 47516 24612 47572
rect 26796 63922 26852 63924
rect 26796 63870 26798 63922
rect 26798 63870 26850 63922
rect 26850 63870 26852 63922
rect 26796 63868 26852 63870
rect 35196 69802 35252 69804
rect 35196 69750 35198 69802
rect 35198 69750 35250 69802
rect 35250 69750 35252 69802
rect 35196 69748 35252 69750
rect 35300 69802 35356 69804
rect 35300 69750 35302 69802
rect 35302 69750 35354 69802
rect 35354 69750 35356 69802
rect 35300 69748 35356 69750
rect 35404 69802 35460 69804
rect 35404 69750 35406 69802
rect 35406 69750 35458 69802
rect 35458 69750 35460 69802
rect 35404 69748 35460 69750
rect 28252 68514 28308 68516
rect 28252 68462 28254 68514
rect 28254 68462 28306 68514
rect 28306 68462 28308 68514
rect 28252 68460 28308 68462
rect 28924 68124 28980 68180
rect 35196 68234 35252 68236
rect 35196 68182 35198 68234
rect 35198 68182 35250 68234
rect 35250 68182 35252 68234
rect 35196 68180 35252 68182
rect 35300 68234 35356 68236
rect 35300 68182 35302 68234
rect 35302 68182 35354 68234
rect 35354 68182 35356 68234
rect 35300 68180 35356 68182
rect 35404 68234 35460 68236
rect 35404 68182 35406 68234
rect 35406 68182 35458 68234
rect 35458 68182 35460 68234
rect 35404 68180 35460 68182
rect 28588 66892 28644 66948
rect 35196 66666 35252 66668
rect 35196 66614 35198 66666
rect 35198 66614 35250 66666
rect 35250 66614 35252 66666
rect 35196 66612 35252 66614
rect 35300 66666 35356 66668
rect 35300 66614 35302 66666
rect 35302 66614 35354 66666
rect 35354 66614 35356 66666
rect 35300 66612 35356 66614
rect 35404 66666 35460 66668
rect 35404 66614 35406 66666
rect 35406 66614 35458 66666
rect 35458 66614 35460 66666
rect 35404 66612 35460 66614
rect 35196 65098 35252 65100
rect 35196 65046 35198 65098
rect 35198 65046 35250 65098
rect 35250 65046 35252 65098
rect 35196 65044 35252 65046
rect 35300 65098 35356 65100
rect 35300 65046 35302 65098
rect 35302 65046 35354 65098
rect 35354 65046 35356 65098
rect 35300 65044 35356 65046
rect 35404 65098 35460 65100
rect 35404 65046 35406 65098
rect 35406 65046 35458 65098
rect 35458 65046 35460 65098
rect 35404 65044 35460 65046
rect 28476 63868 28532 63924
rect 26796 62972 26852 63028
rect 26796 62076 26852 62132
rect 27020 62412 27076 62468
rect 27132 58716 27188 58772
rect 38220 63868 38276 63924
rect 29036 62354 29092 62356
rect 29036 62302 29038 62354
rect 29038 62302 29090 62354
rect 29090 62302 29092 62354
rect 29036 62300 29092 62302
rect 35196 63530 35252 63532
rect 35196 63478 35198 63530
rect 35198 63478 35250 63530
rect 35250 63478 35252 63530
rect 35196 63476 35252 63478
rect 35300 63530 35356 63532
rect 35300 63478 35302 63530
rect 35302 63478 35354 63530
rect 35354 63478 35356 63530
rect 35300 63476 35356 63478
rect 35404 63530 35460 63532
rect 35404 63478 35406 63530
rect 35406 63478 35458 63530
rect 35458 63478 35460 63530
rect 35404 63476 35460 63478
rect 29596 62076 29652 62132
rect 35196 61962 35252 61964
rect 35196 61910 35198 61962
rect 35198 61910 35250 61962
rect 35250 61910 35252 61962
rect 35196 61908 35252 61910
rect 35300 61962 35356 61964
rect 35300 61910 35302 61962
rect 35302 61910 35354 61962
rect 35354 61910 35356 61962
rect 35300 61908 35356 61910
rect 35404 61962 35460 61964
rect 35404 61910 35406 61962
rect 35406 61910 35458 61962
rect 35458 61910 35460 61962
rect 35404 61908 35460 61910
rect 27804 60674 27860 60676
rect 27804 60622 27806 60674
rect 27806 60622 27858 60674
rect 27858 60622 27860 60674
rect 27804 60620 27860 60622
rect 35196 60394 35252 60396
rect 35196 60342 35198 60394
rect 35198 60342 35250 60394
rect 35250 60342 35252 60394
rect 35196 60340 35252 60342
rect 35300 60394 35356 60396
rect 35300 60342 35302 60394
rect 35302 60342 35354 60394
rect 35354 60342 35356 60394
rect 35300 60340 35356 60342
rect 35404 60394 35460 60396
rect 35404 60342 35406 60394
rect 35406 60342 35458 60394
rect 35458 60342 35460 60394
rect 35404 60340 35460 60342
rect 35196 58826 35252 58828
rect 35196 58774 35198 58826
rect 35198 58774 35250 58826
rect 35250 58774 35252 58826
rect 35196 58772 35252 58774
rect 35300 58826 35356 58828
rect 35300 58774 35302 58826
rect 35302 58774 35354 58826
rect 35354 58774 35356 58826
rect 35300 58772 35356 58774
rect 35404 58826 35460 58828
rect 35404 58774 35406 58826
rect 35406 58774 35458 58826
rect 35458 58774 35460 58826
rect 35404 58772 35460 58774
rect 26796 57036 26852 57092
rect 27356 56700 27412 56756
rect 26908 56140 26964 56196
rect 27356 55804 27412 55860
rect 27132 53676 27188 53732
rect 26908 53452 26964 53508
rect 26796 53004 26852 53060
rect 27356 53506 27412 53508
rect 27356 53454 27358 53506
rect 27358 53454 27410 53506
rect 27410 53454 27412 53506
rect 27356 53452 27412 53454
rect 27356 52780 27412 52836
rect 26908 51490 26964 51492
rect 26908 51438 26910 51490
rect 26910 51438 26962 51490
rect 26962 51438 26964 51490
rect 26908 51436 26964 51438
rect 26460 48972 26516 49028
rect 26124 48466 26180 48468
rect 26124 48414 26126 48466
rect 26126 48414 26178 48466
rect 26178 48414 26180 48466
rect 26124 48412 26180 48414
rect 25340 48242 25396 48244
rect 25340 48190 25342 48242
rect 25342 48190 25394 48242
rect 25394 48190 25396 48242
rect 25340 48188 25396 48190
rect 25340 47570 25396 47572
rect 25340 47518 25342 47570
rect 25342 47518 25394 47570
rect 25394 47518 25396 47570
rect 25340 47516 25396 47518
rect 26124 46508 26180 46564
rect 25676 46396 25732 46452
rect 24780 44210 24836 44212
rect 24780 44158 24782 44210
rect 24782 44158 24834 44210
rect 24834 44158 24836 44210
rect 24780 44156 24836 44158
rect 24892 43596 24948 43652
rect 25564 45330 25620 45332
rect 25564 45278 25566 45330
rect 25566 45278 25618 45330
rect 25618 45278 25620 45330
rect 25564 45276 25620 45278
rect 25564 43148 25620 43204
rect 24780 41074 24836 41076
rect 24780 41022 24782 41074
rect 24782 41022 24834 41074
rect 24834 41022 24836 41074
rect 24780 41020 24836 41022
rect 23996 40460 24052 40516
rect 23660 38834 23716 38836
rect 23660 38782 23662 38834
rect 23662 38782 23714 38834
rect 23714 38782 23716 38834
rect 23660 38780 23716 38782
rect 24444 38668 24500 38724
rect 24220 38444 24276 38500
rect 24780 38668 24836 38724
rect 24780 38274 24836 38276
rect 24780 38222 24782 38274
rect 24782 38222 24834 38274
rect 24834 38222 24836 38274
rect 24780 38220 24836 38222
rect 23436 35196 23492 35252
rect 24892 37996 24948 38052
rect 24444 35196 24500 35252
rect 25452 41746 25508 41748
rect 25452 41694 25454 41746
rect 25454 41694 25506 41746
rect 25506 41694 25508 41746
rect 25452 41692 25508 41694
rect 25228 41020 25284 41076
rect 26012 45330 26068 45332
rect 26012 45278 26014 45330
rect 26014 45278 26066 45330
rect 26066 45278 26068 45330
rect 26012 45276 26068 45278
rect 26124 42924 26180 42980
rect 26796 48354 26852 48356
rect 26796 48302 26798 48354
rect 26798 48302 26850 48354
rect 26850 48302 26852 48354
rect 26796 48300 26852 48302
rect 26460 48242 26516 48244
rect 26460 48190 26462 48242
rect 26462 48190 26514 48242
rect 26514 48190 26516 48242
rect 26460 48188 26516 48190
rect 25676 41858 25732 41860
rect 25676 41806 25678 41858
rect 25678 41806 25730 41858
rect 25730 41806 25732 41858
rect 25676 41804 25732 41806
rect 25788 40908 25844 40964
rect 25900 41020 25956 41076
rect 25900 40572 25956 40628
rect 25340 39116 25396 39172
rect 25228 38834 25284 38836
rect 25228 38782 25230 38834
rect 25230 38782 25282 38834
rect 25282 38782 25284 38834
rect 25228 38780 25284 38782
rect 26236 41804 26292 41860
rect 26348 41746 26404 41748
rect 26348 41694 26350 41746
rect 26350 41694 26402 41746
rect 26402 41694 26404 41746
rect 26348 41692 26404 41694
rect 26236 40908 26292 40964
rect 26796 43148 26852 43204
rect 26796 42924 26852 42980
rect 25564 38444 25620 38500
rect 26460 38556 26516 38612
rect 25452 38220 25508 38276
rect 25228 36876 25284 36932
rect 25228 35532 25284 35588
rect 25004 34972 25060 35028
rect 25340 35420 25396 35476
rect 24668 34354 24724 34356
rect 24668 34302 24670 34354
rect 24670 34302 24722 34354
rect 24722 34302 24724 34354
rect 24668 34300 24724 34302
rect 26796 41074 26852 41076
rect 26796 41022 26798 41074
rect 26798 41022 26850 41074
rect 26850 41022 26852 41074
rect 26796 41020 26852 41022
rect 27020 49026 27076 49028
rect 27020 48974 27022 49026
rect 27022 48974 27074 49026
rect 27074 48974 27076 49026
rect 27020 48972 27076 48974
rect 27132 48188 27188 48244
rect 27244 48300 27300 48356
rect 27132 47180 27188 47236
rect 27580 56812 27636 56868
rect 28476 57538 28532 57540
rect 28476 57486 28478 57538
rect 28478 57486 28530 57538
rect 28530 57486 28532 57538
rect 28476 57484 28532 57486
rect 28028 57090 28084 57092
rect 28028 57038 28030 57090
rect 28030 57038 28082 57090
rect 28082 57038 28084 57090
rect 28028 57036 28084 57038
rect 28252 56866 28308 56868
rect 28252 56814 28254 56866
rect 28254 56814 28306 56866
rect 28306 56814 28308 56866
rect 28252 56812 28308 56814
rect 27580 56028 27636 56084
rect 28364 55356 28420 55412
rect 35196 57258 35252 57260
rect 35196 57206 35198 57258
rect 35198 57206 35250 57258
rect 35250 57206 35252 57258
rect 35196 57204 35252 57206
rect 35300 57258 35356 57260
rect 35300 57206 35302 57258
rect 35302 57206 35354 57258
rect 35354 57206 35356 57258
rect 35300 57204 35356 57206
rect 35404 57258 35460 57260
rect 35404 57206 35406 57258
rect 35406 57206 35458 57258
rect 35458 57206 35460 57258
rect 35404 57204 35460 57206
rect 29036 56700 29092 56756
rect 29372 56140 29428 56196
rect 29260 55410 29316 55412
rect 29260 55358 29262 55410
rect 29262 55358 29314 55410
rect 29314 55358 29316 55410
rect 29260 55356 29316 55358
rect 29932 56140 29988 56196
rect 35196 55690 35252 55692
rect 35196 55638 35198 55690
rect 35198 55638 35250 55690
rect 35250 55638 35252 55690
rect 35196 55636 35252 55638
rect 35300 55690 35356 55692
rect 35300 55638 35302 55690
rect 35302 55638 35354 55690
rect 35354 55638 35356 55690
rect 35300 55636 35356 55638
rect 35404 55690 35460 55692
rect 35404 55638 35406 55690
rect 35406 55638 35458 55690
rect 35458 55638 35460 55690
rect 35404 55636 35460 55638
rect 29596 55298 29652 55300
rect 29596 55246 29598 55298
rect 29598 55246 29650 55298
rect 29650 55246 29652 55298
rect 29596 55244 29652 55246
rect 35196 54122 35252 54124
rect 35196 54070 35198 54122
rect 35198 54070 35250 54122
rect 35250 54070 35252 54122
rect 35196 54068 35252 54070
rect 35300 54122 35356 54124
rect 35300 54070 35302 54122
rect 35302 54070 35354 54122
rect 35354 54070 35356 54122
rect 35300 54068 35356 54070
rect 35404 54122 35460 54124
rect 35404 54070 35406 54122
rect 35406 54070 35458 54122
rect 35458 54070 35460 54122
rect 35404 54068 35460 54070
rect 28476 53676 28532 53732
rect 28476 52892 28532 52948
rect 33068 52946 33124 52948
rect 33068 52894 33070 52946
rect 33070 52894 33122 52946
rect 33122 52894 33124 52946
rect 33068 52892 33124 52894
rect 28700 52834 28756 52836
rect 28700 52782 28702 52834
rect 28702 52782 28754 52834
rect 28754 52782 28756 52834
rect 28700 52780 28756 52782
rect 32956 52108 33012 52164
rect 33740 52162 33796 52164
rect 33740 52110 33742 52162
rect 33742 52110 33794 52162
rect 33794 52110 33796 52162
rect 33740 52108 33796 52110
rect 37996 53116 38052 53172
rect 35196 52554 35252 52556
rect 35196 52502 35198 52554
rect 35198 52502 35250 52554
rect 35250 52502 35252 52554
rect 35196 52500 35252 52502
rect 35300 52554 35356 52556
rect 35300 52502 35302 52554
rect 35302 52502 35354 52554
rect 35354 52502 35356 52554
rect 35300 52500 35356 52502
rect 35404 52554 35460 52556
rect 35404 52502 35406 52554
rect 35406 52502 35458 52554
rect 35458 52502 35460 52554
rect 35404 52500 35460 52502
rect 35196 50986 35252 50988
rect 35196 50934 35198 50986
rect 35198 50934 35250 50986
rect 35250 50934 35252 50986
rect 35196 50932 35252 50934
rect 35300 50986 35356 50988
rect 35300 50934 35302 50986
rect 35302 50934 35354 50986
rect 35354 50934 35356 50986
rect 35300 50932 35356 50934
rect 35404 50986 35460 50988
rect 35404 50934 35406 50986
rect 35406 50934 35458 50986
rect 35458 50934 35460 50986
rect 35404 50932 35460 50934
rect 27468 48354 27524 48356
rect 27468 48302 27470 48354
rect 27470 48302 27522 48354
rect 27522 48302 27524 48354
rect 27468 48300 27524 48302
rect 27356 46562 27412 46564
rect 27356 46510 27358 46562
rect 27358 46510 27410 46562
rect 27410 46510 27412 46562
rect 27356 46508 27412 46510
rect 27580 45276 27636 45332
rect 27916 48972 27972 49028
rect 28028 48130 28084 48132
rect 28028 48078 28030 48130
rect 28030 48078 28082 48130
rect 28082 48078 28084 48130
rect 28028 48076 28084 48078
rect 30492 49698 30548 49700
rect 30492 49646 30494 49698
rect 30494 49646 30546 49698
rect 30546 49646 30548 49698
rect 30492 49644 30548 49646
rect 29148 49138 29204 49140
rect 29148 49086 29150 49138
rect 29150 49086 29202 49138
rect 29202 49086 29204 49138
rect 29148 49084 29204 49086
rect 30268 49084 30324 49140
rect 29932 48076 29988 48132
rect 28364 47068 28420 47124
rect 29260 47068 29316 47124
rect 28588 46060 28644 46116
rect 27020 39116 27076 39172
rect 27020 38668 27076 38724
rect 26012 38274 26068 38276
rect 26012 38222 26014 38274
rect 26014 38222 26066 38274
rect 26066 38222 26068 38274
rect 26012 38220 26068 38222
rect 26236 38050 26292 38052
rect 26236 37998 26238 38050
rect 26238 37998 26290 38050
rect 26290 37998 26292 38050
rect 26236 37996 26292 37998
rect 26460 37378 26516 37380
rect 26460 37326 26462 37378
rect 26462 37326 26514 37378
rect 26514 37326 26516 37378
rect 26460 37324 26516 37326
rect 26684 37996 26740 38052
rect 26908 38274 26964 38276
rect 26908 38222 26910 38274
rect 26910 38222 26962 38274
rect 26962 38222 26964 38274
rect 26908 38220 26964 38222
rect 26796 36876 26852 36932
rect 26908 36988 26964 37044
rect 25452 34300 25508 34356
rect 25564 35084 25620 35140
rect 24668 33740 24724 33796
rect 23548 32732 23604 32788
rect 24220 32786 24276 32788
rect 24220 32734 24222 32786
rect 24222 32734 24274 32786
rect 24274 32734 24276 32786
rect 24220 32732 24276 32734
rect 23212 32562 23268 32564
rect 23212 32510 23214 32562
rect 23214 32510 23266 32562
rect 23266 32510 23268 32562
rect 23212 32508 23268 32510
rect 24332 32562 24388 32564
rect 24332 32510 24334 32562
rect 24334 32510 24386 32562
rect 24386 32510 24388 32562
rect 24332 32508 24388 32510
rect 23212 31948 23268 32004
rect 26348 33404 26404 33460
rect 26796 33458 26852 33460
rect 26796 33406 26798 33458
rect 26798 33406 26850 33458
rect 26850 33406 26852 33458
rect 26796 33404 26852 33406
rect 26124 33122 26180 33124
rect 26124 33070 26126 33122
rect 26126 33070 26178 33122
rect 26178 33070 26180 33122
rect 26124 33068 26180 33070
rect 25452 31948 25508 32004
rect 26236 31948 26292 32004
rect 24668 30994 24724 30996
rect 24668 30942 24670 30994
rect 24670 30942 24722 30994
rect 24722 30942 24724 30994
rect 24668 30940 24724 30942
rect 25228 30994 25284 30996
rect 25228 30942 25230 30994
rect 25230 30942 25282 30994
rect 25282 30942 25284 30994
rect 25228 30940 25284 30942
rect 26348 32508 26404 32564
rect 27132 38556 27188 38612
rect 27132 36652 27188 36708
rect 27132 35196 27188 35252
rect 27468 43650 27524 43652
rect 27468 43598 27470 43650
rect 27470 43598 27522 43650
rect 27522 43598 27524 43650
rect 27468 43596 27524 43598
rect 27580 42924 27636 42980
rect 27804 41244 27860 41300
rect 27804 41020 27860 41076
rect 28028 43596 28084 43652
rect 30156 46620 30212 46676
rect 29932 46060 29988 46116
rect 28700 43538 28756 43540
rect 28700 43486 28702 43538
rect 28702 43486 28754 43538
rect 28754 43486 28756 43538
rect 28700 43484 28756 43486
rect 28140 42812 28196 42868
rect 29596 43708 29652 43764
rect 28700 42924 28756 42980
rect 29260 42700 29316 42756
rect 28364 42588 28420 42644
rect 28252 42140 28308 42196
rect 28476 42028 28532 42084
rect 28924 42252 28980 42308
rect 28364 41468 28420 41524
rect 29148 42028 29204 42084
rect 28364 41074 28420 41076
rect 28364 41022 28366 41074
rect 28366 41022 28418 41074
rect 28418 41022 28420 41074
rect 28364 41020 28420 41022
rect 29596 42924 29652 42980
rect 29484 42588 29540 42644
rect 29372 42364 29428 42420
rect 29596 42476 29652 42532
rect 29372 41692 29428 41748
rect 29484 41468 29540 41524
rect 29260 40684 29316 40740
rect 28476 40572 28532 40628
rect 27692 38108 27748 38164
rect 27356 37324 27412 37380
rect 27356 36204 27412 36260
rect 27580 36652 27636 36708
rect 28028 38220 28084 38276
rect 29820 42252 29876 42308
rect 32396 49644 32452 49700
rect 32396 49138 32452 49140
rect 32396 49086 32398 49138
rect 32398 49086 32450 49138
rect 32450 49086 32452 49138
rect 32396 49084 32452 49086
rect 31164 48972 31220 49028
rect 31948 49026 32004 49028
rect 31948 48974 31950 49026
rect 31950 48974 32002 49026
rect 32002 48974 32004 49026
rect 31948 48972 32004 48974
rect 31276 48300 31332 48356
rect 32060 48860 32116 48916
rect 31836 48242 31892 48244
rect 31836 48190 31838 48242
rect 31838 48190 31890 48242
rect 31890 48190 31892 48242
rect 31836 48188 31892 48190
rect 31836 47852 31892 47908
rect 31500 47180 31556 47236
rect 30828 45218 30884 45220
rect 30828 45166 30830 45218
rect 30830 45166 30882 45218
rect 30882 45166 30884 45218
rect 30828 45164 30884 45166
rect 30044 43538 30100 43540
rect 30044 43486 30046 43538
rect 30046 43486 30098 43538
rect 30098 43486 30100 43538
rect 30044 43484 30100 43486
rect 30044 42252 30100 42308
rect 30268 42812 30324 42868
rect 30604 42754 30660 42756
rect 30604 42702 30606 42754
rect 30606 42702 30658 42754
rect 30658 42702 30660 42754
rect 30604 42700 30660 42702
rect 29932 42140 29988 42196
rect 29708 42028 29764 42084
rect 30044 41580 30100 41636
rect 30044 41020 30100 41076
rect 30380 41804 30436 41860
rect 31724 46786 31780 46788
rect 31724 46734 31726 46786
rect 31726 46734 31778 46786
rect 31778 46734 31780 46786
rect 31724 46732 31780 46734
rect 31612 46674 31668 46676
rect 31612 46622 31614 46674
rect 31614 46622 31666 46674
rect 31666 46622 31668 46674
rect 31612 46620 31668 46622
rect 32508 48466 32564 48468
rect 32508 48414 32510 48466
rect 32510 48414 32562 48466
rect 32562 48414 32564 48466
rect 32508 48412 32564 48414
rect 32396 48300 32452 48356
rect 31948 46786 32004 46788
rect 31948 46734 31950 46786
rect 31950 46734 32002 46786
rect 32002 46734 32004 46786
rect 31948 46732 32004 46734
rect 32620 48188 32676 48244
rect 32956 47740 33012 47796
rect 33292 49084 33348 49140
rect 36764 49756 36820 49812
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 34860 48972 34916 49028
rect 35084 49026 35140 49028
rect 35084 48974 35086 49026
rect 35086 48974 35138 49026
rect 35138 48974 35140 49026
rect 35084 48972 35140 48974
rect 35420 49026 35476 49028
rect 35420 48974 35422 49026
rect 35422 48974 35474 49026
rect 35474 48974 35476 49026
rect 35420 48972 35476 48974
rect 34412 48914 34468 48916
rect 34412 48862 34414 48914
rect 34414 48862 34466 48914
rect 34466 48862 34468 48914
rect 34412 48860 34468 48862
rect 35980 48860 36036 48916
rect 33740 48802 33796 48804
rect 33740 48750 33742 48802
rect 33742 48750 33794 48802
rect 33794 48750 33796 48802
rect 33740 48748 33796 48750
rect 34524 48748 34580 48804
rect 33516 48300 33572 48356
rect 33180 47852 33236 47908
rect 34076 47852 34132 47908
rect 32956 46732 33012 46788
rect 33180 47404 33236 47460
rect 31612 45164 31668 45220
rect 32508 46674 32564 46676
rect 32508 46622 32510 46674
rect 32510 46622 32562 46674
rect 32562 46622 32564 46674
rect 32508 46620 32564 46622
rect 31948 44994 32004 44996
rect 31948 44942 31950 44994
rect 31950 44942 32002 44994
rect 32002 44942 32004 44994
rect 31948 44940 32004 44942
rect 31388 43484 31444 43540
rect 30940 42530 30996 42532
rect 30940 42478 30942 42530
rect 30942 42478 30994 42530
rect 30994 42478 30996 42530
rect 30940 42476 30996 42478
rect 30828 41916 30884 41972
rect 30716 41356 30772 41412
rect 30492 40572 30548 40628
rect 30716 41020 30772 41076
rect 30604 40402 30660 40404
rect 30604 40350 30606 40402
rect 30606 40350 30658 40402
rect 30658 40350 30660 40402
rect 30604 40348 30660 40350
rect 29596 39730 29652 39732
rect 29596 39678 29598 39730
rect 29598 39678 29650 39730
rect 29650 39678 29652 39730
rect 29596 39676 29652 39678
rect 31052 41580 31108 41636
rect 31276 42642 31332 42644
rect 31276 42590 31278 42642
rect 31278 42590 31330 42642
rect 31330 42590 31332 42642
rect 31276 42588 31332 42590
rect 31276 42364 31332 42420
rect 31276 42140 31332 42196
rect 31724 42866 31780 42868
rect 31724 42814 31726 42866
rect 31726 42814 31778 42866
rect 31778 42814 31780 42866
rect 31724 42812 31780 42814
rect 31612 42642 31668 42644
rect 31612 42590 31614 42642
rect 31614 42590 31666 42642
rect 31666 42590 31668 42642
rect 31612 42588 31668 42590
rect 32060 43148 32116 43204
rect 32396 46396 32452 46452
rect 31836 42140 31892 42196
rect 31948 42700 32004 42756
rect 32284 46060 32340 46116
rect 32396 45106 32452 45108
rect 32396 45054 32398 45106
rect 32398 45054 32450 45106
rect 32450 45054 32452 45106
rect 32396 45052 32452 45054
rect 32172 42588 32228 42644
rect 33292 46396 33348 46452
rect 33292 45276 33348 45332
rect 33180 45164 33236 45220
rect 33292 45106 33348 45108
rect 33292 45054 33294 45106
rect 33294 45054 33346 45106
rect 33346 45054 33348 45106
rect 33292 45052 33348 45054
rect 34300 47740 34356 47796
rect 33740 46674 33796 46676
rect 33740 46622 33742 46674
rect 33742 46622 33794 46674
rect 33794 46622 33796 46674
rect 33740 46620 33796 46622
rect 34860 48802 34916 48804
rect 34860 48750 34862 48802
rect 34862 48750 34914 48802
rect 34914 48750 34916 48802
rect 34860 48748 34916 48750
rect 34748 47628 34804 47684
rect 34412 45276 34468 45332
rect 34076 45164 34132 45220
rect 34300 45106 34356 45108
rect 34300 45054 34302 45106
rect 34302 45054 34354 45106
rect 34354 45054 34356 45106
rect 34300 45052 34356 45054
rect 33180 44940 33236 44996
rect 31388 41298 31444 41300
rect 31388 41246 31390 41298
rect 31390 41246 31442 41298
rect 31442 41246 31444 41298
rect 31388 41244 31444 41246
rect 31724 41356 31780 41412
rect 31836 41468 31892 41524
rect 31052 40908 31108 40964
rect 31500 40962 31556 40964
rect 31500 40910 31502 40962
rect 31502 40910 31554 40962
rect 31554 40910 31556 40962
rect 31500 40908 31556 40910
rect 31388 40796 31444 40852
rect 30940 40572 30996 40628
rect 31948 41020 32004 41076
rect 32060 40908 32116 40964
rect 31836 40796 31892 40852
rect 32060 40402 32116 40404
rect 32060 40350 32062 40402
rect 32062 40350 32114 40402
rect 32114 40350 32116 40402
rect 32060 40348 32116 40350
rect 30828 39676 30884 39732
rect 32284 42252 32340 42308
rect 33180 42700 33236 42756
rect 33292 43484 33348 43540
rect 34748 46396 34804 46452
rect 34748 44882 34804 44884
rect 34748 44830 34750 44882
rect 34750 44830 34802 44882
rect 34802 44830 34804 44882
rect 34748 44828 34804 44830
rect 35644 48802 35700 48804
rect 35644 48750 35646 48802
rect 35646 48750 35698 48802
rect 35698 48750 35700 48802
rect 35644 48748 35700 48750
rect 34972 44940 35028 44996
rect 35084 48636 35140 48692
rect 35868 48412 35924 48468
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 36092 47628 36148 47684
rect 36876 47068 36932 47124
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 33404 42754 33460 42756
rect 33404 42702 33406 42754
rect 33406 42702 33458 42754
rect 33458 42702 33460 42754
rect 33404 42700 33460 42702
rect 32396 41692 32452 41748
rect 32620 42252 32676 42308
rect 32844 42364 32900 42420
rect 32956 42588 33012 42644
rect 33180 42530 33236 42532
rect 33180 42478 33182 42530
rect 33182 42478 33234 42530
rect 33234 42478 33236 42530
rect 33180 42476 33236 42478
rect 33292 42364 33348 42420
rect 32732 42140 32788 42196
rect 33964 43538 34020 43540
rect 33964 43486 33966 43538
rect 33966 43486 34018 43538
rect 34018 43486 34020 43538
rect 33964 43484 34020 43486
rect 33516 41916 33572 41972
rect 32956 41804 33012 41860
rect 33180 41692 33236 41748
rect 33964 41916 34020 41972
rect 34076 42476 34132 42532
rect 33740 41804 33796 41860
rect 33628 41692 33684 41748
rect 32956 40962 33012 40964
rect 32956 40910 32958 40962
rect 32958 40910 33010 40962
rect 33010 40910 33012 40962
rect 32956 40908 33012 40910
rect 32508 40796 32564 40852
rect 32396 40684 32452 40740
rect 36428 44940 36484 44996
rect 38220 44994 38276 44996
rect 38220 44942 38222 44994
rect 38222 44942 38274 44994
rect 38274 44942 38276 44994
rect 38220 44940 38276 44942
rect 36092 44828 36148 44884
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 34748 42700 34804 42756
rect 34636 42140 34692 42196
rect 34636 41970 34692 41972
rect 34636 41918 34638 41970
rect 34638 41918 34690 41970
rect 34690 41918 34692 41970
rect 34636 41916 34692 41918
rect 35420 42530 35476 42532
rect 35420 42478 35422 42530
rect 35422 42478 35474 42530
rect 35474 42478 35476 42530
rect 35420 42476 35476 42478
rect 36092 42140 36148 42196
rect 36316 42252 36372 42308
rect 36092 41858 36148 41860
rect 36092 41806 36094 41858
rect 36094 41806 36146 41858
rect 36146 41806 36148 41858
rect 36092 41804 36148 41806
rect 34972 41692 35028 41748
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 38220 42252 38276 42308
rect 36428 41804 36484 41860
rect 38220 41858 38276 41860
rect 38220 41806 38222 41858
rect 38222 41806 38274 41858
rect 38274 41806 38276 41858
rect 38220 41804 38276 41806
rect 34188 40908 34244 40964
rect 35980 40348 36036 40404
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 34972 39004 35028 39060
rect 32396 38556 32452 38612
rect 33404 38556 33460 38612
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 32396 38108 32452 38164
rect 27692 36988 27748 37044
rect 28028 36258 28084 36260
rect 28028 36206 28030 36258
rect 28030 36206 28082 36258
rect 28082 36206 28084 36258
rect 28028 36204 28084 36206
rect 27244 33404 27300 33460
rect 27468 33068 27524 33124
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 38220 36370 38276 36372
rect 38220 36318 38222 36370
rect 38222 36318 38274 36370
rect 38274 36318 38276 36370
rect 38220 36316 38276 36318
rect 28924 36204 28980 36260
rect 29820 36204 29876 36260
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 28140 32562 28196 32564
rect 28140 32510 28142 32562
rect 28142 32510 28194 32562
rect 28194 32510 28196 32562
rect 28140 32508 28196 32510
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 27020 30940 27076 30996
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 23212 30268 23268 30324
rect 24220 30322 24276 30324
rect 24220 30270 24222 30322
rect 24222 30270 24274 30322
rect 24274 30270 24276 30322
rect 24220 30268 24276 30270
rect 38220 30268 38276 30324
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 38220 22876 38276 22932
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
<< metal3 >>
rect 4466 96404 4476 96460
rect 4532 96404 4580 96460
rect 4636 96404 4684 96460
rect 4740 96404 4750 96460
rect 35186 96404 35196 96460
rect 35252 96404 35300 96460
rect 35356 96404 35404 96460
rect 35460 96404 35470 96460
rect 19826 95620 19836 95676
rect 19892 95620 19940 95676
rect 19996 95620 20044 95676
rect 20100 95620 20110 95676
rect 4466 94836 4476 94892
rect 4532 94836 4580 94892
rect 4636 94836 4684 94892
rect 4740 94836 4750 94892
rect 35186 94836 35196 94892
rect 35252 94836 35300 94892
rect 35356 94836 35404 94892
rect 35460 94836 35470 94892
rect 19826 94052 19836 94108
rect 19892 94052 19940 94108
rect 19996 94052 20044 94108
rect 20100 94052 20110 94108
rect 4466 93268 4476 93324
rect 4532 93268 4580 93324
rect 4636 93268 4684 93324
rect 4740 93268 4750 93324
rect 35186 93268 35196 93324
rect 35252 93268 35300 93324
rect 35356 93268 35404 93324
rect 35460 93268 35470 93324
rect 19826 92484 19836 92540
rect 19892 92484 19940 92540
rect 19996 92484 20044 92540
rect 20100 92484 20110 92540
rect 4466 91700 4476 91756
rect 4532 91700 4580 91756
rect 4636 91700 4684 91756
rect 4740 91700 4750 91756
rect 35186 91700 35196 91756
rect 35252 91700 35300 91756
rect 35356 91700 35404 91756
rect 35460 91700 35470 91756
rect 19826 90916 19836 90972
rect 19892 90916 19940 90972
rect 19996 90916 20044 90972
rect 20100 90916 20110 90972
rect 4466 90132 4476 90188
rect 4532 90132 4580 90188
rect 4636 90132 4684 90188
rect 4740 90132 4750 90188
rect 35186 90132 35196 90188
rect 35252 90132 35300 90188
rect 35356 90132 35404 90188
rect 35460 90132 35470 90188
rect 19826 89348 19836 89404
rect 19892 89348 19940 89404
rect 19996 89348 20044 89404
rect 20100 89348 20110 89404
rect 4466 88564 4476 88620
rect 4532 88564 4580 88620
rect 4636 88564 4684 88620
rect 4740 88564 4750 88620
rect 35186 88564 35196 88620
rect 35252 88564 35300 88620
rect 35356 88564 35404 88620
rect 35460 88564 35470 88620
rect 19826 87780 19836 87836
rect 19892 87780 19940 87836
rect 19996 87780 20044 87836
rect 20100 87780 20110 87836
rect 4466 86996 4476 87052
rect 4532 86996 4580 87052
rect 4636 86996 4684 87052
rect 4740 86996 4750 87052
rect 35186 86996 35196 87052
rect 35252 86996 35300 87052
rect 35356 86996 35404 87052
rect 35460 86996 35470 87052
rect 19826 86212 19836 86268
rect 19892 86212 19940 86268
rect 19996 86212 20044 86268
rect 20100 86212 20110 86268
rect 4466 85428 4476 85484
rect 4532 85428 4580 85484
rect 4636 85428 4684 85484
rect 4740 85428 4750 85484
rect 35186 85428 35196 85484
rect 35252 85428 35300 85484
rect 35356 85428 35404 85484
rect 35460 85428 35470 85484
rect 19826 84644 19836 84700
rect 19892 84644 19940 84700
rect 19996 84644 20044 84700
rect 20100 84644 20110 84700
rect 4466 83860 4476 83916
rect 4532 83860 4580 83916
rect 4636 83860 4684 83916
rect 4740 83860 4750 83916
rect 35186 83860 35196 83916
rect 35252 83860 35300 83916
rect 35356 83860 35404 83916
rect 35460 83860 35470 83916
rect 19826 83076 19836 83132
rect 19892 83076 19940 83132
rect 19996 83076 20044 83132
rect 20100 83076 20110 83132
rect 4466 82292 4476 82348
rect 4532 82292 4580 82348
rect 4636 82292 4684 82348
rect 4740 82292 4750 82348
rect 35186 82292 35196 82348
rect 35252 82292 35300 82348
rect 35356 82292 35404 82348
rect 35460 82292 35470 82348
rect 19826 81508 19836 81564
rect 19892 81508 19940 81564
rect 19996 81508 20044 81564
rect 20100 81508 20110 81564
rect 4466 80724 4476 80780
rect 4532 80724 4580 80780
rect 4636 80724 4684 80780
rect 4740 80724 4750 80780
rect 35186 80724 35196 80780
rect 35252 80724 35300 80780
rect 35356 80724 35404 80780
rect 35460 80724 35470 80780
rect 19826 79940 19836 79996
rect 19892 79940 19940 79996
rect 19996 79940 20044 79996
rect 20100 79940 20110 79996
rect 4466 79156 4476 79212
rect 4532 79156 4580 79212
rect 4636 79156 4684 79212
rect 4740 79156 4750 79212
rect 35186 79156 35196 79212
rect 35252 79156 35300 79212
rect 35356 79156 35404 79212
rect 35460 79156 35470 79212
rect 19826 78372 19836 78428
rect 19892 78372 19940 78428
rect 19996 78372 20044 78428
rect 20100 78372 20110 78428
rect 4466 77588 4476 77644
rect 4532 77588 4580 77644
rect 4636 77588 4684 77644
rect 4740 77588 4750 77644
rect 35186 77588 35196 77644
rect 35252 77588 35300 77644
rect 35356 77588 35404 77644
rect 35460 77588 35470 77644
rect 19826 76804 19836 76860
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 20100 76804 20110 76860
rect 4466 76020 4476 76076
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4740 76020 4750 76076
rect 35186 76020 35196 76076
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35460 76020 35470 76076
rect 19826 75236 19836 75292
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 20100 75236 20110 75292
rect 4466 74452 4476 74508
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4740 74452 4750 74508
rect 35186 74452 35196 74508
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35460 74452 35470 74508
rect 19826 73668 19836 73724
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 20100 73668 20110 73724
rect 4466 72884 4476 72940
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4740 72884 4750 72940
rect 35186 72884 35196 72940
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35460 72884 35470 72940
rect 19826 72100 19836 72156
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 20100 72100 20110 72156
rect 4466 71316 4476 71372
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4740 71316 4750 71372
rect 35186 71316 35196 71372
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35460 71316 35470 71372
rect 19826 70532 19836 70588
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 20100 70532 20110 70588
rect 25554 70028 25564 70084
rect 25620 70028 26124 70084
rect 26180 70028 27692 70084
rect 27748 70028 27758 70084
rect 24434 69916 24444 69972
rect 24500 69916 25228 69972
rect 25284 69916 25294 69972
rect 4466 69748 4476 69804
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4740 69748 4750 69804
rect 35186 69748 35196 69804
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35460 69748 35470 69804
rect 19506 69580 19516 69636
rect 19572 69580 19852 69636
rect 19908 69580 20636 69636
rect 20692 69580 20702 69636
rect 20066 69468 20076 69524
rect 20132 69468 20412 69524
rect 20468 69468 22316 69524
rect 22372 69468 23548 69524
rect 23604 69468 23614 69524
rect 13010 69356 13020 69412
rect 13076 69356 15260 69412
rect 15316 69356 17612 69412
rect 17668 69356 18172 69412
rect 18228 69356 18238 69412
rect 19826 68964 19836 69020
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 20100 68964 20110 69020
rect 19618 68796 19628 68852
rect 19684 68796 20412 68852
rect 20468 68796 20478 68852
rect 24444 68796 25228 68852
rect 25284 68796 26124 68852
rect 26180 68796 26190 68852
rect 24444 68740 24500 68796
rect 2034 68684 2044 68740
rect 2100 68684 9660 68740
rect 9716 68684 9726 68740
rect 20132 68684 24500 68740
rect 24658 68684 24668 68740
rect 24724 68684 25788 68740
rect 25844 68684 25854 68740
rect 20132 68628 20188 68684
rect 8306 68572 8316 68628
rect 8372 68572 9772 68628
rect 9828 68572 9838 68628
rect 18946 68572 18956 68628
rect 19012 68572 20188 68628
rect 1698 68460 1708 68516
rect 1764 68460 2492 68516
rect 2548 68460 2558 68516
rect 13234 68460 13244 68516
rect 13300 68460 15820 68516
rect 15876 68460 15886 68516
rect 17714 68460 17724 68516
rect 17780 68460 19628 68516
rect 19684 68460 19694 68516
rect 20514 68460 20524 68516
rect 20580 68460 21084 68516
rect 21140 68460 24332 68516
rect 24388 68460 24398 68516
rect 24658 68460 24668 68516
rect 24724 68460 25452 68516
rect 25508 68460 25518 68516
rect 26674 68460 26684 68516
rect 26740 68460 28252 68516
rect 28308 68460 28318 68516
rect 9762 68348 9772 68404
rect 9828 68348 11788 68404
rect 11844 68348 11854 68404
rect 17602 68348 17612 68404
rect 17668 68348 20076 68404
rect 20132 68348 20142 68404
rect 4466 68180 4476 68236
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4740 68180 4750 68236
rect 35186 68180 35196 68236
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35460 68180 35470 68236
rect 23986 68124 23996 68180
rect 24052 68124 25116 68180
rect 25172 68124 25788 68180
rect 25844 68124 28924 68180
rect 28980 68124 28990 68180
rect 0 67956 800 67984
rect 0 67900 1708 67956
rect 1764 67900 1774 67956
rect 7634 67900 7644 67956
rect 7700 67900 8764 67956
rect 8820 67900 16716 67956
rect 16772 67900 17388 67956
rect 17444 67900 17836 67956
rect 17892 67900 17902 67956
rect 24546 67900 24556 67956
rect 24612 67900 25452 67956
rect 25508 67900 25518 67956
rect 0 67872 800 67900
rect 14130 67788 14140 67844
rect 14196 67788 15484 67844
rect 15540 67788 15550 67844
rect 15810 67788 15820 67844
rect 15876 67788 17724 67844
rect 17780 67788 17790 67844
rect 10098 67676 10108 67732
rect 10164 67676 11452 67732
rect 11508 67676 12348 67732
rect 12404 67676 12414 67732
rect 12898 67676 12908 67732
rect 12964 67676 14476 67732
rect 14532 67676 15148 67732
rect 16594 67676 16604 67732
rect 16660 67676 18172 67732
rect 18228 67676 18238 67732
rect 23874 67676 23884 67732
rect 23940 67676 24668 67732
rect 24724 67676 24734 67732
rect 15092 67620 15148 67676
rect 12786 67564 12796 67620
rect 12852 67564 13580 67620
rect 13636 67564 13646 67620
rect 15092 67564 17948 67620
rect 18004 67564 18508 67620
rect 18564 67564 18574 67620
rect 19826 67396 19836 67452
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 20100 67396 20110 67452
rect 2034 67340 2044 67396
rect 2100 67340 8204 67396
rect 8260 67340 8270 67396
rect 0 67284 800 67312
rect 0 67228 1708 67284
rect 1764 67228 2492 67284
rect 2548 67228 2558 67284
rect 0 67200 800 67228
rect 2034 67116 2044 67172
rect 2100 67116 9884 67172
rect 9940 67116 9950 67172
rect 8642 67004 8652 67060
rect 8708 67004 9436 67060
rect 9492 67004 9502 67060
rect 23538 67004 23548 67060
rect 23604 67004 25228 67060
rect 25284 67004 25294 67060
rect 25666 67004 25676 67060
rect 25732 67004 26236 67060
rect 26292 67004 26796 67060
rect 26852 67004 26862 67060
rect 18386 66892 18396 66948
rect 18452 66892 25788 66948
rect 25844 66892 27580 66948
rect 27636 66892 28588 66948
rect 28644 66892 28654 66948
rect 13906 66780 13916 66836
rect 13972 66780 16716 66836
rect 16772 66780 19516 66836
rect 19572 66780 19582 66836
rect 26450 66780 26460 66836
rect 26516 66780 27356 66836
rect 27412 66780 27422 66836
rect 0 66612 800 66640
rect 4466 66612 4476 66668
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4740 66612 4750 66668
rect 35186 66612 35196 66668
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35460 66612 35470 66668
rect 0 66556 1708 66612
rect 1764 66556 2492 66612
rect 2548 66556 2558 66612
rect 0 66528 800 66556
rect 11218 66444 11228 66500
rect 11284 66444 12572 66500
rect 12628 66444 12638 66500
rect 19826 65828 19836 65884
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 20100 65828 20110 65884
rect 9426 65548 9436 65604
rect 9492 65548 10892 65604
rect 10948 65548 10958 65604
rect 22978 65436 22988 65492
rect 23044 65436 23884 65492
rect 23940 65436 23950 65492
rect 24658 65436 24668 65492
rect 24724 65436 25340 65492
rect 25396 65436 25406 65492
rect 4466 65044 4476 65100
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4740 65044 4750 65100
rect 35186 65044 35196 65100
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35460 65044 35470 65100
rect 8866 64764 8876 64820
rect 8932 64764 11340 64820
rect 11396 64764 11406 64820
rect 0 64596 800 64624
rect 0 64540 2380 64596
rect 2436 64540 2446 64596
rect 2706 64540 2716 64596
rect 2772 64540 8652 64596
rect 8708 64540 8718 64596
rect 0 64512 800 64540
rect 1810 64428 1820 64484
rect 1876 64428 3164 64484
rect 3220 64428 3230 64484
rect 10108 64372 10164 64764
rect 13346 64652 13356 64708
rect 13412 64652 14140 64708
rect 14196 64652 14206 64708
rect 24434 64428 24444 64484
rect 24500 64428 25340 64484
rect 25396 64428 25676 64484
rect 25732 64428 25742 64484
rect 10098 64316 10108 64372
rect 10164 64316 10174 64372
rect 19826 64260 19836 64316
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 20100 64260 20110 64316
rect 8978 63980 8988 64036
rect 9044 63980 10220 64036
rect 10276 63980 10286 64036
rect 25442 63980 25452 64036
rect 25508 63980 26236 64036
rect 26292 63980 26302 64036
rect 0 63924 800 63952
rect 39200 63924 40000 63952
rect 0 63868 1820 63924
rect 1876 63868 1886 63924
rect 9986 63868 9996 63924
rect 10052 63868 10892 63924
rect 10948 63868 10958 63924
rect 13906 63868 13916 63924
rect 13972 63868 14588 63924
rect 14644 63868 14654 63924
rect 24322 63868 24332 63924
rect 24388 63868 25900 63924
rect 25956 63868 26796 63924
rect 26852 63868 28476 63924
rect 28532 63868 28542 63924
rect 38210 63868 38220 63924
rect 38276 63868 40000 63924
rect 0 63840 800 63868
rect 39200 63840 40000 63868
rect 2034 63756 2044 63812
rect 2100 63756 13692 63812
rect 13748 63756 13758 63812
rect 18274 63756 18284 63812
rect 18340 63756 21420 63812
rect 21476 63756 21486 63812
rect 4466 63476 4476 63532
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4740 63476 4750 63532
rect 35186 63476 35196 63532
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35460 63476 35470 63532
rect 2146 63308 2156 63364
rect 2212 63308 14364 63364
rect 14420 63308 14430 63364
rect 18050 63308 18060 63364
rect 18116 63308 18956 63364
rect 19012 63308 19964 63364
rect 20020 63308 20030 63364
rect 0 63252 800 63280
rect 0 63196 1708 63252
rect 1764 63196 2492 63252
rect 2548 63196 2558 63252
rect 17826 63196 17836 63252
rect 17892 63196 20188 63252
rect 20244 63196 21532 63252
rect 21588 63196 21598 63252
rect 0 63168 800 63196
rect 19394 63084 19404 63140
rect 19460 63084 20188 63140
rect 21410 63084 21420 63140
rect 21476 63084 22764 63140
rect 22820 63084 22830 63140
rect 24322 63084 24332 63140
rect 24388 63084 24892 63140
rect 24948 63084 26012 63140
rect 26068 63084 26078 63140
rect 2034 62972 2044 63028
rect 2100 62972 8876 63028
rect 8932 62972 8942 63028
rect 15698 62972 15708 63028
rect 15764 62972 16492 63028
rect 16548 62972 17276 63028
rect 17332 62972 18396 63028
rect 18452 62972 18462 63028
rect 20132 62916 20188 63084
rect 23884 62972 26236 63028
rect 26292 62972 26796 63028
rect 26852 62972 26862 63028
rect 23884 62916 23940 62972
rect 17378 62860 17388 62916
rect 17444 62860 18844 62916
rect 18900 62860 18910 62916
rect 20132 62860 23884 62916
rect 23940 62860 23950 62916
rect 24658 62860 24668 62916
rect 24724 62860 25564 62916
rect 25620 62860 25630 62916
rect 12674 62748 12684 62804
rect 12740 62748 14924 62804
rect 14980 62748 16044 62804
rect 16100 62748 16110 62804
rect 19826 62692 19836 62748
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 20100 62692 20110 62748
rect 15092 62636 17836 62692
rect 17892 62636 17902 62692
rect 0 62580 800 62608
rect 15092 62580 15148 62636
rect 0 62524 1708 62580
rect 1764 62524 2492 62580
rect 2548 62524 2558 62580
rect 8082 62524 8092 62580
rect 8148 62524 8988 62580
rect 9044 62524 9054 62580
rect 11442 62524 11452 62580
rect 11508 62524 14700 62580
rect 14756 62524 15148 62580
rect 16818 62524 16828 62580
rect 16884 62524 17948 62580
rect 18004 62524 18014 62580
rect 0 62496 800 62524
rect 10210 62412 10220 62468
rect 10276 62412 11004 62468
rect 11060 62412 13244 62468
rect 13300 62412 13916 62468
rect 13972 62412 13982 62468
rect 15596 62412 18732 62468
rect 18788 62412 19516 62468
rect 19572 62412 19582 62468
rect 22082 62412 22092 62468
rect 22148 62412 23324 62468
rect 23380 62412 24556 62468
rect 24612 62412 25900 62468
rect 25956 62412 27020 62468
rect 27076 62412 27086 62468
rect 15596 62356 15652 62412
rect 14354 62300 14364 62356
rect 14420 62300 15596 62356
rect 15652 62300 15662 62356
rect 17714 62300 17724 62356
rect 17780 62300 18956 62356
rect 19012 62300 19022 62356
rect 19590 62300 19628 62356
rect 19684 62300 19694 62356
rect 24210 62300 24220 62356
rect 24276 62300 25452 62356
rect 25508 62300 29036 62356
rect 29092 62300 29102 62356
rect 8866 62188 8876 62244
rect 8932 62188 10332 62244
rect 10388 62188 10398 62244
rect 13804 62188 17612 62244
rect 17668 62188 17678 62244
rect 13804 62132 13860 62188
rect 13794 62076 13804 62132
rect 13860 62076 13870 62132
rect 19618 62076 19628 62132
rect 19684 62076 20412 62132
rect 20468 62076 20478 62132
rect 26786 62076 26796 62132
rect 26852 62076 29596 62132
rect 29652 62076 29662 62132
rect 4466 61908 4476 61964
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4740 61908 4750 61964
rect 35186 61908 35196 61964
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35460 61908 35470 61964
rect 18946 61852 18956 61908
rect 19012 61852 19292 61908
rect 19348 61852 19964 61908
rect 20020 61852 20188 61908
rect 20244 61852 20254 61908
rect 8754 61740 8764 61796
rect 8820 61740 10108 61796
rect 10164 61740 10174 61796
rect 19506 61740 19516 61796
rect 19572 61740 19740 61796
rect 19796 61740 19806 61796
rect 18162 61516 18172 61572
rect 18228 61516 20188 61572
rect 20244 61516 20254 61572
rect 10434 61404 10444 61460
rect 10500 61404 13804 61460
rect 13860 61404 13870 61460
rect 17602 61404 17612 61460
rect 17668 61404 18732 61460
rect 18788 61404 18798 61460
rect 20738 61404 20748 61460
rect 20804 61404 23324 61460
rect 23380 61404 25228 61460
rect 25284 61404 25676 61460
rect 25732 61404 25742 61460
rect 9650 61292 9660 61348
rect 9716 61292 10332 61348
rect 10388 61292 10398 61348
rect 12450 61292 12460 61348
rect 12516 61292 13580 61348
rect 13636 61292 14812 61348
rect 14868 61292 14878 61348
rect 19394 61292 19404 61348
rect 19460 61292 23212 61348
rect 23268 61292 24444 61348
rect 24500 61292 24510 61348
rect 19590 61180 19628 61236
rect 19684 61180 19694 61236
rect 19826 61124 19836 61180
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 20100 61124 20110 61180
rect 21074 60956 21084 61012
rect 21140 60956 22204 61012
rect 22260 60956 22270 61012
rect 19478 60844 19516 60900
rect 19572 60844 19582 60900
rect 18722 60732 18732 60788
rect 18788 60732 19404 60788
rect 19460 60732 19470 60788
rect 19618 60620 19628 60676
rect 19684 60620 20076 60676
rect 20132 60620 20142 60676
rect 26562 60620 26572 60676
rect 26628 60620 27804 60676
rect 27860 60620 27870 60676
rect 19954 60508 19964 60564
rect 20020 60508 21308 60564
rect 21364 60508 21374 60564
rect 6066 60396 6076 60452
rect 6132 60396 9436 60452
rect 9492 60396 11788 60452
rect 11844 60396 12236 60452
rect 12292 60396 13244 60452
rect 13300 60396 13310 60452
rect 24770 60396 24780 60452
rect 24836 60396 25340 60452
rect 25396 60396 25406 60452
rect 4466 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4750 60396
rect 35186 60340 35196 60396
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35460 60340 35470 60396
rect 18162 59948 18172 60004
rect 18228 59948 19292 60004
rect 19348 59948 19358 60004
rect 24770 59948 24780 60004
rect 24836 59948 25676 60004
rect 25732 59948 25742 60004
rect 1698 59836 1708 59892
rect 1764 59836 2492 59892
rect 2548 59836 2558 59892
rect 3332 59836 13468 59892
rect 13524 59836 13534 59892
rect 14466 59836 14476 59892
rect 14532 59836 15036 59892
rect 15092 59836 17388 59892
rect 17444 59836 17454 59892
rect 3332 59780 3388 59836
rect 2034 59724 2044 59780
rect 2100 59724 3388 59780
rect 9202 59724 9212 59780
rect 9268 59724 9772 59780
rect 9828 59724 9838 59780
rect 13346 59724 13356 59780
rect 13412 59724 13692 59780
rect 13748 59724 13758 59780
rect 19826 59556 19836 59612
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 20100 59556 20110 59612
rect 9538 59388 9548 59444
rect 9604 59388 10332 59444
rect 10388 59388 11116 59444
rect 11172 59388 11182 59444
rect 0 59220 800 59248
rect 0 59164 1708 59220
rect 1764 59164 1774 59220
rect 8194 59164 8204 59220
rect 8260 59164 9436 59220
rect 9492 59164 9502 59220
rect 16818 59164 16828 59220
rect 16884 59164 17612 59220
rect 17668 59164 18508 59220
rect 18564 59164 18574 59220
rect 0 59136 800 59164
rect 25890 59052 25900 59108
rect 25956 59052 26460 59108
rect 26516 59052 26526 59108
rect 4466 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4750 58828
rect 35186 58772 35196 58828
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35460 58772 35470 58828
rect 26338 58716 26348 58772
rect 26404 58716 27132 58772
rect 27188 58716 27198 58772
rect 11442 58604 11452 58660
rect 11508 58604 13692 58660
rect 13748 58604 13758 58660
rect 25526 58492 25564 58548
rect 25620 58492 25630 58548
rect 14242 58380 14252 58436
rect 14308 58380 17836 58436
rect 17892 58380 17902 58436
rect 25638 58380 25676 58436
rect 25732 58380 25742 58436
rect 2034 58156 2044 58212
rect 2100 58156 7756 58212
rect 7812 58156 7822 58212
rect 8642 58156 8652 58212
rect 8708 58156 9772 58212
rect 9828 58156 10108 58212
rect 10164 58156 10174 58212
rect 12898 58156 12908 58212
rect 12964 58156 13468 58212
rect 13524 58156 13534 58212
rect 17490 58156 17500 58212
rect 17556 58156 18956 58212
rect 19012 58156 19022 58212
rect 23650 58156 23660 58212
rect 23716 58156 25564 58212
rect 25620 58156 25630 58212
rect 19826 57988 19836 58044
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20100 57988 20110 58044
rect 0 57876 800 57904
rect 0 57820 1708 57876
rect 1764 57820 2492 57876
rect 2548 57820 2558 57876
rect 0 57792 800 57820
rect 2034 57708 2044 57764
rect 2100 57708 13020 57764
rect 13076 57708 13086 57764
rect 16706 57596 16716 57652
rect 16772 57596 17724 57652
rect 17780 57596 17790 57652
rect 24434 57596 24444 57652
rect 24500 57596 24510 57652
rect 24444 57540 24500 57596
rect 24444 57484 28476 57540
rect 28532 57484 28542 57540
rect 15026 57372 15036 57428
rect 15092 57372 17612 57428
rect 17668 57372 17678 57428
rect 18610 57372 18620 57428
rect 18676 57372 18844 57428
rect 18900 57372 18910 57428
rect 25106 57372 25116 57428
rect 25172 57372 26348 57428
rect 26404 57372 26414 57428
rect 0 57204 800 57232
rect 4466 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4750 57260
rect 35186 57204 35196 57260
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35460 57204 35470 57260
rect 0 57148 1708 57204
rect 1764 57148 2492 57204
rect 2548 57148 2558 57204
rect 0 57120 800 57148
rect 18386 57036 18396 57092
rect 18452 57036 21420 57092
rect 21476 57036 21486 57092
rect 26226 57036 26236 57092
rect 26292 57036 26796 57092
rect 26852 57036 28028 57092
rect 28084 57036 28094 57092
rect 16594 56924 16604 56980
rect 16660 56924 17276 56980
rect 17332 56924 18060 56980
rect 18116 56924 23212 56980
rect 23268 56924 25676 56980
rect 25732 56924 25742 56980
rect 12898 56812 12908 56868
rect 12964 56812 14028 56868
rect 14084 56812 14094 56868
rect 21522 56812 21532 56868
rect 21588 56812 21868 56868
rect 21924 56812 22652 56868
rect 22708 56812 22718 56868
rect 27570 56812 27580 56868
rect 27636 56812 28252 56868
rect 28308 56812 28318 56868
rect 14242 56700 14252 56756
rect 14308 56700 15148 56756
rect 24770 56700 24780 56756
rect 24836 56700 25676 56756
rect 25732 56700 27356 56756
rect 27412 56700 29036 56756
rect 29092 56700 29102 56756
rect 15092 56644 15148 56700
rect 12674 56588 12684 56644
rect 12740 56588 13468 56644
rect 13524 56588 13534 56644
rect 15092 56588 15484 56644
rect 15540 56588 17164 56644
rect 17220 56588 17230 56644
rect 25554 56588 25564 56644
rect 25620 56588 25676 56644
rect 25732 56588 25742 56644
rect 0 56532 800 56560
rect 0 56476 1708 56532
rect 1764 56476 2492 56532
rect 2548 56476 2558 56532
rect 23650 56476 23660 56532
rect 23716 56476 24444 56532
rect 24500 56476 25116 56532
rect 25172 56476 25788 56532
rect 25844 56476 25854 56532
rect 0 56448 800 56476
rect 19826 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20110 56476
rect 2034 56252 2044 56308
rect 2100 56252 7420 56308
rect 7476 56252 7486 56308
rect 2146 56140 2156 56196
rect 2212 56140 3388 56196
rect 8530 56140 8540 56196
rect 8596 56140 10108 56196
rect 10164 56140 10174 56196
rect 18722 56140 18732 56196
rect 18788 56140 24556 56196
rect 24612 56140 26908 56196
rect 26964 56140 29372 56196
rect 29428 56140 29932 56196
rect 29988 56140 29998 56196
rect 0 55860 800 55888
rect 3332 55860 3388 56140
rect 8194 56028 8204 56084
rect 8260 56028 9436 56084
rect 9492 56028 9502 56084
rect 9986 56028 9996 56084
rect 10052 56028 17500 56084
rect 17556 56028 17566 56084
rect 21746 56028 21756 56084
rect 21812 56028 22764 56084
rect 22820 56028 22830 56084
rect 25890 56028 25900 56084
rect 25956 56028 27580 56084
rect 27636 56028 27646 56084
rect 6626 55916 6636 55972
rect 6692 55916 9660 55972
rect 9716 55916 9726 55972
rect 0 55804 1708 55860
rect 1764 55804 2492 55860
rect 2548 55804 2558 55860
rect 3332 55804 7588 55860
rect 9090 55804 9100 55860
rect 9156 55804 9772 55860
rect 9828 55804 9838 55860
rect 16594 55804 16604 55860
rect 16660 55804 17836 55860
rect 17892 55804 18396 55860
rect 18452 55804 18462 55860
rect 25778 55804 25788 55860
rect 25844 55804 27356 55860
rect 27412 55804 27422 55860
rect 0 55776 800 55804
rect 7532 55748 7588 55804
rect 7532 55692 7644 55748
rect 7700 55692 7710 55748
rect 4466 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4750 55692
rect 35186 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35470 55692
rect 6290 55468 6300 55524
rect 6356 55468 12012 55524
rect 12068 55468 12078 55524
rect 8306 55356 8316 55412
rect 8372 55356 9324 55412
rect 9380 55356 9390 55412
rect 11554 55356 11564 55412
rect 11620 55356 12236 55412
rect 12292 55356 12302 55412
rect 17714 55356 17724 55412
rect 17780 55356 21980 55412
rect 22036 55356 22046 55412
rect 28354 55356 28364 55412
rect 28420 55356 29260 55412
rect 29316 55356 29326 55412
rect 2034 55244 2044 55300
rect 2100 55244 8652 55300
rect 8708 55244 8718 55300
rect 9202 55244 9212 55300
rect 9268 55244 9660 55300
rect 9716 55244 9726 55300
rect 17378 55244 17388 55300
rect 17444 55244 19068 55300
rect 19124 55244 19134 55300
rect 22082 55244 22092 55300
rect 22148 55244 24444 55300
rect 24500 55244 29596 55300
rect 29652 55244 29662 55300
rect 0 55188 800 55216
rect 0 55132 1708 55188
rect 1764 55132 2492 55188
rect 2548 55132 2558 55188
rect 6962 55132 6972 55188
rect 7028 55132 8092 55188
rect 8148 55132 8158 55188
rect 17154 55132 17164 55188
rect 17220 55132 19292 55188
rect 19348 55132 19358 55188
rect 0 55104 800 55132
rect 10546 55020 10556 55076
rect 10612 55020 11004 55076
rect 11060 55020 11900 55076
rect 11956 55020 11966 55076
rect 19826 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20110 54908
rect 12450 54796 12460 54852
rect 12516 54796 13692 54852
rect 13748 54796 13758 54852
rect 8866 54684 8876 54740
rect 8932 54684 9772 54740
rect 9828 54684 9838 54740
rect 14914 54572 14924 54628
rect 14980 54572 15484 54628
rect 15540 54572 17724 54628
rect 17780 54572 18844 54628
rect 18900 54572 18910 54628
rect 8642 54460 8652 54516
rect 8708 54460 9100 54516
rect 9156 54460 9166 54516
rect 18274 54460 18284 54516
rect 18340 54460 18956 54516
rect 19012 54460 20076 54516
rect 20132 54460 20142 54516
rect 4466 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4750 54124
rect 35186 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35470 54124
rect 7858 53676 7868 53732
rect 7924 53676 9548 53732
rect 9604 53676 9614 53732
rect 18162 53676 18172 53732
rect 18228 53676 19180 53732
rect 19236 53676 19246 53732
rect 19730 53676 19740 53732
rect 19796 53676 21420 53732
rect 21476 53676 21486 53732
rect 21746 53676 21756 53732
rect 21812 53676 23884 53732
rect 23940 53676 23950 53732
rect 25890 53676 25900 53732
rect 25956 53676 27132 53732
rect 27188 53676 28476 53732
rect 28532 53676 28542 53732
rect 8754 53564 8764 53620
rect 8820 53564 16380 53620
rect 16436 53564 16446 53620
rect 16930 53564 16940 53620
rect 16996 53564 19292 53620
rect 19348 53564 19358 53620
rect 23090 53564 23100 53620
rect 23156 53564 25340 53620
rect 25396 53564 25406 53620
rect 16940 53508 16996 53564
rect 16482 53452 16492 53508
rect 16548 53452 16996 53508
rect 18162 53452 18172 53508
rect 18228 53452 18396 53508
rect 18452 53452 19516 53508
rect 19572 53452 19582 53508
rect 20738 53452 20748 53508
rect 20804 53452 22092 53508
rect 22148 53452 24444 53508
rect 24500 53452 24510 53508
rect 26898 53452 26908 53508
rect 26964 53452 27356 53508
rect 27412 53452 27422 53508
rect 19826 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20110 53340
rect 15250 53228 15260 53284
rect 15316 53228 18956 53284
rect 19012 53228 19022 53284
rect 0 53172 800 53200
rect 39200 53172 40000 53200
rect 0 53116 1708 53172
rect 1764 53116 2492 53172
rect 2548 53116 2558 53172
rect 16034 53116 16044 53172
rect 16100 53116 18732 53172
rect 18788 53116 18798 53172
rect 37986 53116 37996 53172
rect 38052 53116 40000 53172
rect 0 53088 800 53116
rect 39200 53088 40000 53116
rect 15138 53004 15148 53060
rect 15204 53004 16604 53060
rect 16660 53004 16670 53060
rect 21522 53004 21532 53060
rect 21588 53004 23772 53060
rect 23828 53004 24108 53060
rect 24164 53004 26796 53060
rect 26852 53004 26862 53060
rect 15026 52892 15036 52948
rect 15092 52836 15148 52948
rect 16370 52892 16380 52948
rect 16436 52892 17388 52948
rect 17444 52892 17454 52948
rect 20962 52892 20972 52948
rect 21028 52892 21980 52948
rect 22036 52892 24220 52948
rect 24276 52892 24286 52948
rect 28466 52892 28476 52948
rect 28532 52892 33068 52948
rect 33124 52892 33134 52948
rect 15092 52780 16268 52836
rect 16324 52780 18172 52836
rect 18228 52780 18238 52836
rect 22166 52780 22204 52836
rect 22260 52780 22270 52836
rect 27346 52780 27356 52836
rect 27412 52780 28700 52836
rect 28756 52780 28766 52836
rect 15586 52668 15596 52724
rect 15652 52668 20076 52724
rect 20132 52668 20142 52724
rect 4466 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4750 52556
rect 35186 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35470 52556
rect 2034 52108 2044 52164
rect 2100 52108 11452 52164
rect 11508 52108 11518 52164
rect 11778 52108 11788 52164
rect 11844 52108 12124 52164
rect 12180 52108 12190 52164
rect 16706 52108 16716 52164
rect 16772 52108 20748 52164
rect 20804 52108 20814 52164
rect 21830 52108 21868 52164
rect 21924 52108 21934 52164
rect 32946 52108 32956 52164
rect 33012 52108 33740 52164
rect 33796 52108 33806 52164
rect 2146 51996 2156 52052
rect 2212 51996 8540 52052
rect 8596 51996 8606 52052
rect 12898 51996 12908 52052
rect 12964 51996 15596 52052
rect 15652 51996 18620 52052
rect 18676 51996 18686 52052
rect 22306 51996 22316 52052
rect 22372 51996 24444 52052
rect 24500 51996 24510 52052
rect 9762 51884 9772 51940
rect 9828 51884 10220 51940
rect 10276 51884 10286 51940
rect 11666 51884 11676 51940
rect 11732 51884 12236 51940
rect 12292 51884 12302 51940
rect 12460 51884 16492 51940
rect 16548 51884 16558 51940
rect 16706 51884 16716 51940
rect 16772 51884 17948 51940
rect 18004 51884 18508 51940
rect 18564 51884 18574 51940
rect 0 51828 800 51856
rect 12460 51828 12516 51884
rect 0 51772 1708 51828
rect 1764 51772 2492 51828
rect 2548 51772 2558 51828
rect 8978 51772 8988 51828
rect 9044 51772 9436 51828
rect 9492 51772 12516 51828
rect 15092 51772 17836 51828
rect 17892 51772 17902 51828
rect 20738 51772 20748 51828
rect 20804 51772 22092 51828
rect 22148 51772 25228 51828
rect 25284 51772 25294 51828
rect 0 51744 800 51772
rect 15092 51716 15148 51772
rect 19826 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20110 51772
rect 9986 51660 9996 51716
rect 10052 51660 15148 51716
rect 2034 51436 2044 51492
rect 2100 51436 11452 51492
rect 11508 51436 11518 51492
rect 14802 51436 14812 51492
rect 14868 51436 16604 51492
rect 16660 51436 16670 51492
rect 21074 51436 21084 51492
rect 21140 51436 23100 51492
rect 23156 51436 23166 51492
rect 25666 51436 25676 51492
rect 25732 51436 26908 51492
rect 26964 51436 26974 51492
rect 8530 51324 8540 51380
rect 8596 51324 9772 51380
rect 9828 51324 9838 51380
rect 22418 51324 22428 51380
rect 22484 51324 24668 51380
rect 24724 51324 24734 51380
rect 14578 51212 14588 51268
rect 14644 51212 15708 51268
rect 15764 51212 15774 51268
rect 0 51156 800 51184
rect 0 51100 1708 51156
rect 1764 51100 2492 51156
rect 2548 51100 2558 51156
rect 21746 51100 21756 51156
rect 21812 51100 22428 51156
rect 22484 51100 22494 51156
rect 0 51072 800 51100
rect 4466 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4750 50988
rect 35186 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35470 50988
rect 19730 50764 19740 50820
rect 19796 50764 21084 50820
rect 21140 50764 21150 50820
rect 2706 50540 2716 50596
rect 2772 50540 9660 50596
rect 9716 50540 9726 50596
rect 11666 50540 11676 50596
rect 11732 50540 12124 50596
rect 12180 50540 12190 50596
rect 16258 50540 16268 50596
rect 16324 50540 17724 50596
rect 17780 50540 17790 50596
rect 0 50484 800 50512
rect 0 50428 1708 50484
rect 1764 50428 2492 50484
rect 2548 50428 2558 50484
rect 7746 50428 7756 50484
rect 7812 50428 9548 50484
rect 9604 50428 9614 50484
rect 9762 50428 9772 50484
rect 9828 50428 10668 50484
rect 10724 50428 11452 50484
rect 11508 50428 12684 50484
rect 12740 50428 12750 50484
rect 12898 50428 12908 50484
rect 12964 50428 15148 50484
rect 15204 50428 15214 50484
rect 15698 50428 15708 50484
rect 15764 50428 16380 50484
rect 16436 50428 16446 50484
rect 18498 50428 18508 50484
rect 18564 50428 18956 50484
rect 19012 50428 19022 50484
rect 20626 50428 20636 50484
rect 20692 50428 25228 50484
rect 25284 50428 25294 50484
rect 0 50400 800 50428
rect 2034 50316 2044 50372
rect 2100 50316 11228 50372
rect 11284 50316 11294 50372
rect 8754 50204 8764 50260
rect 8820 50204 10332 50260
rect 10388 50204 10398 50260
rect 14802 50204 14812 50260
rect 14868 50204 15260 50260
rect 15316 50204 15326 50260
rect 19826 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20110 50204
rect 8372 49980 15708 50036
rect 15764 49980 17836 50036
rect 17892 49980 18396 50036
rect 18452 49980 18462 50036
rect 2034 49868 2044 49924
rect 2100 49868 7196 49924
rect 7252 49868 7262 49924
rect 0 49812 800 49840
rect 8372 49812 8428 49980
rect 22642 49868 22652 49924
rect 22708 49868 24556 49924
rect 24612 49868 24622 49924
rect 39200 49812 40000 49840
rect 0 49756 2380 49812
rect 2436 49756 3164 49812
rect 3220 49756 3230 49812
rect 8194 49756 8204 49812
rect 8260 49756 8428 49812
rect 9090 49756 9100 49812
rect 9156 49756 10220 49812
rect 10276 49756 10286 49812
rect 21634 49756 21644 49812
rect 21700 49756 22764 49812
rect 22820 49756 22830 49812
rect 36754 49756 36764 49812
rect 36820 49756 40000 49812
rect 0 49728 800 49756
rect 9772 49700 9828 49756
rect 39200 49728 40000 49756
rect 1698 49644 1708 49700
rect 1764 49644 2940 49700
rect 2996 49644 3006 49700
rect 9762 49644 9772 49700
rect 9828 49644 9838 49700
rect 30482 49644 30492 49700
rect 30548 49644 32396 49700
rect 32452 49644 32462 49700
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 14802 49308 14812 49364
rect 14868 49308 18172 49364
rect 18228 49308 18238 49364
rect 0 49140 800 49168
rect 0 49084 1708 49140
rect 1764 49084 1774 49140
rect 29138 49084 29148 49140
rect 29204 49084 30268 49140
rect 30324 49084 30334 49140
rect 32386 49084 32396 49140
rect 32452 49084 33292 49140
rect 33348 49084 33358 49140
rect 0 49056 800 49084
rect 18050 48972 18060 49028
rect 18116 48972 20412 49028
rect 20468 48972 26460 49028
rect 26516 48972 26526 49028
rect 27010 48972 27020 49028
rect 27076 48972 27916 49028
rect 27972 48972 31164 49028
rect 31220 48972 31948 49028
rect 32004 48972 34860 49028
rect 34916 48972 34926 49028
rect 35074 48972 35084 49028
rect 35140 48972 35420 49028
rect 35476 48972 35486 49028
rect 2034 48860 2044 48916
rect 2100 48860 6636 48916
rect 6692 48860 6702 48916
rect 20850 48860 20860 48916
rect 20916 48860 21420 48916
rect 21476 48860 22876 48916
rect 22932 48860 22942 48916
rect 32050 48860 32060 48916
rect 32116 48860 34412 48916
rect 34468 48860 35980 48916
rect 36036 48860 36046 48916
rect 7074 48748 7084 48804
rect 7140 48748 8428 48804
rect 8484 48748 8494 48804
rect 21186 48748 21196 48804
rect 21252 48748 21756 48804
rect 21812 48748 23660 48804
rect 23716 48748 24220 48804
rect 24276 48748 24286 48804
rect 33730 48748 33740 48804
rect 33796 48748 34524 48804
rect 34580 48748 34860 48804
rect 34916 48748 35644 48804
rect 35700 48748 35710 48804
rect 34850 48636 34860 48692
rect 34916 48636 35084 48692
rect 35140 48636 35150 48692
rect 19826 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20110 48636
rect 0 48468 800 48496
rect 0 48412 1708 48468
rect 1764 48412 2492 48468
rect 2548 48412 2558 48468
rect 5954 48412 5964 48468
rect 6020 48412 6636 48468
rect 6692 48412 6702 48468
rect 10546 48412 10556 48468
rect 10612 48412 15148 48468
rect 18386 48412 18396 48468
rect 18452 48412 19068 48468
rect 19124 48412 19134 48468
rect 20290 48412 20300 48468
rect 20356 48412 22764 48468
rect 22820 48412 22830 48468
rect 23986 48412 23996 48468
rect 24052 48412 25004 48468
rect 25060 48412 26124 48468
rect 26180 48412 26190 48468
rect 32498 48412 32508 48468
rect 32564 48412 35868 48468
rect 35924 48412 35934 48468
rect 0 48384 800 48412
rect 15092 48356 15148 48412
rect 2034 48300 2044 48356
rect 2100 48300 7980 48356
rect 8036 48300 8046 48356
rect 15092 48300 26796 48356
rect 26852 48300 27244 48356
rect 27300 48300 27468 48356
rect 27524 48300 27534 48356
rect 31266 48300 31276 48356
rect 31332 48300 32396 48356
rect 32452 48300 33516 48356
rect 33572 48300 33582 48356
rect 11890 48188 11900 48244
rect 11956 48188 15484 48244
rect 15540 48188 15550 48244
rect 16258 48188 16268 48244
rect 16324 48188 17500 48244
rect 17556 48188 18732 48244
rect 18788 48188 18798 48244
rect 21522 48188 21532 48244
rect 21588 48188 22316 48244
rect 22372 48188 22382 48244
rect 24658 48188 24668 48244
rect 24724 48188 25340 48244
rect 25396 48188 25406 48244
rect 26450 48188 26460 48244
rect 26516 48188 27132 48244
rect 27188 48188 27198 48244
rect 31826 48188 31836 48244
rect 31892 48188 32620 48244
rect 32676 48188 32686 48244
rect 18498 48076 18508 48132
rect 18564 48076 19180 48132
rect 19236 48076 19246 48132
rect 28018 48076 28028 48132
rect 28084 48076 29932 48132
rect 29988 48076 29998 48132
rect 16594 47964 16604 48020
rect 16660 47964 20524 48020
rect 20580 47964 23100 48020
rect 23156 47964 23166 48020
rect 31826 47852 31836 47908
rect 31892 47852 33180 47908
rect 33236 47852 34076 47908
rect 34132 47852 34142 47908
rect 0 47796 800 47824
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 0 47740 1708 47796
rect 1764 47740 2492 47796
rect 2548 47740 2558 47796
rect 32946 47740 32956 47796
rect 33012 47740 34300 47796
rect 34356 47740 34366 47796
rect 0 47712 800 47740
rect 20738 47628 20748 47684
rect 20804 47628 22764 47684
rect 22820 47628 22830 47684
rect 24098 47516 24108 47572
rect 24164 47516 24556 47572
rect 24612 47516 25340 47572
rect 25396 47516 25406 47572
rect 33180 47460 33236 47740
rect 34738 47628 34748 47684
rect 34804 47628 36092 47684
rect 36148 47628 36158 47684
rect 33170 47404 33180 47460
rect 33236 47404 33246 47460
rect 8866 47292 8876 47348
rect 8932 47292 10220 47348
rect 10276 47292 11340 47348
rect 11396 47292 11406 47348
rect 15474 47292 15484 47348
rect 15540 47292 17948 47348
rect 18004 47292 18014 47348
rect 19506 47292 19516 47348
rect 19572 47292 20412 47348
rect 20468 47292 20478 47348
rect 18162 47180 18172 47236
rect 18228 47180 20300 47236
rect 20356 47180 20366 47236
rect 27122 47180 27132 47236
rect 27188 47180 31500 47236
rect 31556 47180 31566 47236
rect 39200 47124 40000 47152
rect 21858 47068 21868 47124
rect 21924 47068 21934 47124
rect 28354 47068 28364 47124
rect 28420 47068 29260 47124
rect 29316 47068 29326 47124
rect 36866 47068 36876 47124
rect 36932 47068 40000 47124
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 21868 47012 21924 47068
rect 39200 47040 40000 47068
rect 8866 46956 8876 47012
rect 8932 46956 9660 47012
rect 9716 46956 9726 47012
rect 21868 46956 22204 47012
rect 22260 46956 23996 47012
rect 24052 46956 24062 47012
rect 10770 46844 10780 46900
rect 10836 46844 11340 46900
rect 11396 46844 11406 46900
rect 8754 46732 8764 46788
rect 8820 46732 9436 46788
rect 9492 46732 9502 46788
rect 31714 46732 31724 46788
rect 31780 46732 31948 46788
rect 32004 46732 32956 46788
rect 33012 46732 33022 46788
rect 8978 46620 8988 46676
rect 9044 46620 10780 46676
rect 10836 46620 10846 46676
rect 19142 46620 19180 46676
rect 19236 46620 19246 46676
rect 22054 46620 22092 46676
rect 22148 46620 22158 46676
rect 30146 46620 30156 46676
rect 30212 46620 31612 46676
rect 31668 46620 31678 46676
rect 32498 46620 32508 46676
rect 32564 46620 33740 46676
rect 33796 46620 33806 46676
rect 7298 46508 7308 46564
rect 7364 46508 8540 46564
rect 8596 46508 8606 46564
rect 26114 46508 26124 46564
rect 26180 46508 27356 46564
rect 27412 46508 27422 46564
rect 39200 46452 40000 46480
rect 22418 46396 22428 46452
rect 22484 46396 25676 46452
rect 25732 46396 25742 46452
rect 32386 46396 32396 46452
rect 32452 46396 33292 46452
rect 33348 46396 33358 46452
rect 34738 46396 34748 46452
rect 34804 46396 40000 46452
rect 39200 46368 40000 46396
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 21634 46060 21644 46116
rect 21700 46060 22428 46116
rect 22484 46060 22494 46116
rect 28578 46060 28588 46116
rect 28644 46060 29932 46116
rect 29988 46060 32284 46116
rect 32340 46060 32350 46116
rect 14914 45948 14924 46004
rect 14980 45948 16940 46004
rect 16996 45948 17500 46004
rect 17556 45948 17566 46004
rect 14242 45836 14252 45892
rect 14308 45836 15036 45892
rect 15092 45836 15372 45892
rect 15428 45836 15438 45892
rect 21634 45836 21644 45892
rect 21700 45836 21980 45892
rect 22036 45836 22046 45892
rect 9650 45724 9660 45780
rect 9716 45724 10780 45780
rect 10836 45724 10846 45780
rect 22082 45724 22092 45780
rect 22148 45724 24108 45780
rect 24164 45724 24174 45780
rect 12898 45612 12908 45668
rect 12964 45612 13916 45668
rect 13972 45612 14588 45668
rect 14644 45612 14654 45668
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 9202 45276 9212 45332
rect 9268 45276 9884 45332
rect 9940 45276 9950 45332
rect 14802 45276 14812 45332
rect 14868 45276 15148 45332
rect 17938 45276 17948 45332
rect 18004 45276 18620 45332
rect 18676 45276 18686 45332
rect 19954 45276 19964 45332
rect 20020 45276 21868 45332
rect 21924 45276 21934 45332
rect 25554 45276 25564 45332
rect 25620 45276 26012 45332
rect 26068 45276 27580 45332
rect 27636 45276 27646 45332
rect 33282 45276 33292 45332
rect 33348 45276 34412 45332
rect 34468 45276 34478 45332
rect 15092 45220 15148 45276
rect 2034 45164 2044 45220
rect 2100 45164 6636 45220
rect 6692 45164 6702 45220
rect 8754 45164 8764 45220
rect 8820 45164 10220 45220
rect 10276 45164 10286 45220
rect 15092 45164 15484 45220
rect 15540 45164 18396 45220
rect 18452 45164 18462 45220
rect 22082 45164 22092 45220
rect 22148 45164 22988 45220
rect 23044 45164 23054 45220
rect 30818 45164 30828 45220
rect 30884 45164 31612 45220
rect 31668 45164 33180 45220
rect 33236 45164 34076 45220
rect 34132 45164 34142 45220
rect 10882 45052 10892 45108
rect 10948 45052 12572 45108
rect 12628 45052 14476 45108
rect 14532 45052 16604 45108
rect 16660 45052 16670 45108
rect 17714 45052 17724 45108
rect 17780 45052 18060 45108
rect 18116 45052 18844 45108
rect 18900 45052 18910 45108
rect 19618 45052 19628 45108
rect 19684 45052 19852 45108
rect 19908 45052 19918 45108
rect 32386 45052 32396 45108
rect 32452 45052 33292 45108
rect 33348 45052 34300 45108
rect 34356 45052 34366 45108
rect 1698 44940 1708 44996
rect 1764 44940 2492 44996
rect 2548 44940 2558 44996
rect 31938 44940 31948 44996
rect 32004 44940 33180 44996
rect 33236 44940 34972 44996
rect 35028 44940 35038 44996
rect 36418 44940 36428 44996
rect 36484 44940 38220 44996
rect 38276 44940 38286 44996
rect 5954 44828 5964 44884
rect 6020 44828 6860 44884
rect 6916 44828 6926 44884
rect 20178 44828 20188 44884
rect 20244 44828 20860 44884
rect 20916 44828 20926 44884
rect 34738 44828 34748 44884
rect 34804 44828 36092 44884
rect 36148 44828 36158 44884
rect 6962 44716 6972 44772
rect 7028 44716 8092 44772
rect 8148 44716 8158 44772
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 17042 44492 17052 44548
rect 17108 44492 18508 44548
rect 18564 44492 18574 44548
rect 20738 44492 20748 44548
rect 20804 44492 21420 44548
rect 21476 44492 21486 44548
rect 0 44436 800 44464
rect 0 44380 1708 44436
rect 1764 44380 1774 44436
rect 0 44352 800 44380
rect 12898 44268 12908 44324
rect 12964 44268 13580 44324
rect 13636 44268 13646 44324
rect 14018 44268 14028 44324
rect 14084 44268 15708 44324
rect 15764 44268 15774 44324
rect 18386 44268 18396 44324
rect 18452 44268 21756 44324
rect 21812 44268 21822 44324
rect 9426 44156 9436 44212
rect 9492 44156 13916 44212
rect 13972 44156 16156 44212
rect 16212 44156 16222 44212
rect 18610 44156 18620 44212
rect 18676 44156 19180 44212
rect 19236 44156 19246 44212
rect 23426 44156 23436 44212
rect 23492 44156 24780 44212
rect 24836 44156 24846 44212
rect 2034 44044 2044 44100
rect 2100 44044 7644 44100
rect 7700 44044 7710 44100
rect 15362 44044 15372 44100
rect 15428 44044 17276 44100
rect 17332 44044 17342 44100
rect 17714 44044 17724 44100
rect 17780 44044 18284 44100
rect 18340 44044 18350 44100
rect 18722 44044 18732 44100
rect 18788 44044 19404 44100
rect 19460 44044 19470 44100
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 0 43764 800 43792
rect 0 43708 1708 43764
rect 1764 43708 2492 43764
rect 2548 43708 2558 43764
rect 8194 43708 8204 43764
rect 8260 43708 14028 43764
rect 14084 43708 14094 43764
rect 15698 43708 15708 43764
rect 15764 43708 19852 43764
rect 19908 43708 19918 43764
rect 24322 43708 24332 43764
rect 24388 43708 29596 43764
rect 29652 43708 29662 43764
rect 0 43680 800 43708
rect 20290 43596 20300 43652
rect 20356 43596 21420 43652
rect 21476 43596 21486 43652
rect 21858 43596 21868 43652
rect 21924 43596 22204 43652
rect 22260 43596 22270 43652
rect 24882 43596 24892 43652
rect 24948 43596 26908 43652
rect 27458 43596 27468 43652
rect 27524 43596 28028 43652
rect 28084 43596 28094 43652
rect 26852 43540 26908 43596
rect 5282 43484 5292 43540
rect 5348 43484 6524 43540
rect 6580 43484 6590 43540
rect 16146 43484 16156 43540
rect 16212 43484 18284 43540
rect 18340 43484 18350 43540
rect 22194 43484 22204 43540
rect 22260 43484 22876 43540
rect 22932 43484 22942 43540
rect 26852 43484 28700 43540
rect 28756 43484 28766 43540
rect 30034 43484 30044 43540
rect 30100 43484 31388 43540
rect 31444 43484 31454 43540
rect 33282 43484 33292 43540
rect 33348 43484 33964 43540
rect 34020 43484 34030 43540
rect 14130 43372 14140 43428
rect 14196 43372 15596 43428
rect 15652 43372 15932 43428
rect 15988 43372 18620 43428
rect 18676 43372 18686 43428
rect 18946 43260 18956 43316
rect 19012 43260 19628 43316
rect 19684 43260 19694 43316
rect 23538 43148 23548 43204
rect 23604 43148 25564 43204
rect 25620 43148 26796 43204
rect 26852 43148 26862 43204
rect 31948 43148 32060 43204
rect 32116 43148 32126 43204
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 22418 43036 22428 43092
rect 22484 43036 22988 43092
rect 23044 43036 23054 43092
rect 26114 42924 26124 42980
rect 26180 42924 26796 42980
rect 26852 42924 27580 42980
rect 27636 42924 27646 42980
rect 28690 42924 28700 42980
rect 28756 42924 29596 42980
rect 29652 42924 29662 42980
rect 9874 42812 9884 42868
rect 9940 42812 10556 42868
rect 10612 42812 21644 42868
rect 21700 42812 21710 42868
rect 22978 42812 22988 42868
rect 23044 42812 23660 42868
rect 23716 42812 23726 42868
rect 28130 42812 28140 42868
rect 28196 42812 30268 42868
rect 30324 42812 31724 42868
rect 31780 42812 31790 42868
rect 31948 42756 32004 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 6514 42700 6524 42756
rect 6580 42700 7084 42756
rect 7140 42700 10108 42756
rect 10164 42700 10174 42756
rect 29250 42700 29260 42756
rect 29316 42700 30604 42756
rect 30660 42700 30670 42756
rect 31938 42700 31948 42756
rect 32004 42700 32014 42756
rect 33170 42700 33180 42756
rect 33236 42700 33404 42756
rect 33460 42700 34748 42756
rect 34804 42700 34814 42756
rect 14690 42588 14700 42644
rect 14756 42588 16380 42644
rect 16436 42588 16446 42644
rect 28354 42588 28364 42644
rect 28420 42588 29484 42644
rect 29540 42588 29550 42644
rect 31266 42588 31276 42644
rect 31332 42588 31612 42644
rect 31668 42588 31678 42644
rect 32162 42588 32172 42644
rect 32228 42588 32956 42644
rect 33012 42588 33022 42644
rect 8306 42476 8316 42532
rect 8372 42476 10556 42532
rect 10612 42476 10622 42532
rect 29586 42476 29596 42532
rect 29652 42476 30940 42532
rect 30996 42476 31006 42532
rect 33170 42476 33180 42532
rect 33236 42476 34076 42532
rect 34132 42476 34142 42532
rect 35410 42476 35420 42532
rect 35476 42476 35486 42532
rect 35420 42420 35476 42476
rect 39200 42420 40000 42448
rect 29362 42364 29372 42420
rect 29428 42364 31276 42420
rect 31332 42364 31342 42420
rect 32834 42364 32844 42420
rect 32900 42364 33292 42420
rect 33348 42364 33358 42420
rect 35420 42364 40000 42420
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 39200 42336 40000 42364
rect 28914 42252 28924 42308
rect 28980 42252 29820 42308
rect 29876 42252 29886 42308
rect 30034 42252 30044 42308
rect 30100 42252 32284 42308
rect 32340 42252 32620 42308
rect 32676 42252 32686 42308
rect 36306 42252 36316 42308
rect 36372 42252 38220 42308
rect 38276 42252 38286 42308
rect 14242 42140 14252 42196
rect 14308 42140 16604 42196
rect 16660 42140 16670 42196
rect 18162 42140 18172 42196
rect 18228 42140 19852 42196
rect 19908 42140 19918 42196
rect 28242 42140 28252 42196
rect 28308 42140 29932 42196
rect 29988 42140 29998 42196
rect 31266 42140 31276 42196
rect 31332 42140 31836 42196
rect 31892 42140 32732 42196
rect 32788 42140 32798 42196
rect 34626 42140 34636 42196
rect 34692 42140 36092 42196
rect 36148 42140 36158 42196
rect 22866 42028 22876 42084
rect 22932 42028 23548 42084
rect 23604 42028 23614 42084
rect 28466 42028 28476 42084
rect 28532 42028 29148 42084
rect 29204 42028 29708 42084
rect 29764 42028 29774 42084
rect 18722 41916 18732 41972
rect 18788 41916 20636 41972
rect 20692 41916 20702 41972
rect 22082 41916 22092 41972
rect 22148 41916 30828 41972
rect 30884 41916 30894 41972
rect 33506 41916 33516 41972
rect 33572 41916 33964 41972
rect 34020 41916 34636 41972
rect 34692 41916 34702 41972
rect 16706 41804 16716 41860
rect 16772 41804 19964 41860
rect 20020 41804 20030 41860
rect 21746 41804 21756 41860
rect 21812 41804 25676 41860
rect 25732 41804 26236 41860
rect 26292 41804 26302 41860
rect 30370 41804 30380 41860
rect 30436 41804 32956 41860
rect 33012 41804 33022 41860
rect 33730 41804 33740 41860
rect 33796 41804 36092 41860
rect 36148 41804 36158 41860
rect 36418 41804 36428 41860
rect 36484 41804 38220 41860
rect 38276 41804 38286 41860
rect 39200 41748 40000 41776
rect 16594 41692 16604 41748
rect 16660 41692 17500 41748
rect 17556 41692 18732 41748
rect 18788 41692 18844 41748
rect 18900 41692 18910 41748
rect 19170 41692 19180 41748
rect 19236 41692 20636 41748
rect 20692 41692 22092 41748
rect 22148 41692 22158 41748
rect 22530 41692 22540 41748
rect 22596 41692 22988 41748
rect 23044 41692 23054 41748
rect 24098 41692 24108 41748
rect 24164 41692 25452 41748
rect 25508 41692 25518 41748
rect 26338 41692 26348 41748
rect 26404 41692 29372 41748
rect 29428 41692 29438 41748
rect 32386 41692 32396 41748
rect 32452 41692 33180 41748
rect 33236 41692 33628 41748
rect 33684 41692 33694 41748
rect 34962 41692 34972 41748
rect 35028 41692 40000 41748
rect 39200 41664 40000 41692
rect 30034 41580 30044 41636
rect 30100 41580 31052 41636
rect 31108 41580 31118 41636
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 22726 41468 22764 41524
rect 22820 41468 22830 41524
rect 28354 41468 28364 41524
rect 28420 41468 29484 41524
rect 29540 41468 31836 41524
rect 31892 41468 31902 41524
rect 21634 41356 21644 41412
rect 21700 41356 22428 41412
rect 22484 41356 22494 41412
rect 30706 41356 30716 41412
rect 30772 41356 31724 41412
rect 31780 41356 31790 41412
rect 9202 41244 9212 41300
rect 9268 41244 10444 41300
rect 10500 41244 10510 41300
rect 27794 41244 27804 41300
rect 27860 41244 31388 41300
rect 31444 41244 31454 41300
rect 11218 41132 11228 41188
rect 11284 41132 11900 41188
rect 11956 41132 11966 41188
rect 1810 41020 1820 41076
rect 1876 41020 2492 41076
rect 2548 41020 2558 41076
rect 10098 41020 10108 41076
rect 10164 41020 14140 41076
rect 14196 41020 14206 41076
rect 19282 41020 19292 41076
rect 19348 41020 21756 41076
rect 21812 41020 21822 41076
rect 24742 41020 24780 41076
rect 24836 41020 25228 41076
rect 25284 41020 25294 41076
rect 25890 41020 25900 41076
rect 25956 41020 26796 41076
rect 26852 41020 26862 41076
rect 27794 41020 27804 41076
rect 27860 41020 28364 41076
rect 28420 41020 30044 41076
rect 30100 41020 30110 41076
rect 30706 41020 30716 41076
rect 30772 41020 31948 41076
rect 32004 41020 32014 41076
rect 2034 40908 2044 40964
rect 2100 40908 9660 40964
rect 9716 40908 9726 40964
rect 19170 40908 19180 40964
rect 19236 40908 19516 40964
rect 19572 40908 19582 40964
rect 21858 40908 21868 40964
rect 21924 40908 23436 40964
rect 23492 40908 23502 40964
rect 25778 40908 25788 40964
rect 25844 40908 26236 40964
rect 26292 40908 26302 40964
rect 31042 40908 31052 40964
rect 31108 40908 31500 40964
rect 31556 40908 31566 40964
rect 32050 40908 32060 40964
rect 32116 40908 32956 40964
rect 33012 40908 34188 40964
rect 34244 40908 34254 40964
rect 31378 40796 31388 40852
rect 31444 40796 31836 40852
rect 31892 40796 32508 40852
rect 32564 40796 32574 40852
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 19058 40684 19068 40740
rect 19124 40684 19628 40740
rect 19684 40684 19694 40740
rect 29250 40684 29260 40740
rect 29316 40684 32396 40740
rect 32452 40684 32462 40740
rect 9762 40572 9772 40628
rect 9828 40572 10332 40628
rect 10388 40572 10398 40628
rect 20178 40572 20188 40628
rect 20244 40572 21868 40628
rect 21924 40572 21934 40628
rect 22418 40572 22428 40628
rect 22484 40572 25900 40628
rect 25956 40572 25966 40628
rect 28466 40572 28476 40628
rect 28532 40572 30492 40628
rect 30548 40572 30940 40628
rect 30996 40572 31006 40628
rect 11554 40460 11564 40516
rect 11620 40460 12908 40516
rect 12964 40460 13468 40516
rect 13524 40460 13534 40516
rect 17154 40460 17164 40516
rect 17220 40460 23324 40516
rect 23380 40460 23996 40516
rect 24052 40460 24062 40516
rect 0 40404 800 40432
rect 0 40348 1820 40404
rect 1876 40348 1886 40404
rect 21522 40348 21532 40404
rect 21588 40348 23100 40404
rect 23156 40348 23166 40404
rect 30594 40348 30604 40404
rect 30660 40348 32060 40404
rect 32116 40348 35980 40404
rect 36036 40348 36046 40404
rect 0 40320 800 40348
rect 1698 40236 1708 40292
rect 1764 40236 2492 40292
rect 2548 40236 2558 40292
rect 18582 40236 18620 40292
rect 18676 40236 18686 40292
rect 20962 40236 20972 40292
rect 21028 40236 21756 40292
rect 21812 40236 21822 40292
rect 9762 40124 9772 40180
rect 9828 40124 11228 40180
rect 11284 40124 11294 40180
rect 15698 40124 15708 40180
rect 15764 40124 21420 40180
rect 21476 40124 21486 40180
rect 21970 40124 21980 40180
rect 22036 40124 22764 40180
rect 22820 40124 22830 40180
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 19618 39900 19628 39956
rect 19684 39900 21308 39956
rect 21364 39900 21374 39956
rect 19478 39788 19516 39844
rect 19572 39788 19582 39844
rect 19842 39788 19852 39844
rect 19908 39788 19918 39844
rect 20066 39788 20076 39844
rect 20132 39788 20636 39844
rect 20692 39788 20702 39844
rect 0 39732 800 39760
rect 0 39676 1708 39732
rect 1764 39676 1774 39732
rect 0 39648 800 39676
rect 19852 39620 19908 39788
rect 29586 39676 29596 39732
rect 29652 39676 30828 39732
rect 30884 39676 30894 39732
rect 2034 39564 2044 39620
rect 2100 39564 9548 39620
rect 9604 39564 9614 39620
rect 19852 39564 20300 39620
rect 20356 39564 20366 39620
rect 21522 39564 21532 39620
rect 21588 39564 22988 39620
rect 23044 39564 23054 39620
rect 6962 39452 6972 39508
rect 7028 39452 8204 39508
rect 8260 39452 13692 39508
rect 13748 39452 16044 39508
rect 16100 39452 17388 39508
rect 17444 39452 17454 39508
rect 19394 39452 19404 39508
rect 19460 39452 19852 39508
rect 19908 39452 19918 39508
rect 20626 39452 20636 39508
rect 20692 39452 22428 39508
rect 22484 39452 22494 39508
rect 22754 39452 22764 39508
rect 22820 39452 23324 39508
rect 23380 39452 23390 39508
rect 2034 39340 2044 39396
rect 2100 39340 8092 39396
rect 8148 39340 8158 39396
rect 19628 39340 19740 39396
rect 19796 39340 19806 39396
rect 14018 39228 14028 39284
rect 14084 39228 17388 39284
rect 17444 39228 19180 39284
rect 19236 39228 19246 39284
rect 19628 39172 19684 39340
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 8194 39116 8204 39172
rect 8260 39116 9660 39172
rect 9716 39116 10332 39172
rect 10388 39116 10398 39172
rect 19618 39116 19628 39172
rect 19684 39116 19694 39172
rect 23202 39116 23212 39172
rect 23268 39116 25340 39172
rect 25396 39116 25406 39172
rect 27010 39116 27020 39172
rect 27076 39116 27086 39172
rect 0 39060 800 39088
rect 0 39004 1708 39060
rect 1764 39004 2492 39060
rect 2548 39004 2558 39060
rect 7522 39004 7532 39060
rect 7588 39004 9436 39060
rect 9492 39004 9502 39060
rect 9762 39004 9772 39060
rect 9828 39004 10892 39060
rect 10948 39004 12572 39060
rect 12628 39004 13244 39060
rect 13300 39004 13310 39060
rect 18386 39004 18396 39060
rect 18452 39004 19516 39060
rect 19572 39004 20636 39060
rect 20692 39004 20702 39060
rect 0 38976 800 39004
rect 7634 38892 7644 38948
rect 7700 38892 9884 38948
rect 9940 38892 9950 38948
rect 12674 38892 12684 38948
rect 12740 38892 14028 38948
rect 14084 38892 14700 38948
rect 14756 38892 14766 38948
rect 17826 38892 17836 38948
rect 17892 38892 19068 38948
rect 19124 38892 19134 38948
rect 8418 38780 8428 38836
rect 8484 38780 8764 38836
rect 8820 38780 8830 38836
rect 16258 38780 16268 38836
rect 16324 38780 18284 38836
rect 18340 38780 18844 38836
rect 18900 38780 18910 38836
rect 19618 38780 19628 38836
rect 19684 38780 20412 38836
rect 20468 38780 20478 38836
rect 22754 38780 22764 38836
rect 22820 38780 23660 38836
rect 23716 38780 25228 38836
rect 25284 38780 25294 38836
rect 27020 38724 27076 39116
rect 39200 39060 40000 39088
rect 34962 39004 34972 39060
rect 35028 39004 40000 39060
rect 39200 38976 40000 39004
rect 22082 38668 22092 38724
rect 22148 38668 24444 38724
rect 24500 38668 24780 38724
rect 24836 38668 24846 38724
rect 27010 38668 27020 38724
rect 27076 38668 27086 38724
rect 26450 38556 26460 38612
rect 26516 38556 27132 38612
rect 27188 38556 27198 38612
rect 32386 38556 32396 38612
rect 32452 38556 33404 38612
rect 33460 38556 33470 38612
rect 17938 38444 17948 38500
rect 18004 38444 19180 38500
rect 19236 38444 19246 38500
rect 24210 38444 24220 38500
rect 24276 38444 25564 38500
rect 25620 38444 25630 38500
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 24742 38220 24780 38276
rect 24836 38220 24846 38276
rect 25442 38220 25452 38276
rect 25508 38220 26012 38276
rect 26068 38220 26908 38276
rect 26964 38220 28028 38276
rect 28084 38220 28094 38276
rect 14914 38108 14924 38164
rect 14980 38108 15148 38164
rect 20066 38108 20076 38164
rect 20132 38108 20748 38164
rect 20804 38108 22092 38164
rect 22148 38108 22158 38164
rect 27682 38108 27692 38164
rect 27748 38108 32396 38164
rect 32452 38108 32462 38164
rect 15092 38052 15148 38108
rect 13122 37996 13132 38052
rect 13188 37996 14028 38052
rect 14084 37996 14094 38052
rect 15092 37996 22652 38052
rect 22708 37996 22718 38052
rect 24882 37996 24892 38052
rect 24948 37996 26236 38052
rect 26292 37996 26684 38052
rect 26740 37996 26750 38052
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 7858 37436 7868 37492
rect 7924 37436 8764 37492
rect 8820 37436 8830 37492
rect 20132 37436 21308 37492
rect 21364 37436 21374 37492
rect 20132 37156 20188 37436
rect 26450 37324 26460 37380
rect 26516 37324 27356 37380
rect 27412 37324 27422 37380
rect 19954 37100 19964 37156
rect 20020 37100 20188 37156
rect 26898 36988 26908 37044
rect 26964 36988 27692 37044
rect 27748 36988 27758 37044
rect 25218 36876 25228 36932
rect 25284 36876 26796 36932
rect 26852 36876 26862 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 27122 36652 27132 36708
rect 27188 36652 27580 36708
rect 27636 36652 27646 36708
rect 39200 36372 40000 36400
rect 38210 36316 38220 36372
rect 38276 36316 40000 36372
rect 39200 36288 40000 36316
rect 8082 36204 8092 36260
rect 8148 36204 10332 36260
rect 10388 36204 11340 36260
rect 11396 36204 11406 36260
rect 27346 36204 27356 36260
rect 27412 36204 28028 36260
rect 28084 36204 28924 36260
rect 28980 36204 29820 36260
rect 29876 36204 29886 36260
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 21858 35868 21868 35924
rect 21924 35868 22540 35924
rect 22596 35868 22606 35924
rect 15092 35756 15260 35812
rect 15316 35756 16156 35812
rect 16212 35756 16222 35812
rect 15092 35588 15148 35756
rect 14354 35532 14364 35588
rect 14420 35532 15148 35588
rect 15810 35532 15820 35588
rect 15876 35532 25228 35588
rect 25284 35532 25294 35588
rect 22194 35420 22204 35476
rect 22260 35420 25340 35476
rect 25396 35420 25406 35476
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 22194 35196 22204 35252
rect 22260 35196 22876 35252
rect 22932 35196 23100 35252
rect 23156 35196 23436 35252
rect 23492 35196 23502 35252
rect 24434 35196 24444 35252
rect 24500 35196 27132 35252
rect 27188 35196 27198 35252
rect 12226 35084 12236 35140
rect 12292 35084 13468 35140
rect 13524 35084 13534 35140
rect 22754 35084 22764 35140
rect 22820 35084 25564 35140
rect 25620 35084 25630 35140
rect 22642 34972 22652 35028
rect 22708 34972 25004 35028
rect 25060 34972 25070 35028
rect 14354 34860 14364 34916
rect 14420 34860 15260 34916
rect 15316 34860 15326 34916
rect 16818 34860 16828 34916
rect 16884 34860 17388 34916
rect 17444 34860 17454 34916
rect 13570 34748 13580 34804
rect 13636 34748 14252 34804
rect 14308 34748 14318 34804
rect 14130 34636 14140 34692
rect 14196 34636 15036 34692
rect 15092 34636 15102 34692
rect 15250 34636 15260 34692
rect 15316 34636 16380 34692
rect 16436 34636 16940 34692
rect 16996 34636 19628 34692
rect 19684 34636 19694 34692
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 21074 34300 21084 34356
rect 21140 34300 21756 34356
rect 21812 34300 21822 34356
rect 24658 34300 24668 34356
rect 24724 34300 25452 34356
rect 25508 34300 25518 34356
rect 15362 34188 15372 34244
rect 15428 34188 16380 34244
rect 16436 34188 16446 34244
rect 20066 34188 20076 34244
rect 20132 34188 21924 34244
rect 16034 34076 16044 34132
rect 16100 34076 16828 34132
rect 16884 34076 16894 34132
rect 20132 34076 20636 34132
rect 20692 34076 21644 34132
rect 21700 34076 21710 34132
rect 20132 34020 20188 34076
rect 21868 34020 21924 34188
rect 14690 33964 14700 34020
rect 14756 33964 15372 34020
rect 15428 33964 16268 34020
rect 16324 33964 16334 34020
rect 16594 33964 16604 34020
rect 16660 33964 17724 34020
rect 17780 33964 17790 34020
rect 19142 33964 19180 34020
rect 19236 33964 20188 34020
rect 21410 33964 21420 34020
rect 21476 33964 22092 34020
rect 22148 33964 22158 34020
rect 14466 33852 14476 33908
rect 14532 33852 15596 33908
rect 15652 33852 15662 33908
rect 20626 33852 20636 33908
rect 20692 33852 22428 33908
rect 22484 33852 22494 33908
rect 20132 33740 21420 33796
rect 21476 33740 24668 33796
rect 24724 33740 24734 33796
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 17154 33628 17164 33684
rect 17220 33628 19068 33684
rect 19124 33628 19740 33684
rect 19796 33628 19806 33684
rect 20132 33572 20188 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 20514 33628 20524 33684
rect 20580 33628 21532 33684
rect 21588 33628 21598 33684
rect 12562 33516 12572 33572
rect 12628 33516 13916 33572
rect 13972 33516 13982 33572
rect 17826 33516 17836 33572
rect 17892 33516 18732 33572
rect 18788 33516 20188 33572
rect 13682 33404 13692 33460
rect 13748 33404 14028 33460
rect 14084 33404 15484 33460
rect 15540 33404 15550 33460
rect 19282 33404 19292 33460
rect 19348 33404 20076 33460
rect 20132 33404 20142 33460
rect 26338 33404 26348 33460
rect 26404 33404 26796 33460
rect 26852 33404 27244 33460
rect 27300 33404 27310 33460
rect 14130 33292 14140 33348
rect 14196 33292 14812 33348
rect 14868 33292 16828 33348
rect 16884 33292 16894 33348
rect 18946 33292 18956 33348
rect 19012 33292 20300 33348
rect 20356 33292 20366 33348
rect 14242 33180 14252 33236
rect 14308 33180 14924 33236
rect 14980 33180 14990 33236
rect 1698 33068 1708 33124
rect 1764 33068 1774 33124
rect 20066 33068 20076 33124
rect 20132 33068 20300 33124
rect 20356 33068 20366 33124
rect 26114 33068 26124 33124
rect 26180 33068 27468 33124
rect 27524 33068 27534 33124
rect 0 33012 800 33040
rect 1708 33012 1764 33068
rect 0 32956 1764 33012
rect 0 32928 800 32956
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 22754 32732 22764 32788
rect 22820 32732 23548 32788
rect 23604 32732 24220 32788
rect 24276 32732 24286 32788
rect 23202 32508 23212 32564
rect 23268 32508 24332 32564
rect 24388 32508 24398 32564
rect 26338 32508 26348 32564
rect 26404 32508 28140 32564
rect 28196 32508 28206 32564
rect 18610 32396 18620 32452
rect 18676 32396 19628 32452
rect 19684 32396 19694 32452
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 14914 31948 14924 32004
rect 14980 31948 15260 32004
rect 15316 31948 22540 32004
rect 22596 31948 23212 32004
rect 23268 31948 23278 32004
rect 25442 31948 25452 32004
rect 25508 31948 26236 32004
rect 26292 31948 26302 32004
rect 18610 31836 18620 31892
rect 18676 31836 20748 31892
rect 20804 31836 21756 31892
rect 21812 31836 21822 31892
rect 14466 31724 14476 31780
rect 14532 31724 15484 31780
rect 15540 31724 15550 31780
rect 12114 31612 12124 31668
rect 12180 31612 14364 31668
rect 14420 31612 14430 31668
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 39200 30996 40000 31024
rect 11442 30940 11452 30996
rect 11508 30940 14700 30996
rect 14756 30940 14766 30996
rect 17490 30940 17500 30996
rect 17556 30940 18620 30996
rect 18676 30940 18686 30996
rect 24658 30940 24668 30996
rect 24724 30940 25228 30996
rect 25284 30940 25294 30996
rect 27010 30940 27020 30996
rect 27076 30940 40000 30996
rect 39200 30912 40000 30940
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 39200 30324 40000 30352
rect 23202 30268 23212 30324
rect 23268 30268 24220 30324
rect 24276 30268 24286 30324
rect 38210 30268 38220 30324
rect 38276 30268 40000 30324
rect 39200 30240 40000 30268
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 39200 22932 40000 22960
rect 38210 22876 38220 22932
rect 38276 22876 40000 22932
rect 39200 22848 40000 22876
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
<< via3 >>
rect 4476 96404 4532 96460
rect 4580 96404 4636 96460
rect 4684 96404 4740 96460
rect 35196 96404 35252 96460
rect 35300 96404 35356 96460
rect 35404 96404 35460 96460
rect 19836 95620 19892 95676
rect 19940 95620 19996 95676
rect 20044 95620 20100 95676
rect 4476 94836 4532 94892
rect 4580 94836 4636 94892
rect 4684 94836 4740 94892
rect 35196 94836 35252 94892
rect 35300 94836 35356 94892
rect 35404 94836 35460 94892
rect 19836 94052 19892 94108
rect 19940 94052 19996 94108
rect 20044 94052 20100 94108
rect 4476 93268 4532 93324
rect 4580 93268 4636 93324
rect 4684 93268 4740 93324
rect 35196 93268 35252 93324
rect 35300 93268 35356 93324
rect 35404 93268 35460 93324
rect 19836 92484 19892 92540
rect 19940 92484 19996 92540
rect 20044 92484 20100 92540
rect 4476 91700 4532 91756
rect 4580 91700 4636 91756
rect 4684 91700 4740 91756
rect 35196 91700 35252 91756
rect 35300 91700 35356 91756
rect 35404 91700 35460 91756
rect 19836 90916 19892 90972
rect 19940 90916 19996 90972
rect 20044 90916 20100 90972
rect 4476 90132 4532 90188
rect 4580 90132 4636 90188
rect 4684 90132 4740 90188
rect 35196 90132 35252 90188
rect 35300 90132 35356 90188
rect 35404 90132 35460 90188
rect 19836 89348 19892 89404
rect 19940 89348 19996 89404
rect 20044 89348 20100 89404
rect 4476 88564 4532 88620
rect 4580 88564 4636 88620
rect 4684 88564 4740 88620
rect 35196 88564 35252 88620
rect 35300 88564 35356 88620
rect 35404 88564 35460 88620
rect 19836 87780 19892 87836
rect 19940 87780 19996 87836
rect 20044 87780 20100 87836
rect 4476 86996 4532 87052
rect 4580 86996 4636 87052
rect 4684 86996 4740 87052
rect 35196 86996 35252 87052
rect 35300 86996 35356 87052
rect 35404 86996 35460 87052
rect 19836 86212 19892 86268
rect 19940 86212 19996 86268
rect 20044 86212 20100 86268
rect 4476 85428 4532 85484
rect 4580 85428 4636 85484
rect 4684 85428 4740 85484
rect 35196 85428 35252 85484
rect 35300 85428 35356 85484
rect 35404 85428 35460 85484
rect 19836 84644 19892 84700
rect 19940 84644 19996 84700
rect 20044 84644 20100 84700
rect 4476 83860 4532 83916
rect 4580 83860 4636 83916
rect 4684 83860 4740 83916
rect 35196 83860 35252 83916
rect 35300 83860 35356 83916
rect 35404 83860 35460 83916
rect 19836 83076 19892 83132
rect 19940 83076 19996 83132
rect 20044 83076 20100 83132
rect 4476 82292 4532 82348
rect 4580 82292 4636 82348
rect 4684 82292 4740 82348
rect 35196 82292 35252 82348
rect 35300 82292 35356 82348
rect 35404 82292 35460 82348
rect 19836 81508 19892 81564
rect 19940 81508 19996 81564
rect 20044 81508 20100 81564
rect 4476 80724 4532 80780
rect 4580 80724 4636 80780
rect 4684 80724 4740 80780
rect 35196 80724 35252 80780
rect 35300 80724 35356 80780
rect 35404 80724 35460 80780
rect 19836 79940 19892 79996
rect 19940 79940 19996 79996
rect 20044 79940 20100 79996
rect 4476 79156 4532 79212
rect 4580 79156 4636 79212
rect 4684 79156 4740 79212
rect 35196 79156 35252 79212
rect 35300 79156 35356 79212
rect 35404 79156 35460 79212
rect 19836 78372 19892 78428
rect 19940 78372 19996 78428
rect 20044 78372 20100 78428
rect 4476 77588 4532 77644
rect 4580 77588 4636 77644
rect 4684 77588 4740 77644
rect 35196 77588 35252 77644
rect 35300 77588 35356 77644
rect 35404 77588 35460 77644
rect 19836 76804 19892 76860
rect 19940 76804 19996 76860
rect 20044 76804 20100 76860
rect 4476 76020 4532 76076
rect 4580 76020 4636 76076
rect 4684 76020 4740 76076
rect 35196 76020 35252 76076
rect 35300 76020 35356 76076
rect 35404 76020 35460 76076
rect 19836 75236 19892 75292
rect 19940 75236 19996 75292
rect 20044 75236 20100 75292
rect 4476 74452 4532 74508
rect 4580 74452 4636 74508
rect 4684 74452 4740 74508
rect 35196 74452 35252 74508
rect 35300 74452 35356 74508
rect 35404 74452 35460 74508
rect 19836 73668 19892 73724
rect 19940 73668 19996 73724
rect 20044 73668 20100 73724
rect 4476 72884 4532 72940
rect 4580 72884 4636 72940
rect 4684 72884 4740 72940
rect 35196 72884 35252 72940
rect 35300 72884 35356 72940
rect 35404 72884 35460 72940
rect 19836 72100 19892 72156
rect 19940 72100 19996 72156
rect 20044 72100 20100 72156
rect 4476 71316 4532 71372
rect 4580 71316 4636 71372
rect 4684 71316 4740 71372
rect 35196 71316 35252 71372
rect 35300 71316 35356 71372
rect 35404 71316 35460 71372
rect 19836 70532 19892 70588
rect 19940 70532 19996 70588
rect 20044 70532 20100 70588
rect 4476 69748 4532 69804
rect 4580 69748 4636 69804
rect 4684 69748 4740 69804
rect 35196 69748 35252 69804
rect 35300 69748 35356 69804
rect 35404 69748 35460 69804
rect 19836 68964 19892 69020
rect 19940 68964 19996 69020
rect 20044 68964 20100 69020
rect 4476 68180 4532 68236
rect 4580 68180 4636 68236
rect 4684 68180 4740 68236
rect 35196 68180 35252 68236
rect 35300 68180 35356 68236
rect 35404 68180 35460 68236
rect 19836 67396 19892 67452
rect 19940 67396 19996 67452
rect 20044 67396 20100 67452
rect 4476 66612 4532 66668
rect 4580 66612 4636 66668
rect 4684 66612 4740 66668
rect 35196 66612 35252 66668
rect 35300 66612 35356 66668
rect 35404 66612 35460 66668
rect 19836 65828 19892 65884
rect 19940 65828 19996 65884
rect 20044 65828 20100 65884
rect 4476 65044 4532 65100
rect 4580 65044 4636 65100
rect 4684 65044 4740 65100
rect 35196 65044 35252 65100
rect 35300 65044 35356 65100
rect 35404 65044 35460 65100
rect 19836 64260 19892 64316
rect 19940 64260 19996 64316
rect 20044 64260 20100 64316
rect 4476 63476 4532 63532
rect 4580 63476 4636 63532
rect 4684 63476 4740 63532
rect 35196 63476 35252 63532
rect 35300 63476 35356 63532
rect 35404 63476 35460 63532
rect 19836 62692 19892 62748
rect 19940 62692 19996 62748
rect 20044 62692 20100 62748
rect 19628 62300 19684 62356
rect 4476 61908 4532 61964
rect 4580 61908 4636 61964
rect 4684 61908 4740 61964
rect 35196 61908 35252 61964
rect 35300 61908 35356 61964
rect 35404 61908 35460 61964
rect 19516 61740 19572 61796
rect 19628 61180 19684 61236
rect 19836 61124 19892 61180
rect 19940 61124 19996 61180
rect 20044 61124 20100 61180
rect 19516 60844 19572 60900
rect 19628 60620 19684 60676
rect 4476 60340 4532 60396
rect 4580 60340 4636 60396
rect 4684 60340 4740 60396
rect 35196 60340 35252 60396
rect 35300 60340 35356 60396
rect 35404 60340 35460 60396
rect 19836 59556 19892 59612
rect 19940 59556 19996 59612
rect 20044 59556 20100 59612
rect 4476 58772 4532 58828
rect 4580 58772 4636 58828
rect 4684 58772 4740 58828
rect 35196 58772 35252 58828
rect 35300 58772 35356 58828
rect 35404 58772 35460 58828
rect 25564 58492 25620 58548
rect 25676 58380 25732 58436
rect 19836 57988 19892 58044
rect 19940 57988 19996 58044
rect 20044 57988 20100 58044
rect 18844 57372 18900 57428
rect 4476 57204 4532 57260
rect 4580 57204 4636 57260
rect 4684 57204 4740 57260
rect 35196 57204 35252 57260
rect 35300 57204 35356 57260
rect 35404 57204 35460 57260
rect 25676 56700 25732 56756
rect 25564 56588 25620 56644
rect 19836 56420 19892 56476
rect 19940 56420 19996 56476
rect 20044 56420 20100 56476
rect 4476 55636 4532 55692
rect 4580 55636 4636 55692
rect 4684 55636 4740 55692
rect 35196 55636 35252 55692
rect 35300 55636 35356 55692
rect 35404 55636 35460 55692
rect 19836 54852 19892 54908
rect 19940 54852 19996 54908
rect 20044 54852 20100 54908
rect 4476 54068 4532 54124
rect 4580 54068 4636 54124
rect 4684 54068 4740 54124
rect 35196 54068 35252 54124
rect 35300 54068 35356 54124
rect 35404 54068 35460 54124
rect 19836 53284 19892 53340
rect 19940 53284 19996 53340
rect 20044 53284 20100 53340
rect 22204 52780 22260 52836
rect 4476 52500 4532 52556
rect 4580 52500 4636 52556
rect 4684 52500 4740 52556
rect 35196 52500 35252 52556
rect 35300 52500 35356 52556
rect 35404 52500 35460 52556
rect 21868 52108 21924 52164
rect 22092 51772 22148 51828
rect 19836 51716 19892 51772
rect 19940 51716 19996 51772
rect 20044 51716 20100 51772
rect 4476 50932 4532 50988
rect 4580 50932 4636 50988
rect 4684 50932 4740 50988
rect 35196 50932 35252 50988
rect 35300 50932 35356 50988
rect 35404 50932 35460 50988
rect 19836 50148 19892 50204
rect 19940 50148 19996 50204
rect 20044 50148 20100 50204
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 34860 48972 34916 49028
rect 34860 48636 34916 48692
rect 19836 48580 19892 48636
rect 19940 48580 19996 48636
rect 20044 48580 20100 48636
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 19180 46620 19236 46676
rect 22092 46620 22148 46676
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 21868 45276 21924 45332
rect 19628 45052 19684 45108
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 18620 44156 18676 44212
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 22204 43596 22260 43652
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 18844 41692 18900 41748
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 22764 41468 22820 41524
rect 24780 41020 24836 41076
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 18620 40236 18676 40292
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 19516 39788 19572 39844
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 19516 39004 19572 39060
rect 22764 38780 22820 38836
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 24780 38220 24836 38276
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 19180 33964 19236 34020
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 96460 4768 96492
rect 4448 96404 4476 96460
rect 4532 96404 4580 96460
rect 4636 96404 4684 96460
rect 4740 96404 4768 96460
rect 4448 94892 4768 96404
rect 4448 94836 4476 94892
rect 4532 94836 4580 94892
rect 4636 94836 4684 94892
rect 4740 94836 4768 94892
rect 4448 93324 4768 94836
rect 4448 93268 4476 93324
rect 4532 93268 4580 93324
rect 4636 93268 4684 93324
rect 4740 93268 4768 93324
rect 4448 91756 4768 93268
rect 4448 91700 4476 91756
rect 4532 91700 4580 91756
rect 4636 91700 4684 91756
rect 4740 91700 4768 91756
rect 4448 90188 4768 91700
rect 4448 90132 4476 90188
rect 4532 90132 4580 90188
rect 4636 90132 4684 90188
rect 4740 90132 4768 90188
rect 4448 88620 4768 90132
rect 4448 88564 4476 88620
rect 4532 88564 4580 88620
rect 4636 88564 4684 88620
rect 4740 88564 4768 88620
rect 4448 87052 4768 88564
rect 4448 86996 4476 87052
rect 4532 86996 4580 87052
rect 4636 86996 4684 87052
rect 4740 86996 4768 87052
rect 4448 85484 4768 86996
rect 4448 85428 4476 85484
rect 4532 85428 4580 85484
rect 4636 85428 4684 85484
rect 4740 85428 4768 85484
rect 4448 83916 4768 85428
rect 4448 83860 4476 83916
rect 4532 83860 4580 83916
rect 4636 83860 4684 83916
rect 4740 83860 4768 83916
rect 4448 82348 4768 83860
rect 4448 82292 4476 82348
rect 4532 82292 4580 82348
rect 4636 82292 4684 82348
rect 4740 82292 4768 82348
rect 4448 80780 4768 82292
rect 4448 80724 4476 80780
rect 4532 80724 4580 80780
rect 4636 80724 4684 80780
rect 4740 80724 4768 80780
rect 4448 79212 4768 80724
rect 4448 79156 4476 79212
rect 4532 79156 4580 79212
rect 4636 79156 4684 79212
rect 4740 79156 4768 79212
rect 4448 77644 4768 79156
rect 4448 77588 4476 77644
rect 4532 77588 4580 77644
rect 4636 77588 4684 77644
rect 4740 77588 4768 77644
rect 4448 76076 4768 77588
rect 4448 76020 4476 76076
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4740 76020 4768 76076
rect 4448 74508 4768 76020
rect 4448 74452 4476 74508
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4740 74452 4768 74508
rect 4448 72940 4768 74452
rect 4448 72884 4476 72940
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4740 72884 4768 72940
rect 4448 71372 4768 72884
rect 4448 71316 4476 71372
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4740 71316 4768 71372
rect 4448 69804 4768 71316
rect 4448 69748 4476 69804
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4740 69748 4768 69804
rect 4448 68236 4768 69748
rect 4448 68180 4476 68236
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4740 68180 4768 68236
rect 4448 66668 4768 68180
rect 4448 66612 4476 66668
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4740 66612 4768 66668
rect 4448 65100 4768 66612
rect 4448 65044 4476 65100
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4740 65044 4768 65100
rect 4448 63532 4768 65044
rect 4448 63476 4476 63532
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4740 63476 4768 63532
rect 4448 61964 4768 63476
rect 19808 95676 20128 96492
rect 19808 95620 19836 95676
rect 19892 95620 19940 95676
rect 19996 95620 20044 95676
rect 20100 95620 20128 95676
rect 19808 94108 20128 95620
rect 19808 94052 19836 94108
rect 19892 94052 19940 94108
rect 19996 94052 20044 94108
rect 20100 94052 20128 94108
rect 19808 92540 20128 94052
rect 19808 92484 19836 92540
rect 19892 92484 19940 92540
rect 19996 92484 20044 92540
rect 20100 92484 20128 92540
rect 19808 90972 20128 92484
rect 19808 90916 19836 90972
rect 19892 90916 19940 90972
rect 19996 90916 20044 90972
rect 20100 90916 20128 90972
rect 19808 89404 20128 90916
rect 19808 89348 19836 89404
rect 19892 89348 19940 89404
rect 19996 89348 20044 89404
rect 20100 89348 20128 89404
rect 19808 87836 20128 89348
rect 19808 87780 19836 87836
rect 19892 87780 19940 87836
rect 19996 87780 20044 87836
rect 20100 87780 20128 87836
rect 19808 86268 20128 87780
rect 19808 86212 19836 86268
rect 19892 86212 19940 86268
rect 19996 86212 20044 86268
rect 20100 86212 20128 86268
rect 19808 84700 20128 86212
rect 19808 84644 19836 84700
rect 19892 84644 19940 84700
rect 19996 84644 20044 84700
rect 20100 84644 20128 84700
rect 19808 83132 20128 84644
rect 19808 83076 19836 83132
rect 19892 83076 19940 83132
rect 19996 83076 20044 83132
rect 20100 83076 20128 83132
rect 19808 81564 20128 83076
rect 19808 81508 19836 81564
rect 19892 81508 19940 81564
rect 19996 81508 20044 81564
rect 20100 81508 20128 81564
rect 19808 79996 20128 81508
rect 19808 79940 19836 79996
rect 19892 79940 19940 79996
rect 19996 79940 20044 79996
rect 20100 79940 20128 79996
rect 19808 78428 20128 79940
rect 19808 78372 19836 78428
rect 19892 78372 19940 78428
rect 19996 78372 20044 78428
rect 20100 78372 20128 78428
rect 19808 76860 20128 78372
rect 19808 76804 19836 76860
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 20100 76804 20128 76860
rect 19808 75292 20128 76804
rect 19808 75236 19836 75292
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 20100 75236 20128 75292
rect 19808 73724 20128 75236
rect 19808 73668 19836 73724
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 20100 73668 20128 73724
rect 19808 72156 20128 73668
rect 19808 72100 19836 72156
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 20100 72100 20128 72156
rect 19808 70588 20128 72100
rect 19808 70532 19836 70588
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 20100 70532 20128 70588
rect 19808 69020 20128 70532
rect 19808 68964 19836 69020
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 20100 68964 20128 69020
rect 19808 67452 20128 68964
rect 19808 67396 19836 67452
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 20100 67396 20128 67452
rect 19808 65884 20128 67396
rect 19808 65828 19836 65884
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 20100 65828 20128 65884
rect 19808 64316 20128 65828
rect 19808 64260 19836 64316
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 20100 64260 20128 64316
rect 19808 62748 20128 64260
rect 19808 62692 19836 62748
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 20100 62692 20128 62748
rect 4448 61908 4476 61964
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4740 61908 4768 61964
rect 4448 60396 4768 61908
rect 19628 62356 19684 62366
rect 19516 61796 19572 61806
rect 19516 60900 19572 61740
rect 19628 61236 19684 62300
rect 19628 61170 19684 61180
rect 19808 61180 20128 62692
rect 19516 60834 19572 60844
rect 19808 61124 19836 61180
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 20100 61124 20128 61180
rect 4448 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4768 60396
rect 4448 58828 4768 60340
rect 4448 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4768 58828
rect 4448 57260 4768 58772
rect 19628 60676 19684 60686
rect 4448 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4768 57260
rect 4448 55692 4768 57204
rect 4448 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4768 55692
rect 4448 54124 4768 55636
rect 4448 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4768 54124
rect 4448 52556 4768 54068
rect 4448 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4768 52556
rect 4448 50988 4768 52500
rect 4448 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4768 50988
rect 4448 49420 4768 50932
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 4448 47852 4768 49364
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4448 46284 4768 47796
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 18844 57428 18900 57438
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 18620 44212 18676 44222
rect 18620 40292 18676 44156
rect 18844 41748 18900 57372
rect 18844 41682 18900 41692
rect 19180 46676 19236 46686
rect 18620 40226 18676 40236
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 19180 34020 19236 46620
rect 19628 45108 19684 60620
rect 19628 45042 19684 45052
rect 19808 59612 20128 61124
rect 19808 59556 19836 59612
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 20100 59556 20128 59612
rect 19808 58044 20128 59556
rect 35168 96460 35488 96492
rect 35168 96404 35196 96460
rect 35252 96404 35300 96460
rect 35356 96404 35404 96460
rect 35460 96404 35488 96460
rect 35168 94892 35488 96404
rect 35168 94836 35196 94892
rect 35252 94836 35300 94892
rect 35356 94836 35404 94892
rect 35460 94836 35488 94892
rect 35168 93324 35488 94836
rect 35168 93268 35196 93324
rect 35252 93268 35300 93324
rect 35356 93268 35404 93324
rect 35460 93268 35488 93324
rect 35168 91756 35488 93268
rect 35168 91700 35196 91756
rect 35252 91700 35300 91756
rect 35356 91700 35404 91756
rect 35460 91700 35488 91756
rect 35168 90188 35488 91700
rect 35168 90132 35196 90188
rect 35252 90132 35300 90188
rect 35356 90132 35404 90188
rect 35460 90132 35488 90188
rect 35168 88620 35488 90132
rect 35168 88564 35196 88620
rect 35252 88564 35300 88620
rect 35356 88564 35404 88620
rect 35460 88564 35488 88620
rect 35168 87052 35488 88564
rect 35168 86996 35196 87052
rect 35252 86996 35300 87052
rect 35356 86996 35404 87052
rect 35460 86996 35488 87052
rect 35168 85484 35488 86996
rect 35168 85428 35196 85484
rect 35252 85428 35300 85484
rect 35356 85428 35404 85484
rect 35460 85428 35488 85484
rect 35168 83916 35488 85428
rect 35168 83860 35196 83916
rect 35252 83860 35300 83916
rect 35356 83860 35404 83916
rect 35460 83860 35488 83916
rect 35168 82348 35488 83860
rect 35168 82292 35196 82348
rect 35252 82292 35300 82348
rect 35356 82292 35404 82348
rect 35460 82292 35488 82348
rect 35168 80780 35488 82292
rect 35168 80724 35196 80780
rect 35252 80724 35300 80780
rect 35356 80724 35404 80780
rect 35460 80724 35488 80780
rect 35168 79212 35488 80724
rect 35168 79156 35196 79212
rect 35252 79156 35300 79212
rect 35356 79156 35404 79212
rect 35460 79156 35488 79212
rect 35168 77644 35488 79156
rect 35168 77588 35196 77644
rect 35252 77588 35300 77644
rect 35356 77588 35404 77644
rect 35460 77588 35488 77644
rect 35168 76076 35488 77588
rect 35168 76020 35196 76076
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35460 76020 35488 76076
rect 35168 74508 35488 76020
rect 35168 74452 35196 74508
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35460 74452 35488 74508
rect 35168 72940 35488 74452
rect 35168 72884 35196 72940
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35460 72884 35488 72940
rect 35168 71372 35488 72884
rect 35168 71316 35196 71372
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35460 71316 35488 71372
rect 35168 69804 35488 71316
rect 35168 69748 35196 69804
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35460 69748 35488 69804
rect 35168 68236 35488 69748
rect 35168 68180 35196 68236
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35460 68180 35488 68236
rect 35168 66668 35488 68180
rect 35168 66612 35196 66668
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35460 66612 35488 66668
rect 35168 65100 35488 66612
rect 35168 65044 35196 65100
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35460 65044 35488 65100
rect 35168 63532 35488 65044
rect 35168 63476 35196 63532
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35460 63476 35488 63532
rect 35168 61964 35488 63476
rect 35168 61908 35196 61964
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35460 61908 35488 61964
rect 35168 60396 35488 61908
rect 35168 60340 35196 60396
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35460 60340 35488 60396
rect 35168 58828 35488 60340
rect 35168 58772 35196 58828
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35460 58772 35488 58828
rect 19808 57988 19836 58044
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20100 57988 20128 58044
rect 19808 56476 20128 57988
rect 25564 58548 25620 58558
rect 25564 56644 25620 58492
rect 25676 58436 25732 58446
rect 25676 56756 25732 58380
rect 25676 56690 25732 56700
rect 35168 57260 35488 58772
rect 35168 57204 35196 57260
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35460 57204 35488 57260
rect 25564 56578 25620 56588
rect 19808 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20128 56476
rect 19808 54908 20128 56420
rect 19808 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20128 54908
rect 19808 53340 20128 54852
rect 19808 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20128 53340
rect 19808 51772 20128 53284
rect 35168 55692 35488 57204
rect 35168 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35488 55692
rect 35168 54124 35488 55636
rect 35168 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35488 54124
rect 22204 52836 22260 52846
rect 19808 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20128 51772
rect 19808 50204 20128 51716
rect 19808 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20128 50204
rect 19808 48636 20128 50148
rect 19808 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20128 48636
rect 19808 47068 20128 48580
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 19808 45500 20128 47012
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19808 43932 20128 45444
rect 21868 52164 21924 52174
rect 21868 45332 21924 52108
rect 22092 51828 22148 51838
rect 22092 46676 22148 51772
rect 22092 46610 22148 46620
rect 21868 45266 21924 45276
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 22204 43652 22260 52780
rect 35168 52556 35488 54068
rect 35168 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35488 52556
rect 35168 50988 35488 52500
rect 35168 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35488 50988
rect 35168 49420 35488 50932
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 34860 49028 34916 49038
rect 34860 48692 34916 48972
rect 34860 48626 34916 48636
rect 22204 43586 22260 43596
rect 35168 47852 35488 49364
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 35168 46284 35488 47796
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19516 39844 19572 39854
rect 19516 39060 19572 39788
rect 19516 38994 19572 39004
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19180 33954 19236 33964
rect 19808 37660 20128 39172
rect 22764 41524 22820 41534
rect 22764 38836 22820 41468
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 22764 38770 22820 38780
rect 24780 41076 24836 41086
rect 24780 38276 24836 41020
rect 24780 38210 24836 38220
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _386_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10080 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _387_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 26656 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _388_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 32704 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _389_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 31472 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _390_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19488 0 1 67424
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _391_
timestamp 1698175906
transform 1 0 14672 0 1 59584
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  _392_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16016 0 -1 58016
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _393_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 16800 0 -1 54880
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _394_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 15456 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _395_
timestamp 1698175906
transform -1 0 19152 0 1 53312
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _396_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15680 0 1 50176
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__and3_2  _397_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15344 0 1 48608
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _398_
timestamp 1698175906
transform 1 0 13440 0 1 43904
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _399_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 14336 0 -1 40768
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _400_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15904 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _401_
timestamp 1698175906
transform -1 0 24304 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _402_
timestamp 1698175906
transform 1 0 12432 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _403_
timestamp 1698175906
transform -1 0 16016 0 -1 58016
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _404_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19040 0 -1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _405_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15008 0 -1 50176
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _406_
timestamp 1698175906
transform 1 0 14672 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _407_
timestamp 1698175906
transform 1 0 14672 0 1 39200
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _408_
timestamp 1698175906
transform 1 0 12880 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _409_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13888 0 1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _410_
timestamp 1698175906
transform -1 0 23408 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _411_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 24080 0 1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or3_2  _412_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 23184 0 -1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _413_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 24080 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _414_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 -1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _415_
timestamp 1698175906
transform -1 0 15792 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _416_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16128 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _417_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 17808 0 1 56448
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _418_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 -1 56448
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _419_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21504 0 1 54880
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _420_
timestamp 1698175906
transform 1 0 13328 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _421_
timestamp 1698175906
transform -1 0 15232 0 -1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _422_
timestamp 1698175906
transform 1 0 13776 0 1 67424
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _423_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16352 0 1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or4_2  _424_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 -1 67424
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _425_
timestamp 1698175906
transform 1 0 19824 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _426_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18368 0 1 62720
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _427_
timestamp 1698175906
transform -1 0 15904 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _428_
timestamp 1698175906
transform 1 0 18368 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _429_
timestamp 1698175906
transform 1 0 17248 0 -1 62720
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _430_
timestamp 1698175906
transform 1 0 18928 0 -1 62720
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _431_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17136 0 1 62720
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _432_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20048 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _433_
timestamp 1698175906
transform -1 0 17024 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _434_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 16016 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _435_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20832 0 1 67424
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _436_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20048 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _437_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19712 0 -1 70560
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _438_
timestamp 1698175906
transform 1 0 17248 0 -1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _439_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17920 0 -1 68992
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _440_
timestamp 1698175906
transform 1 0 17808 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _441_
timestamp 1698175906
transform 1 0 17360 0 1 68992
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _442_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 22064 0 -1 67424
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _443_
timestamp 1698175906
transform -1 0 23520 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _444_
timestamp 1698175906
transform 1 0 17248 0 -1 59584
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _445_
timestamp 1698175906
transform -1 0 19488 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _446_
timestamp 1698175906
transform 1 0 17248 0 -1 64288
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _447_
timestamp 1698175906
transform -1 0 20048 0 1 59584
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__or4_2  _448_
timestamp 1698175906
transform 1 0 20496 0 -1 61152
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _449_
timestamp 1698175906
transform 1 0 18256 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _450_
timestamp 1698175906
transform 1 0 17248 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _451_
timestamp 1698175906
transform -1 0 13104 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _452_
timestamp 1698175906
transform 1 0 13776 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _453_
timestamp 1698175906
transform -1 0 14896 0 -1 45472
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _454_
timestamp 1698175906
transform 1 0 18256 0 -1 45472
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _455_
timestamp 1698175906
transform -1 0 16800 0 -1 42336
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _456_
timestamp 1698175906
transform -1 0 14896 0 1 42336
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _457_
timestamp 1698175906
transform 1 0 14448 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _458_
timestamp 1698175906
transform 1 0 16800 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _459_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20272 0 -1 43904
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__and3_2  _460_
timestamp 1698175906
transform 1 0 19040 0 1 43904
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _461_
timestamp 1698175906
transform -1 0 17024 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _462_
timestamp 1698175906
transform -1 0 17024 0 -1 53312
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _463_
timestamp 1698175906
transform 1 0 15904 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _464_
timestamp 1698175906
transform 1 0 14672 0 -1 53312
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _465_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 14896 0 1 51744
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _466_
timestamp 1698175906
transform 1 0 25088 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _467_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 22624 0 -1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _468_
timestamp 1698175906
transform 1 0 21728 0 1 51744
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _469_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 27104 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _470_
timestamp 1698175906
transform 1 0 19040 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _471_
timestamp 1698175906
transform 1 0 19152 0 1 53312
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _472_
timestamp 1698175906
transform 1 0 19152 0 -1 53312
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _473_
timestamp 1698175906
transform 1 0 15232 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _474_
timestamp 1698175906
transform -1 0 18592 0 1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _475_
timestamp 1698175906
transform 1 0 15120 0 1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _476_
timestamp 1698175906
transform 1 0 20160 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _477_
timestamp 1698175906
transform 1 0 21616 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_4  _478_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20944 0 1 50176
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _479_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21840 0 -1 51744
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _480_
timestamp 1698175906
transform 1 0 23744 0 -1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _481_
timestamp 1698175906
transform 1 0 18368 0 -1 54880
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _482_
timestamp 1698175906
transform -1 0 23968 0 1 48608
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _483_
timestamp 1698175906
transform -1 0 14672 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _484_
timestamp 1698175906
transform 1 0 17024 0 1 58016
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _485_
timestamp 1698175906
transform 1 0 21168 0 1 56448
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _486_
timestamp 1698175906
transform 1 0 22288 0 1 53312
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _487_
timestamp 1698175906
transform -1 0 24304 0 -1 50176
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _488_
timestamp 1698175906
transform 1 0 13328 0 -1 39200
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _489_
timestamp 1698175906
transform -1 0 18816 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _490_
timestamp 1698175906
transform -1 0 19040 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _491_
timestamp 1698175906
transform 1 0 17472 0 -1 45472
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _492_
timestamp 1698175906
transform -1 0 17024 0 -1 45472
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _493_
timestamp 1698175906
transform 1 0 19488 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _494_
timestamp 1698175906
transform -1 0 20384 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _495_
timestamp 1698175906
transform 1 0 17248 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _496_
timestamp 1698175906
transform 1 0 18032 0 -1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _497_
timestamp 1698175906
transform 1 0 18816 0 -1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _498_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19824 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _499_
timestamp 1698175906
transform 1 0 21168 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _500_
timestamp 1698175906
transform -1 0 19040 0 1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _501_
timestamp 1698175906
transform 1 0 15680 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_4  _502_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 17024 0 -1 43904
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _503_
timestamp 1698175906
transform 1 0 16016 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _504_
timestamp 1698175906
transform -1 0 18704 0 -1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _505_
timestamp 1698175906
transform 1 0 18704 0 -1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _506_
timestamp 1698175906
transform 1 0 15568 0 1 36064
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _507_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19936 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _508_
timestamp 1698175906
transform 1 0 21168 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _509_
timestamp 1698175906
transform -1 0 15904 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _510_
timestamp 1698175906
transform 1 0 16912 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _511_
timestamp 1698175906
transform 1 0 17584 0 -1 50176
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _512_
timestamp 1698175906
transform 1 0 19488 0 -1 40768
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _513_
timestamp 1698175906
transform 1 0 22848 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _514_
timestamp 1698175906
transform 1 0 17472 0 1 48608
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _515_
timestamp 1698175906
transform 1 0 19936 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _516_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20272 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _517_
timestamp 1698175906
transform -1 0 25536 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _518_
timestamp 1698175906
transform 1 0 21392 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _519_
timestamp 1698175906
transform 1 0 21840 0 1 45472
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _520_
timestamp 1698175906
transform -1 0 19040 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _521_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _522_
timestamp 1698175906
transform -1 0 24864 0 -1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _523_
timestamp 1698175906
transform -1 0 24864 0 -1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or4_2  _524_
timestamp 1698175906
transform 1 0 21168 0 -1 40768
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__or4_2  _525_
timestamp 1698175906
transform 1 0 25088 0 -1 42336
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _526_
timestamp 1698175906
transform -1 0 32256 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _527_
timestamp 1698175906
transform -1 0 31136 0 1 40768
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _528_
timestamp 1698175906
transform -1 0 31696 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _529_
timestamp 1698175906
transform -1 0 30912 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _530_
timestamp 1698175906
transform 1 0 28560 0 -1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _531_
timestamp 1698175906
transform -1 0 28112 0 1 40768
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _532_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 29792 0 -1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and3_2  _533_
timestamp 1698175906
transform 1 0 31360 0 -1 42336
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _534_
timestamp 1698175906
transform 1 0 33040 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _535_
timestamp 1698175906
transform 1 0 27328 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _536_
timestamp 1698175906
transform -1 0 31360 0 -1 42336
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _537_
timestamp 1698175906
transform 1 0 19488 0 1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _538_
timestamp 1698175906
transform 1 0 17696 0 -1 61152
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _539_
timestamp 1698175906
transform 1 0 19600 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _540_
timestamp 1698175906
transform 1 0 20272 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _541_
timestamp 1698175906
transform 1 0 25088 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _542_
timestamp 1698175906
transform 1 0 22624 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _543_
timestamp 1698175906
transform -1 0 22400 0 -1 62720
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _544_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21168 0 -1 53312
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _545_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21056 0 -1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _546_
timestamp 1698175906
transform 1 0 22512 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _547_
timestamp 1698175906
transform -1 0 22288 0 -1 56448
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _548_
timestamp 1698175906
transform -1 0 21840 0 -1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _549_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 26544 0 1 39200
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _550_
timestamp 1698175906
transform -1 0 23072 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _551_
timestamp 1698175906
transform -1 0 22848 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _552_
timestamp 1698175906
transform 1 0 19600 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _553_
timestamp 1698175906
transform 1 0 21168 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _554_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21392 0 1 40768
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _555_
timestamp 1698175906
transform 1 0 20832 0 -1 50176
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _556_
timestamp 1698175906
transform 1 0 21056 0 -1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _557_
timestamp 1698175906
transform -1 0 22064 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _558_
timestamp 1698175906
transform 1 0 20272 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _559_
timestamp 1698175906
transform 1 0 22064 0 -1 48608
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _560_
timestamp 1698175906
transform 1 0 23072 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _561_
timestamp 1698175906
transform -1 0 30912 0 1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _562_
timestamp 1698175906
transform -1 0 32704 0 -1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _563_
timestamp 1698175906
transform 1 0 31472 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _564_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 31136 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _565_
timestamp 1698175906
transform -1 0 28560 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _566_
timestamp 1698175906
transform 1 0 23184 0 -1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _567_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 30688 0 1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _568_
timestamp 1698175906
transform 1 0 31136 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _569_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 31696 0 -1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _570_
timestamp 1698175906
transform 1 0 29008 0 -1 45472
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _571_
timestamp 1698175906
transform 1 0 29792 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _572_
timestamp 1698175906
transform 1 0 30688 0 1 47040
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _573_
timestamp 1698175906
transform 1 0 31920 0 1 42336
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _574_
timestamp 1698175906
transform 1 0 28224 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _575_
timestamp 1698175906
transform 1 0 28224 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _576_
timestamp 1698175906
transform 1 0 29456 0 -1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _577_
timestamp 1698175906
transform 1 0 32928 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _578_
timestamp 1698175906
transform 1 0 32704 0 1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _579_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 33600 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _580_
timestamp 1698175906
transform -1 0 32032 0 -1 48608
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _581_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 33824 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _582_
timestamp 1698175906
transform -1 0 33152 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _583_
timestamp 1698175906
transform 1 0 33600 0 -1 47040
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _584_
timestamp 1698175906
transform 1 0 33152 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _585_
timestamp 1698175906
transform -1 0 31808 0 -1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _586_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 35952 0 1 47040
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _587_
timestamp 1698175906
transform -1 0 33712 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _588_
timestamp 1698175906
transform 1 0 33600 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _589_
timestamp 1698175906
transform 1 0 33040 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _590_
timestamp 1698175906
transform 1 0 32480 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _591_
timestamp 1698175906
transform 1 0 34048 0 -1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or3_4  _592_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 32928 0 -1 48608
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _593_
timestamp 1698175906
transform -1 0 34720 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _594_
timestamp 1698175906
transform -1 0 35056 0 -1 45472
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _595_
timestamp 1698175906
transform 1 0 31808 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _596_
timestamp 1698175906
transform 1 0 34272 0 1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _597_
timestamp 1698175906
transform 1 0 32032 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _598_
timestamp 1698175906
transform -1 0 36288 0 1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _599_
timestamp 1698175906
transform 1 0 10080 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _600_
timestamp 1698175906
transform 1 0 11760 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _601_
timestamp 1698175906
transform 1 0 12432 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _602_
timestamp 1698175906
transform 1 0 9856 0 1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _603_
timestamp 1698175906
transform 1 0 9744 0 1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _604_
timestamp 1698175906
transform 1 0 11872 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _605_
timestamp 1698175906
transform 1 0 14224 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _606_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13552 0 1 64288
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _607_
timestamp 1698175906
transform 1 0 10864 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _608_
timestamp 1698175906
transform -1 0 13104 0 1 65856
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _609_
timestamp 1698175906
transform -1 0 8848 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _610_
timestamp 1698175906
transform 1 0 8176 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _611_
timestamp 1698175906
transform 1 0 9744 0 1 65856
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _612_
timestamp 1698175906
transform 1 0 9520 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _613_
timestamp 1698175906
transform 1 0 10752 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _614_
timestamp 1698175906
transform -1 0 13104 0 1 67424
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _615_
timestamp 1698175906
transform 1 0 7616 0 -1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _616_
timestamp 1698175906
transform 1 0 9520 0 -1 68992
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _617_
timestamp 1698175906
transform 1 0 11648 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _618_
timestamp 1698175906
transform -1 0 10864 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _619_
timestamp 1698175906
transform -1 0 10416 0 -1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _620_
timestamp 1698175906
transform 1 0 8624 0 -1 67424
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _621_
timestamp 1698175906
transform 1 0 8064 0 -1 67424
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _622_
timestamp 1698175906
transform 1 0 9408 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _623_
timestamp 1698175906
transform -1 0 11648 0 -1 64288
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _624_
timestamp 1698175906
transform 1 0 8512 0 1 64288
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _625_
timestamp 1698175906
transform 1 0 10192 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _626_
timestamp 1698175906
transform -1 0 10640 0 1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _627_
timestamp 1698175906
transform 1 0 8736 0 1 62720
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _628_
timestamp 1698175906
transform -1 0 9744 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _629_
timestamp 1698175906
transform -1 0 9184 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _630_
timestamp 1698175906
transform 1 0 13552 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _631_
timestamp 1698175906
transform -1 0 14560 0 -1 62720
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _632_
timestamp 1698175906
transform 1 0 10976 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _633_
timestamp 1698175906
transform 1 0 13328 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _634_
timestamp 1698175906
transform -1 0 14448 0 1 58016
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _635_
timestamp 1698175906
transform 1 0 12880 0 -1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _636_
timestamp 1698175906
transform -1 0 14448 0 1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _637_
timestamp 1698175906
transform -1 0 9968 0 -1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _638_
timestamp 1698175906
transform -1 0 10080 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _639_
timestamp 1698175906
transform 1 0 7616 0 -1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _640_
timestamp 1698175906
transform 1 0 7728 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _641_
timestamp 1698175906
transform -1 0 7840 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _642_
timestamp 1698175906
transform 1 0 7056 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _643_
timestamp 1698175906
transform 1 0 10080 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _644_
timestamp 1698175906
transform 1 0 9744 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _645_
timestamp 1698175906
transform 1 0 9296 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _646_
timestamp 1698175906
transform -1 0 7952 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _647_
timestamp 1698175906
transform -1 0 10304 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _648_
timestamp 1698175906
transform 1 0 8624 0 -1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _649_
timestamp 1698175906
transform 1 0 7616 0 -1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _650_
timestamp 1698175906
transform 1 0 9408 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _651_
timestamp 1698175906
transform 1 0 11312 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _652_
timestamp 1698175906
transform -1 0 13104 0 1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _653_
timestamp 1698175906
transform 1 0 6496 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _654_
timestamp 1698175906
transform -1 0 10864 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _655_
timestamp 1698175906
transform 1 0 8176 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _656_
timestamp 1698175906
transform -1 0 7168 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _657_
timestamp 1698175906
transform -1 0 9856 0 1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _658_
timestamp 1698175906
transform 1 0 7280 0 1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _659_
timestamp 1698175906
transform 1 0 7840 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _660_
timestamp 1698175906
transform 1 0 11312 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _661_
timestamp 1698175906
transform -1 0 13104 0 1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _662_
timestamp 1698175906
transform 1 0 11088 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _663_
timestamp 1698175906
transform -1 0 12096 0 -1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _664_
timestamp 1698175906
transform -1 0 11088 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _665_
timestamp 1698175906
transform 1 0 9408 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _666_
timestamp 1698175906
transform 1 0 10080 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _667_
timestamp 1698175906
transform 1 0 6496 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _668_
timestamp 1698175906
transform 1 0 8064 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _669_
timestamp 1698175906
transform -1 0 7168 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _670_
timestamp 1698175906
transform -1 0 9968 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _671_
timestamp 1698175906
transform 1 0 7840 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _672_
timestamp 1698175906
transform 1 0 8288 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _673_
timestamp 1698175906
transform 1 0 7952 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _674_
timestamp 1698175906
transform 1 0 9968 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _675_
timestamp 1698175906
transform 1 0 8064 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _676_
timestamp 1698175906
transform 1 0 8512 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _677_
timestamp 1698175906
transform 1 0 9408 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _678_
timestamp 1698175906
transform -1 0 9856 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _679_
timestamp 1698175906
transform 1 0 7392 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _680_
timestamp 1698175906
transform 1 0 9520 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _681_
timestamp 1698175906
transform -1 0 11648 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _682_
timestamp 1698175906
transform -1 0 11648 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _683_
timestamp 1698175906
transform 1 0 7392 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _684_
timestamp 1698175906
transform -1 0 10976 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _685_
timestamp 1698175906
transform -1 0 8512 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _686_
timestamp 1698175906
transform 1 0 23408 0 1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _687_
timestamp 1698175906
transform -1 0 28896 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _688_
timestamp 1698175906
transform -1 0 28336 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _689_
timestamp 1698175906
transform -1 0 26320 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _690_
timestamp 1698175906
transform -1 0 25760 0 -1 70560
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _691_
timestamp 1698175906
transform -1 0 26656 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _692_
timestamp 1698175906
transform -1 0 25088 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _693_
timestamp 1698175906
transform 1 0 24192 0 -1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _694_
timestamp 1698175906
transform -1 0 25424 0 1 67424
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _695_
timestamp 1698175906
transform -1 0 24864 0 -1 65856
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _696_
timestamp 1698175906
transform 1 0 22736 0 -1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _697_
timestamp 1698175906
transform -1 0 27664 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _698_
timestamp 1698175906
transform 1 0 25536 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _699_
timestamp 1698175906
transform 1 0 25424 0 1 68992
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _700_
timestamp 1698175906
transform -1 0 25984 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _701_
timestamp 1698175906
transform 1 0 26096 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _702_
timestamp 1698175906
transform -1 0 27104 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _703_
timestamp 1698175906
transform 1 0 25088 0 -1 67424
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _704_
timestamp 1698175906
transform 1 0 27216 0 -1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _705_
timestamp 1698175906
transform -1 0 27216 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _706_
timestamp 1698175906
transform -1 0 24864 0 -1 62720
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _707_
timestamp 1698175906
transform -1 0 25984 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _708_
timestamp 1698175906
transform -1 0 25424 0 1 62720
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _709_
timestamp 1698175906
transform -1 0 24192 0 1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _710_
timestamp 1698175906
transform 1 0 25760 0 1 62720
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _711_
timestamp 1698175906
transform 1 0 27104 0 1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _712_
timestamp 1698175906
transform 1 0 25088 0 1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _713_
timestamp 1698175906
transform -1 0 25312 0 1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _714_
timestamp 1698175906
transform 1 0 23744 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _715_
timestamp 1698175906
transform -1 0 25088 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _716_
timestamp 1698175906
transform 1 0 24640 0 1 59584
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _717_
timestamp 1698175906
transform 1 0 26096 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _718_
timestamp 1698175906
transform 1 0 22960 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _719_
timestamp 1698175906
transform 1 0 23856 0 1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _720_
timestamp 1698175906
transform 1 0 24976 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _721_
timestamp 1698175906
transform 1 0 25312 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _722_
timestamp 1698175906
transform 1 0 26320 0 1 56448
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _723_
timestamp 1698175906
transform 1 0 27104 0 1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _724_
timestamp 1698175906
transform 1 0 24304 0 -1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _725_
timestamp 1698175906
transform 1 0 25200 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _726_
timestamp 1698175906
transform 1 0 29008 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _727_
timestamp 1698175906
transform -1 0 28672 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _728_
timestamp 1698175906
transform -1 0 27776 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _729_
timestamp 1698175906
transform 1 0 24640 0 1 54880
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _730_
timestamp 1698175906
transform -1 0 27328 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _731_
timestamp 1698175906
transform 1 0 24192 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _732_
timestamp 1698175906
transform -1 0 27104 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _733_
timestamp 1698175906
transform -1 0 26432 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _734_
timestamp 1698175906
transform -1 0 26096 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _735_
timestamp 1698175906
transform 1 0 25088 0 1 42336
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _736_
timestamp 1698175906
transform -1 0 26432 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _737_
timestamp 1698175906
transform 1 0 25984 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _738_
timestamp 1698175906
transform 1 0 26880 0 -1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _739_
timestamp 1698175906
transform -1 0 27776 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _740_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 26880 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _741_
timestamp 1698175906
transform 1 0 25088 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _742_
timestamp 1698175906
transform 1 0 25872 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _743_
timestamp 1698175906
transform -1 0 22400 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _744_
timestamp 1698175906
transform -1 0 22512 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _745_
timestamp 1698175906
transform -1 0 21840 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _746_
timestamp 1698175906
transform -1 0 22064 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _747_
timestamp 1698175906
transform 1 0 21504 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _748_
timestamp 1698175906
transform 1 0 23744 0 -1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _749_
timestamp 1698175906
transform 1 0 25088 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _750_
timestamp 1698175906
transform -1 0 20608 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _751_
timestamp 1698175906
transform -1 0 20944 0 -1 34496
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _752_
timestamp 1698175906
transform -1 0 19376 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _753_
timestamp 1698175906
transform 1 0 17248 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _754_
timestamp 1698175906
transform -1 0 17584 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _755_
timestamp 1698175906
transform 1 0 17248 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _756_
timestamp 1698175906
transform -1 0 15456 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _757_
timestamp 1698175906
transform 1 0 14896 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _758_
timestamp 1698175906
transform 1 0 14000 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _759_
timestamp 1698175906
transform -1 0 13776 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _760_
timestamp 1698175906
transform 1 0 14672 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _761_
timestamp 1698175906
transform -1 0 16800 0 -1 34496
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _762_
timestamp 1698175906
transform -1 0 14672 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _763_
timestamp 1698175906
transform -1 0 14560 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _764_
timestamp 1698175906
transform 1 0 14560 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _765_
timestamp 1698175906
transform -1 0 15120 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _766_
timestamp 1698175906
transform 1 0 23072 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _767_
timestamp 1698175906
transform 1 0 22400 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _768_
timestamp 1698175906
transform 1 0 21728 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _769_
timestamp 1698175906
transform -1 0 24528 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _770_
timestamp 1698175906
transform 1 0 23520 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _771_
timestamp 1698175906
transform 1 0 25088 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _772_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 32592 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _773_
timestamp 1698175906
transform -1 0 31472 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _774_
timestamp 1698175906
transform -1 0 32256 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _775_
timestamp 1698175906
transform 1 0 32928 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _776_
timestamp 1698175906
transform 1 0 13552 0 -1 68992
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _777_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10080 0 -1 68992
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _778_
timestamp 1698175906
transform 1 0 10752 0 -1 67424
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _779_
timestamp 1698175906
transform -1 0 10752 0 1 67424
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_4  _780_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9072 0 1 64288
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _781_
timestamp 1698175906
transform 1 0 9408 0 -1 62720
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _782_
timestamp 1698175906
transform 1 0 13328 0 1 62720
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _783_
timestamp 1698175906
transform 1 0 11984 0 -1 59584
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _784_
timestamp 1698175906
transform 1 0 11760 0 -1 54880
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _785_
timestamp 1698175906
transform 1 0 5824 0 1 59584
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _786_
timestamp 1698175906
transform 1 0 5936 0 -1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _787_
timestamp 1698175906
transform 1 0 5712 0 -1 56448
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _788_
timestamp 1698175906
transform 1 0 11536 0 -1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _789_
timestamp 1698175906
transform 1 0 5040 0 -1 50176
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _790_
timestamp 1698175906
transform 1 0 6048 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _791_
timestamp 1698175906
transform 1 0 11760 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _792_
timestamp 1698175906
transform 1 0 9856 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _793_
timestamp 1698175906
transform 1 0 9856 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _794_
timestamp 1698175906
transform 1 0 5040 0 -1 43904
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _795_
timestamp 1698175906
transform 1 0 6384 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _796_
timestamp 1698175906
transform -1 0 10080 0 1 37632
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _797_
timestamp 1698175906
transform 1 0 7840 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _798_
timestamp 1698175906
transform 1 0 9856 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _799_
timestamp 1698175906
transform 1 0 6832 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _800_
timestamp 1698175906
transform -1 0 25424 0 1 68992
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _801_
timestamp 1698175906
transform -1 0 24192 0 -1 68992
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _802_
timestamp 1698175906
transform -1 0 29232 0 -1 68992
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _803_
timestamp 1698175906
transform 1 0 25536 0 1 67424
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _804_
timestamp 1698175906
transform -1 0 24528 0 -1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _805_
timestamp 1698175906
transform 1 0 26544 0 -1 64288
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _806_
timestamp 1698175906
transform -1 0 28784 0 -1 61152
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _807_
timestamp 1698175906
transform -1 0 24640 0 -1 58016
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _808_
timestamp 1698175906
transform 1 0 26880 0 -1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _809_
timestamp 1698175906
transform 1 0 26880 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _810_
timestamp 1698175906
transform 1 0 25648 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _811_
timestamp 1698175906
transform -1 0 27776 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _812_
timestamp 1698175906
transform -1 0 28336 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _813_
timestamp 1698175906
transform 1 0 26768 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _814_
timestamp 1698175906
transform -1 0 28448 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _815_
timestamp 1698175906
transform -1 0 22064 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _816_
timestamp 1698175906
transform -1 0 27328 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _817_
timestamp 1698175906
transform 1 0 17248 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _818_
timestamp 1698175906
transform 1 0 16128 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _819_
timestamp 1698175906
transform 1 0 11312 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _820_
timestamp 1698175906
transform 1 0 11648 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _821_
timestamp 1698175906
transform 1 0 11200 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _822_
timestamp 1698175906
transform 1 0 21168 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _823_
timestamp 1698175906
transform -1 0 26544 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _824_
timestamp 1698175906
transform 1 0 33264 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _825_
timestamp 1698175906
transform 1 0 32928 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _826_
timestamp 1698175906
transform 1 0 35168 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _827_
timestamp 1698175906
transform 1 0 35168 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _828_
timestamp 1698175906
transform 1 0 35168 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _829_
timestamp 1698175906
transform 1 0 35168 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _830_
timestamp 1698175906
transform 1 0 34720 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__386__A2 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9856 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__387__I
timestamp 1698175906
transform -1 0 26656 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__407__A2
timestamp 1698175906
transform 1 0 18816 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__455__I
timestamp 1698175906
transform 1 0 17472 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__479__B2
timestamp 1698175906
transform 1 0 24640 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__484__B
timestamp 1698175906
transform 1 0 18928 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__514__A2
timestamp 1698175906
transform 1 0 20384 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__522__A2
timestamp 1698175906
transform 1 0 23296 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__535__I
timestamp 1698175906
transform -1 0 27328 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__602__I
timestamp 1698175906
transform -1 0 9856 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__606__B
timestamp 1698175906
transform 1 0 13328 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__608__A1
timestamp 1698175906
transform 1 0 12320 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__611__A1
timestamp 1698175906
transform -1 0 9744 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__614__A1
timestamp 1698175906
transform 1 0 13552 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__631__B
timestamp 1698175906
transform 1 0 13216 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__644__I
timestamp 1698175906
transform 1 0 8960 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__666__B
timestamp 1698175906
transform -1 0 11424 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__672__B
timestamp 1698175906
transform 1 0 9184 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__673__A1
timestamp 1698175906
transform 1 0 10640 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__674__I
timestamp 1698175906
transform -1 0 9968 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__677__A1
timestamp 1698175906
transform -1 0 10416 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__680__A1
timestamp 1698175906
transform 1 0 10304 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__681__A1
timestamp 1698175906
transform 1 0 11872 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__684__A2
timestamp 1698175906
transform 1 0 11200 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__689__I
timestamp 1698175906
transform 1 0 26768 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__690__A2
timestamp 1698175906
transform -1 0 26208 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__695__A1
timestamp 1698175906
transform 1 0 25312 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__695__A2
timestamp 1698175906
transform 1 0 25760 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__698__I
timestamp 1698175906
transform 1 0 27328 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__701__A1
timestamp 1698175906
transform 1 0 27216 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__702__I
timestamp 1698175906
transform 1 0 27776 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__708__A1
timestamp 1698175906
transform 1 0 26208 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__708__A2
timestamp 1698175906
transform 1 0 25648 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__711__A1
timestamp 1698175906
transform 1 0 28000 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__716__A1
timestamp 1698175906
transform 1 0 25872 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__716__A2
timestamp 1698175906
transform 1 0 24416 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__723__A1
timestamp 1698175906
transform 1 0 26880 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__730__A3
timestamp 1698175906
transform 1 0 27552 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__731__I
timestamp 1698175906
transform 1 0 24864 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__732__A2
timestamp 1698175906
transform 1 0 28000 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__733__A2
timestamp 1698175906
transform -1 0 25536 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__736__A1
timestamp 1698175906
transform 1 0 25536 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__738__A1
timestamp 1698175906
transform 1 0 28896 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__739__A1
timestamp 1698175906
transform 1 0 26880 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__740__A3
timestamp 1698175906
transform 1 0 28000 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__740__A4
timestamp 1698175906
transform 1 0 28448 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__742__A1
timestamp 1698175906
transform 1 0 26768 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__747__A1
timestamp 1698175906
transform 1 0 23072 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__748__A1
timestamp 1698175906
transform -1 0 25088 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__748__A2
timestamp 1698175906
transform 1 0 25312 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__750__A1
timestamp 1698175906
transform 1 0 22288 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__751__A2
timestamp 1698175906
transform 1 0 22736 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__757__B
timestamp 1698175906
transform 1 0 15792 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__762__A1
timestamp 1698175906
transform -1 0 13776 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__765__A1
timestamp 1698175906
transform -1 0 15568 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__766__B
timestamp 1698175906
transform 1 0 23968 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__771__A1
timestamp 1698175906
transform -1 0 26208 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__796__CLK
timestamp 1698175906
transform 1 0 10304 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__797__CLK
timestamp 1698175906
transform 1 0 11312 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__815__CLK
timestamp 1698175906
transform 1 0 18592 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__817__CLK
timestamp 1698175906
transform 1 0 20720 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__818__CLK
timestamp 1698175906
transform 1 0 19600 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__819__CLK
timestamp 1698175906
transform 1 0 14560 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__820__CLK
timestamp 1698175906
transform 1 0 15120 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__821__CLK
timestamp 1698175906
transform 1 0 14672 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__822__CLK
timestamp 1698175906
transform -1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform 1 0 26992 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_0__f_clk_I
timestamp 1698175906
transform -1 0 22176 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_1__f_clk_I
timestamp 1698175906
transform 1 0 20608 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_2__f_clk_I
timestamp 1698175906
transform 1 0 29568 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_3__f_clk_I
timestamp 1698175906
transform 1 0 30576 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_4__f_clk_I
timestamp 1698175906
transform 1 0 18032 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_5__f_clk_I
timestamp 1698175906
transform 1 0 17472 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_6__f_clk_I
timestamp 1698175906
transform 1 0 25648 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_7__f_clk_I
timestamp 1698175906
transform -1 0 24304 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698175906
transform 1 0 3136 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698175906
transform 1 0 2912 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698175906
transform 1 0 2464 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698175906
transform 1 0 2464 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698175906
transform 1 0 2464 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698175906
transform 1 0 2464 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698175906
transform 1 0 2464 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698175906
transform 1 0 2464 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698175906
transform 1 0 3136 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698175906
transform 1 0 2464 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698175906
transform 1 0 2464 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698175906
transform 1 0 2464 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698175906
transform 1 0 2464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698175906
transform 1 0 2464 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698175906
transform 1 0 2464 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698175906
transform 1 0 2464 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698175906
transform 1 0 2464 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1698175906
transform 1 0 2464 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1698175906
transform -1 0 2240 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1698175906
transform 1 0 2464 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1698175906
transform 1 0 2464 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1698175906
transform 1 0 2464 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1698175906
transform 1 0 2464 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1698175906
transform 1 0 2464 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1698175906
transform 1 0 2464 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1698175906
transform 1 0 2464 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 26768 0 1 50176
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_0__f_clk
timestamp 1698175906
transform -1 0 20944 0 1 37632
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_1__f_clk
timestamp 1698175906
transform -1 0 19376 0 1 40768
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_2__f_clk
timestamp 1698175906
transform 1 0 29792 0 1 39200
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_3__f_clk
timestamp 1698175906
transform 1 0 30800 0 1 43904
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_4__f_clk
timestamp 1698175906
transform -1 0 17024 0 -1 56448
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_5__f_clk
timestamp 1698175906
transform -1 0 17024 0 -1 61152
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_6__f_clk
timestamp 1698175906
transform 1 0 25872 0 -1 58016
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_7__f_clk
timestamp 1698175906
transform -1 0 30688 0 -1 62720
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_2 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_10 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 2464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_12 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 2688 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_17 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 3248 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_33
timestamp 1698175906
transform 1 0 5040 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_138
timestamp 1698175906
transform 1 0 16800 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_172
timestamp 1698175906
transform 1 0 20608 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_206
timestamp 1698175906
transform 1 0 24416 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_308
timestamp 1698175906
transform 1 0 35840 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_324 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 37632 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_328
timestamp 1698175906
transform 1 0 38080 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_330
timestamp 1698175906
transform 1 0 38304 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_142
timestamp 1698175906
transform 1 0 17248 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_206
timestamp 1698175906
transform 1 0 24416 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_212
timestamp 1698175906
transform 1 0 25088 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_276
timestamp 1698175906
transform 1 0 32256 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_282
timestamp 1698175906
transform 1 0 32928 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_314
timestamp 1698175906
transform 1 0 36512 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_330
timestamp 1698175906
transform 1 0 38304 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 21168 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 28336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_317
timestamp 1698175906
transform 1 0 36848 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_325
timestamp 1698175906
transform 1 0 37744 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_329
timestamp 1698175906
transform 1 0 38192 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_282
timestamp 1698175906
transform 1 0 32928 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_314
timestamp 1698175906
transform 1 0 36512 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_330
timestamp 1698175906
transform 1 0 38304 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_317
timestamp 1698175906
transform 1 0 36848 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_325
timestamp 1698175906
transform 1 0 37744 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_329
timestamp 1698175906
transform 1 0 38192 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_282
timestamp 1698175906
transform 1 0 32928 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_314
timestamp 1698175906
transform 1 0 36512 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_330
timestamp 1698175906
transform 1 0 38304 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_317
timestamp 1698175906
transform 1 0 36848 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_325
timestamp 1698175906
transform 1 0 37744 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_329
timestamp 1698175906
transform 1 0 38192 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_282
timestamp 1698175906
transform 1 0 32928 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_314
timestamp 1698175906
transform 1 0 36512 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_330
timestamp 1698175906
transform 1 0 38304 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_317
timestamp 1698175906
transform 1 0 36848 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_325
timestamp 1698175906
transform 1 0 37744 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_329
timestamp 1698175906
transform 1 0 38192 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_282
timestamp 1698175906
transform 1 0 32928 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_314
timestamp 1698175906
transform 1 0 36512 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_330
timestamp 1698175906
transform 1 0 38304 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_317
timestamp 1698175906
transform 1 0 36848 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_325
timestamp 1698175906
transform 1 0 37744 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_329
timestamp 1698175906
transform 1 0 38192 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 17248 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_282
timestamp 1698175906
transform 1 0 32928 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_314
timestamp 1698175906
transform 1 0 36512 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_330
timestamp 1698175906
transform 1 0 38304 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_107
timestamp 1698175906
transform 1 0 13328 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698175906
transform 1 0 20496 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698175906
transform 1 0 21168 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698175906
transform 1 0 28336 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_317
timestamp 1698175906
transform 1 0 36848 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_325
timestamp 1698175906
transform 1 0 37744 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_329
timestamp 1698175906
transform 1 0 38192 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698175906
transform 1 0 9408 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698175906
transform 1 0 16576 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_142
timestamp 1698175906
transform 1 0 17248 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_206
timestamp 1698175906
transform 1 0 24416 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698175906
transform 1 0 25088 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698175906
transform 1 0 32256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_282
timestamp 1698175906
transform 1 0 32928 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_314
timestamp 1698175906
transform 1 0 36512 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_330
timestamp 1698175906
transform 1 0 38304 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_107
timestamp 1698175906
transform 1 0 13328 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_171
timestamp 1698175906
transform 1 0 20496 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_177
timestamp 1698175906
transform 1 0 21168 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_241
timestamp 1698175906
transform 1 0 28336 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 29008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 36176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_317
timestamp 1698175906
transform 1 0 36848 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_325
timestamp 1698175906
transform 1 0 37744 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_329
timestamp 1698175906
transform 1 0 38192 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_72
timestamp 1698175906
transform 1 0 9408 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_136
timestamp 1698175906
transform 1 0 16576 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_142
timestamp 1698175906
transform 1 0 17248 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_206
timestamp 1698175906
transform 1 0 24416 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_212
timestamp 1698175906
transform 1 0 25088 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_276
timestamp 1698175906
transform 1 0 32256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_282
timestamp 1698175906
transform 1 0 32928 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_314
timestamp 1698175906
transform 1 0 36512 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_330
timestamp 1698175906
transform 1 0 38304 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_107
timestamp 1698175906
transform 1 0 13328 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_171
timestamp 1698175906
transform 1 0 20496 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_177
timestamp 1698175906
transform 1 0 21168 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_241
timestamp 1698175906
transform 1 0 28336 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 29008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 36176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_317
timestamp 1698175906
transform 1 0 36848 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_325
timestamp 1698175906
transform 1 0 37744 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_329
timestamp 1698175906
transform 1 0 38192 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698175906
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698175906
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_72
timestamp 1698175906
transform 1 0 9408 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_136
timestamp 1698175906
transform 1 0 16576 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_142
timestamp 1698175906
transform 1 0 17248 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_206
timestamp 1698175906
transform 1 0 24416 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_212
timestamp 1698175906
transform 1 0 25088 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_276
timestamp 1698175906
transform 1 0 32256 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_282
timestamp 1698175906
transform 1 0 32928 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_314
timestamp 1698175906
transform 1 0 36512 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_330
timestamp 1698175906
transform 1 0 38304 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698175906
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_107
timestamp 1698175906
transform 1 0 13328 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_171
timestamp 1698175906
transform 1 0 20496 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_177
timestamp 1698175906
transform 1 0 21168 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_241
timestamp 1698175906
transform 1 0 28336 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 29008 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 36176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_317
timestamp 1698175906
transform 1 0 36848 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_325
timestamp 1698175906
transform 1 0 37744 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_329
timestamp 1698175906
transform 1 0 38192 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_72
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_136
timestamp 1698175906
transform 1 0 16576 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_142
timestamp 1698175906
transform 1 0 17248 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_206
timestamp 1698175906
transform 1 0 24416 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_212
timestamp 1698175906
transform 1 0 25088 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_276
timestamp 1698175906
transform 1 0 32256 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_282
timestamp 1698175906
transform 1 0 32928 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_314
timestamp 1698175906
transform 1 0 36512 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_330
timestamp 1698175906
transform 1 0 38304 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698175906
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698175906
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_107
timestamp 1698175906
transform 1 0 13328 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_171
timestamp 1698175906
transform 1 0 20496 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_177
timestamp 1698175906
transform 1 0 21168 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_241
timestamp 1698175906
transform 1 0 28336 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698175906
transform 1 0 29008 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698175906
transform 1 0 36176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_317
timestamp 1698175906
transform 1 0 36848 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_325
timestamp 1698175906
transform 1 0 37744 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_329
timestamp 1698175906
transform 1 0 38192 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_72
timestamp 1698175906
transform 1 0 9408 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_136
timestamp 1698175906
transform 1 0 16576 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_142
timestamp 1698175906
transform 1 0 17248 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_206
timestamp 1698175906
transform 1 0 24416 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_212
timestamp 1698175906
transform 1 0 25088 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_276
timestamp 1698175906
transform 1 0 32256 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698175906
transform 1 0 32928 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_314
timestamp 1698175906
transform 1 0 36512 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_330
timestamp 1698175906
transform 1 0 38304 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698175906
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698175906
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_107
timestamp 1698175906
transform 1 0 13328 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_171
timestamp 1698175906
transform 1 0 20496 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_177
timestamp 1698175906
transform 1 0 21168 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_241
timestamp 1698175906
transform 1 0 28336 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698175906
transform 1 0 29008 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 36176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_317
timestamp 1698175906
transform 1 0 36848 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_325
timestamp 1698175906
transform 1 0 37744 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_329
timestamp 1698175906
transform 1 0 38192 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_72
timestamp 1698175906
transform 1 0 9408 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_136
timestamp 1698175906
transform 1 0 16576 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_142
timestamp 1698175906
transform 1 0 17248 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_206
timestamp 1698175906
transform 1 0 24416 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_212
timestamp 1698175906
transform 1 0 25088 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_276
timestamp 1698175906
transform 1 0 32256 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 32928 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_314
timestamp 1698175906
transform 1 0 36512 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_330
timestamp 1698175906
transform 1 0 38304 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698175906
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_107
timestamp 1698175906
transform 1 0 13328 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_171
timestamp 1698175906
transform 1 0 20496 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_177
timestamp 1698175906
transform 1 0 21168 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_241
timestamp 1698175906
transform 1 0 28336 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 29008 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 36176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_317
timestamp 1698175906
transform 1 0 36848 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_325
timestamp 1698175906
transform 1 0 37744 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_329
timestamp 1698175906
transform 1 0 38192 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698175906
transform 1 0 1568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698175906
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_72
timestamp 1698175906
transform 1 0 9408 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_136
timestamp 1698175906
transform 1 0 16576 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_142
timestamp 1698175906
transform 1 0 17248 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_206
timestamp 1698175906
transform 1 0 24416 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_212
timestamp 1698175906
transform 1 0 25088 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_276
timestamp 1698175906
transform 1 0 32256 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698175906
transform 1 0 32928 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_314
timestamp 1698175906
transform 1 0 36512 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_322
timestamp 1698175906
transform 1 0 37408 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_326
timestamp 1698175906
transform 1 0 37856 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698175906
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_107
timestamp 1698175906
transform 1 0 13328 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_171
timestamp 1698175906
transform 1 0 20496 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_177
timestamp 1698175906
transform 1 0 21168 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_241
timestamp 1698175906
transform 1 0 28336 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 29008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 36176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_317
timestamp 1698175906
transform 1 0 36848 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_325
timestamp 1698175906
transform 1 0 37744 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_329
timestamp 1698175906
transform 1 0 38192 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_72
timestamp 1698175906
transform 1 0 9408 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_136
timestamp 1698175906
transform 1 0 16576 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_142
timestamp 1698175906
transform 1 0 17248 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_206
timestamp 1698175906
transform 1 0 24416 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_212
timestamp 1698175906
transform 1 0 25088 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_276
timestamp 1698175906
transform 1 0 32256 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_282
timestamp 1698175906
transform 1 0 32928 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_314
timestamp 1698175906
transform 1 0 36512 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_330
timestamp 1698175906
transform 1 0 38304 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698175906
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_107
timestamp 1698175906
transform 1 0 13328 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_171
timestamp 1698175906
transform 1 0 20496 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_177
timestamp 1698175906
transform 1 0 21168 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_241
timestamp 1698175906
transform 1 0 28336 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 29008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 36176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_317
timestamp 1698175906
transform 1 0 36848 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_325
timestamp 1698175906
transform 1 0 37744 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_329
timestamp 1698175906
transform 1 0 38192 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698175906
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698175906
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_72
timestamp 1698175906
transform 1 0 9408 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_136
timestamp 1698175906
transform 1 0 16576 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_142
timestamp 1698175906
transform 1 0 17248 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_206
timestamp 1698175906
transform 1 0 24416 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_212
timestamp 1698175906
transform 1 0 25088 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_276
timestamp 1698175906
transform 1 0 32256 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_282
timestamp 1698175906
transform 1 0 32928 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_314
timestamp 1698175906
transform 1 0 36512 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_330
timestamp 1698175906
transform 1 0 38304 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698175906
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_107
timestamp 1698175906
transform 1 0 13328 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_171
timestamp 1698175906
transform 1 0 20496 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_177
timestamp 1698175906
transform 1 0 21168 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_241
timestamp 1698175906
transform 1 0 28336 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 29008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_317
timestamp 1698175906
transform 1 0 36848 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_325
timestamp 1698175906
transform 1 0 37744 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_329
timestamp 1698175906
transform 1 0 38192 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698175906
transform 1 0 9408 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698175906
transform 1 0 16576 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_142
timestamp 1698175906
transform 1 0 17248 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_206
timestamp 1698175906
transform 1 0 24416 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 25088 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 32256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_282
timestamp 1698175906
transform 1 0 32928 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_314
timestamp 1698175906
transform 1 0 36512 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_330
timestamp 1698175906
transform 1 0 38304 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698175906
transform 1 0 13328 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698175906
transform 1 0 20496 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 21168 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 28336 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 29008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_317
timestamp 1698175906
transform 1 0 36848 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_325
timestamp 1698175906
transform 1 0 37744 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_329
timestamp 1698175906
transform 1 0 38192 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 17248 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_282
timestamp 1698175906
transform 1 0 32928 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_314
timestamp 1698175906
transform 1 0 36512 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_330
timestamp 1698175906
transform 1 0 38304 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 13328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_171
timestamp 1698175906
transform 1 0 20496 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_206
timestamp 1698175906
transform 1 0 24416 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_238
timestamp 1698175906
transform 1 0 28000 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_242
timestamp 1698175906
transform 1 0 28448 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_244
timestamp 1698175906
transform 1 0 28672 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 29008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_317
timestamp 1698175906
transform 1 0 36848 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_325
timestamp 1698175906
transform 1 0 37744 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_329
timestamp 1698175906
transform 1 0 38192 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_72
timestamp 1698175906
transform 1 0 9408 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_117
timestamp 1698175906
transform 1 0 14448 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_121
timestamp 1698175906
transform 1 0 14896 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_137
timestamp 1698175906
transform 1 0 16688 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_139
timestamp 1698175906
transform 1 0 16912 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_171
timestamp 1698175906
transform 1 0 20496 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_175
timestamp 1698175906
transform 1 0 20944 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_179
timestamp 1698175906
transform 1 0 21392 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_181
timestamp 1698175906
transform 1 0 21616 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_186
timestamp 1698175906
transform 1 0 22176 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_190
timestamp 1698175906
transform 1 0 22624 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_197
timestamp 1698175906
transform 1 0 23408 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_218
timestamp 1698175906
transform 1 0 25760 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_222
timestamp 1698175906
transform 1 0 26208 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_254
timestamp 1698175906
transform 1 0 29792 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_270
timestamp 1698175906
transform 1 0 31584 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_278
timestamp 1698175906
transform 1 0 32480 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_282
timestamp 1698175906
transform 1 0 32928 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_314
timestamp 1698175906
transform 1 0 36512 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_322
timestamp 1698175906
transform 1 0 37408 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_326
timestamp 1698175906
transform 1 0 37856 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_107
timestamp 1698175906
transform 1 0 13328 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_123
timestamp 1698175906
transform 1 0 15120 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_127
timestamp 1698175906
transform 1 0 15568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_159
timestamp 1698175906
transform 1 0 19152 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_177
timestamp 1698175906
transform 1 0 21168 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_185
timestamp 1698175906
transform 1 0 22064 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_187
timestamp 1698175906
transform 1 0 22288 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_225
timestamp 1698175906
transform 1 0 26544 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 29008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_317
timestamp 1698175906
transform 1 0 36848 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_325
timestamp 1698175906
transform 1 0 37744 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_329
timestamp 1698175906
transform 1 0 38192 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_72
timestamp 1698175906
transform 1 0 9408 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_104
timestamp 1698175906
transform 1 0 12992 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_126
timestamp 1698175906
transform 1 0 15456 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_134
timestamp 1698175906
transform 1 0 16352 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_138
timestamp 1698175906
transform 1 0 16800 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_142
timestamp 1698175906
transform 1 0 17248 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_150
timestamp 1698175906
transform 1 0 18144 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_185
timestamp 1698175906
transform 1 0 22064 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_193
timestamp 1698175906
transform 1 0 22960 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_207
timestamp 1698175906
transform 1 0 24528 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_209
timestamp 1698175906
transform 1 0 24752 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_212
timestamp 1698175906
transform 1 0 25088 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_242
timestamp 1698175906
transform 1 0 28448 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_274
timestamp 1698175906
transform 1 0 32032 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_278
timestamp 1698175906
transform 1 0 32480 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_282
timestamp 1698175906
transform 1 0 32928 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_314
timestamp 1698175906
transform 1 0 36512 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_330
timestamp 1698175906
transform 1 0 38304 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_6
timestamp 1698175906
transform 1 0 2016 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_22
timestamp 1698175906
transform 1 0 3808 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_30
timestamp 1698175906
transform 1 0 4704 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_107
timestamp 1698175906
transform 1 0 13328 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_127
timestamp 1698175906
transform 1 0 15568 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_135
timestamp 1698175906
transform 1 0 16464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_145
timestamp 1698175906
transform 1 0 17584 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_161
timestamp 1698175906
transform 1 0 19376 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_163
timestamp 1698175906
transform 1 0 19600 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_172
timestamp 1698175906
transform 1 0 20608 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_174
timestamp 1698175906
transform 1 0 20832 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_185
timestamp 1698175906
transform 1 0 22064 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_189
timestamp 1698175906
transform 1 0 22512 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_197
timestamp 1698175906
transform 1 0 23408 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_201
timestamp 1698175906
transform 1 0 23856 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_204
timestamp 1698175906
transform 1 0 24192 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_208
timestamp 1698175906
transform 1 0 24640 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_212
timestamp 1698175906
transform 1 0 25088 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_216
timestamp 1698175906
transform 1 0 25536 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_218
timestamp 1698175906
transform 1 0 25760 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_225
timestamp 1698175906
transform 1 0 26544 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_229
timestamp 1698175906
transform 1 0 26992 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 29008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_317
timestamp 1698175906
transform 1 0 36848 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_325
timestamp 1698175906
transform 1 0 37744 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_329
timestamp 1698175906
transform 1 0 38192 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_72
timestamp 1698175906
transform 1 0 9408 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_88
timestamp 1698175906
transform 1 0 11200 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_121
timestamp 1698175906
transform 1 0 14896 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_125
timestamp 1698175906
transform 1 0 15344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_138
timestamp 1698175906
transform 1 0 16800 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_150
timestamp 1698175906
transform 1 0 18144 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_158
timestamp 1698175906
transform 1 0 19040 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_162
timestamp 1698175906
transform 1 0 19488 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_189
timestamp 1698175906
transform 1 0 22512 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_193
timestamp 1698175906
transform 1 0 22960 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_201
timestamp 1698175906
transform 1 0 23856 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_203
timestamp 1698175906
transform 1 0 24080 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_224
timestamp 1698175906
transform 1 0 26432 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_256
timestamp 1698175906
transform 1 0 30016 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_272
timestamp 1698175906
transform 1 0 31808 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_282
timestamp 1698175906
transform 1 0 32928 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_314
timestamp 1698175906
transform 1 0 36512 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_330
timestamp 1698175906
transform 1 0 38304 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_111
timestamp 1698175906
transform 1 0 13776 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_129
timestamp 1698175906
transform 1 0 15792 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_131
timestamp 1698175906
transform 1 0 16016 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_161
timestamp 1698175906
transform 1 0 19376 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_165
timestamp 1698175906
transform 1 0 19824 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_173
timestamp 1698175906
transform 1 0 20720 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_177
timestamp 1698175906
transform 1 0 21168 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_179
timestamp 1698175906
transform 1 0 21392 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_192
timestamp 1698175906
transform 1 0 22848 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_196
timestamp 1698175906
transform 1 0 23296 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_228
timestamp 1698175906
transform 1 0 26880 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_244
timestamp 1698175906
transform 1 0 28672 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_317
timestamp 1698175906
transform 1 0 36848 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_325
timestamp 1698175906
transform 1 0 37744 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_329
timestamp 1698175906
transform 1 0 38192 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_72
timestamp 1698175906
transform 1 0 9408 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_88
timestamp 1698175906
transform 1 0 11200 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_118
timestamp 1698175906
transform 1 0 14560 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_126
timestamp 1698175906
transform 1 0 15456 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_128
timestamp 1698175906
transform 1 0 15680 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_131
timestamp 1698175906
transform 1 0 16016 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_139
timestamp 1698175906
transform 1 0 16912 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_148
timestamp 1698175906
transform 1 0 17920 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_180
timestamp 1698175906
transform 1 0 21504 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_192
timestamp 1698175906
transform 1 0 22848 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_208
timestamp 1698175906
transform 1 0 24640 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_212
timestamp 1698175906
transform 1 0 25088 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_221
timestamp 1698175906
transform 1 0 26096 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_225
timestamp 1698175906
transform 1 0 26544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_256
timestamp 1698175906
transform 1 0 30016 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_272
timestamp 1698175906
transform 1 0 31808 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_282
timestamp 1698175906
transform 1 0 32928 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_314
timestamp 1698175906
transform 1 0 36512 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_330
timestamp 1698175906
transform 1 0 38304 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_37
timestamp 1698175906
transform 1 0 5488 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_53
timestamp 1698175906
transform 1 0 7280 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_57
timestamp 1698175906
transform 1 0 7728 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_87
timestamp 1698175906
transform 1 0 11088 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_91
timestamp 1698175906
transform 1 0 11536 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_99
timestamp 1698175906
transform 1 0 12432 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_103
timestamp 1698175906
transform 1 0 12880 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_107
timestamp 1698175906
transform 1 0 13328 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_115
timestamp 1698175906
transform 1 0 14224 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_117
timestamp 1698175906
transform 1 0 14448 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_120
timestamp 1698175906
transform 1 0 14784 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_124
timestamp 1698175906
transform 1 0 15232 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_126
timestamp 1698175906
transform 1 0 15456 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_156
timestamp 1698175906
transform 1 0 18816 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_172
timestamp 1698175906
transform 1 0 20608 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_174
timestamp 1698175906
transform 1 0 20832 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_177
timestamp 1698175906
transform 1 0 21168 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_193
timestamp 1698175906
transform 1 0 22960 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_201
timestamp 1698175906
transform 1 0 23856 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_205
timestamp 1698175906
transform 1 0 24304 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_236
timestamp 1698175906
transform 1 0 27776 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_240
timestamp 1698175906
transform 1 0 28224 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_244
timestamp 1698175906
transform 1 0 28672 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 29008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_317
timestamp 1698175906
transform 1 0 36848 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_325
timestamp 1698175906
transform 1 0 37744 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_72
timestamp 1698175906
transform 1 0 9408 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_104
timestamp 1698175906
transform 1 0 12992 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_120
timestamp 1698175906
transform 1 0 14784 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_128
timestamp 1698175906
transform 1 0 15680 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_130
timestamp 1698175906
transform 1 0 15904 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_135
timestamp 1698175906
transform 1 0 16464 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_139
timestamp 1698175906
transform 1 0 16912 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_142
timestamp 1698175906
transform 1 0 17248 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_158
timestamp 1698175906
transform 1 0 19040 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_162
timestamp 1698175906
transform 1 0 19488 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_168
timestamp 1698175906
transform 1 0 20160 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_200
timestamp 1698175906
transform 1 0 23744 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_208
timestamp 1698175906
transform 1 0 24640 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_240
timestamp 1698175906
transform 1 0 28224 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_244
timestamp 1698175906
transform 1 0 28672 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_248
timestamp 1698175906
transform 1 0 29120 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_282
timestamp 1698175906
transform 1 0 32928 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_314
timestamp 1698175906
transform 1 0 36512 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_330
timestamp 1698175906
transform 1 0 38304 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_34
timestamp 1698175906
transform 1 0 5152 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_37
timestamp 1698175906
transform 1 0 5488 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_45
timestamp 1698175906
transform 1 0 6384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_78
timestamp 1698175906
transform 1 0 10080 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_82
timestamp 1698175906
transform 1 0 10528 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_98
timestamp 1698175906
transform 1 0 12320 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_102
timestamp 1698175906
transform 1 0 12768 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_104
timestamp 1698175906
transform 1 0 12992 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_107
timestamp 1698175906
transform 1 0 13328 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_111
timestamp 1698175906
transform 1 0 13776 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_182
timestamp 1698175906
transform 1 0 21728 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_186
timestamp 1698175906
transform 1 0 22176 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_211
timestamp 1698175906
transform 1 0 24976 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_213
timestamp 1698175906
transform 1 0 25200 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 27776 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_240
timestamp 1698175906
transform 1 0 28224 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_244
timestamp 1698175906
transform 1 0 28672 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_247
timestamp 1698175906
transform 1 0 29008 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_249
timestamp 1698175906
transform 1 0 29232 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_279
timestamp 1698175906
transform 1 0 32592 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_287
timestamp 1698175906
transform 1 0 33488 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_317
timestamp 1698175906
transform 1 0 36848 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_325
timestamp 1698175906
transform 1 0 37744 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_329
timestamp 1698175906
transform 1 0 38192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_2
timestamp 1698175906
transform 1 0 1568 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_34
timestamp 1698175906
transform 1 0 5152 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_50
timestamp 1698175906
transform 1 0 6944 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_69
timestamp 1698175906
transform 1 0 9072 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_77
timestamp 1698175906
transform 1 0 9968 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_81
timestamp 1698175906
transform 1 0 10416 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_85
timestamp 1698175906
transform 1 0 10864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_92
timestamp 1698175906
transform 1 0 11648 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_96
timestamp 1698175906
transform 1 0 12096 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_98
timestamp 1698175906
transform 1 0 12320 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_130
timestamp 1698175906
transform 1 0 15904 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_138
timestamp 1698175906
transform 1 0 16800 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_165
timestamp 1698175906
transform 1 0 19824 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_167
timestamp 1698175906
transform 1 0 20048 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_216
timestamp 1698175906
transform 1 0 25536 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_225
timestamp 1698175906
transform 1 0 26544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_227
timestamp 1698175906
transform 1 0 26768 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_230
timestamp 1698175906
transform 1 0 27104 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_262
timestamp 1698175906
transform 1 0 30688 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_278
timestamp 1698175906
transform 1 0 32480 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_282
timestamp 1698175906
transform 1 0 32928 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_284
timestamp 1698175906
transform 1 0 33152 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_314
timestamp 1698175906
transform 1 0 36512 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_330
timestamp 1698175906
transform 1 0 38304 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_8
timestamp 1698175906
transform 1 0 2240 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_12
timestamp 1698175906
transform 1 0 2688 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_28
timestamp 1698175906
transform 1 0 4480 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_32
timestamp 1698175906
transform 1 0 4928 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_34
timestamp 1698175906
transform 1 0 5152 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_37
timestamp 1698175906
transform 1 0 5488 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_53
timestamp 1698175906
transform 1 0 7280 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_57
timestamp 1698175906
transform 1 0 7728 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_59
timestamp 1698175906
transform 1 0 7952 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_107
timestamp 1698175906
transform 1 0 13328 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_115
timestamp 1698175906
transform 1 0 14224 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_156
timestamp 1698175906
transform 1 0 18816 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_174
timestamp 1698175906
transform 1 0 20832 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_177
timestamp 1698175906
transform 1 0 21168 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_185
timestamp 1698175906
transform 1 0 22064 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_225
timestamp 1698175906
transform 1 0 26544 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_241
timestamp 1698175906
transform 1 0 28336 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_247
timestamp 1698175906
transform 1 0 29008 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_251
timestamp 1698175906
transform 1 0 29456 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_304
timestamp 1698175906
transform 1 0 35392 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_312
timestamp 1698175906
transform 1 0 36288 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_314
timestamp 1698175906
transform 1 0 36512 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_317
timestamp 1698175906
transform 1 0 36848 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_325
timestamp 1698175906
transform 1 0 37744 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_329
timestamp 1698175906
transform 1 0 38192 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_8
timestamp 1698175906
transform 1 0 2240 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_47_12
timestamp 1698175906
transform 1 0 2688 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_44
timestamp 1698175906
transform 1 0 6272 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_60
timestamp 1698175906
transform 1 0 8064 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_68
timestamp 1698175906
transform 1 0 8960 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_72
timestamp 1698175906
transform 1 0 9408 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_78
timestamp 1698175906
transform 1 0 10080 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_82
timestamp 1698175906
transform 1 0 10528 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_98
timestamp 1698175906
transform 1 0 12320 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_116
timestamp 1698175906
transform 1 0 14336 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_132
timestamp 1698175906
transform 1 0 16128 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_142
timestamp 1698175906
transform 1 0 17248 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_150
timestamp 1698175906
transform 1 0 18144 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_154
timestamp 1698175906
transform 1 0 18592 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_158
timestamp 1698175906
transform 1 0 19040 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_191
timestamp 1698175906
transform 1 0 22736 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_195
timestamp 1698175906
transform 1 0 23184 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_47_212
timestamp 1698175906
transform 1 0 25088 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_244
timestamp 1698175906
transform 1 0 28672 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_252
timestamp 1698175906
transform 1 0 29568 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_271
timestamp 1698175906
transform 1 0 31696 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_311
timestamp 1698175906
transform 1 0 36176 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_327
timestamp 1698175906
transform 1 0 37968 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_8
timestamp 1698175906
transform 1 0 2240 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_12
timestamp 1698175906
transform 1 0 2688 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_28
timestamp 1698175906
transform 1 0 4480 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_32
timestamp 1698175906
transform 1 0 4928 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_34
timestamp 1698175906
transform 1 0 5152 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_37
timestamp 1698175906
transform 1 0 5488 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_69
timestamp 1698175906
transform 1 0 9072 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_77
timestamp 1698175906
transform 1 0 9968 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_81
timestamp 1698175906
transform 1 0 10416 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_83
timestamp 1698175906
transform 1 0 10640 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_92
timestamp 1698175906
transform 1 0 11648 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_96
timestamp 1698175906
transform 1 0 12096 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_104
timestamp 1698175906
transform 1 0 12992 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_107
timestamp 1698175906
transform 1 0 13328 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_161
timestamp 1698175906
transform 1 0 19376 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_170
timestamp 1698175906
transform 1 0 20384 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_174
timestamp 1698175906
transform 1 0 20832 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_177
timestamp 1698175906
transform 1 0 21168 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_190
timestamp 1698175906
transform 1 0 22624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_200
timestamp 1698175906
transform 1 0 23744 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_239
timestamp 1698175906
transform 1 0 28112 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_276
timestamp 1698175906
transform 1 0 32256 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_317
timestamp 1698175906
transform 1 0 36848 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_325
timestamp 1698175906
transform 1 0 37744 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_329
timestamp 1698175906
transform 1 0 38192 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_2
timestamp 1698175906
transform 1 0 1568 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_34
timestamp 1698175906
transform 1 0 5152 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_50
timestamp 1698175906
transform 1 0 6944 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_58
timestamp 1698175906
transform 1 0 7840 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_64
timestamp 1698175906
transform 1 0 8512 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_68
timestamp 1698175906
transform 1 0 8960 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_72
timestamp 1698175906
transform 1 0 9408 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_104
timestamp 1698175906
transform 1 0 12992 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_112
timestamp 1698175906
transform 1 0 13888 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_116
timestamp 1698175906
transform 1 0 14336 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_118
timestamp 1698175906
transform 1 0 14560 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_123
timestamp 1698175906
transform 1 0 15120 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_138
timestamp 1698175906
transform 1 0 16800 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_142
timestamp 1698175906
transform 1 0 17248 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_146
timestamp 1698175906
transform 1 0 17696 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_158
timestamp 1698175906
transform 1 0 19040 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_172
timestamp 1698175906
transform 1 0 20608 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_188
timestamp 1698175906
transform 1 0 22400 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_194
timestamp 1698175906
transform 1 0 23072 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_226
timestamp 1698175906
transform 1 0 26656 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_234
timestamp 1698175906
transform 1 0 27552 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_279
timestamp 1698175906
transform 1 0 32592 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_290
timestamp 1698175906
transform 1 0 33824 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_301
timestamp 1698175906
transform 1 0 35056 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_2
timestamp 1698175906
transform 1 0 1568 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_34
timestamp 1698175906
transform 1 0 5152 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_37
timestamp 1698175906
transform 1 0 5488 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_45
timestamp 1698175906
transform 1 0 6384 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_86
timestamp 1698175906
transform 1 0 10976 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_90
timestamp 1698175906
transform 1 0 11424 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_98
timestamp 1698175906
transform 1 0 12320 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_102
timestamp 1698175906
transform 1 0 12768 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_104
timestamp 1698175906
transform 1 0 12992 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_127
timestamp 1698175906
transform 1 0 15568 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_129
timestamp 1698175906
transform 1 0 15792 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_162
timestamp 1698175906
transform 1 0 19488 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_164
timestamp 1698175906
transform 1 0 19712 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_182
timestamp 1698175906
transform 1 0 21728 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_198
timestamp 1698175906
transform 1 0 23520 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_206
timestamp 1698175906
transform 1 0 24416 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_210
timestamp 1698175906
transform 1 0 24864 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_225
timestamp 1698175906
transform 1 0 26544 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_229
timestamp 1698175906
transform 1 0 26992 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_237
timestamp 1698175906
transform 1 0 27888 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_239
timestamp 1698175906
transform 1 0 28112 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_247
timestamp 1698175906
transform 1 0 29008 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_317
timestamp 1698175906
transform 1 0 36848 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_325
timestamp 1698175906
transform 1 0 37744 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_329
timestamp 1698175906
transform 1 0 38192 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_2
timestamp 1698175906
transform 1 0 1568 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_18
timestamp 1698175906
transform 1 0 3360 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_26
timestamp 1698175906
transform 1 0 4256 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_30
timestamp 1698175906
transform 1 0 4704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_32
timestamp 1698175906
transform 1 0 4928 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_64
timestamp 1698175906
transform 1 0 8512 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_68
timestamp 1698175906
transform 1 0 8960 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_72
timestamp 1698175906
transform 1 0 9408 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_74
timestamp 1698175906
transform 1 0 9632 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_83
timestamp 1698175906
transform 1 0 10640 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_142
timestamp 1698175906
transform 1 0 17248 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_169
timestamp 1698175906
transform 1 0 20272 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_173
timestamp 1698175906
transform 1 0 20720 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_175
timestamp 1698175906
transform 1 0 20944 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_189
timestamp 1698175906
transform 1 0 22512 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_193
timestamp 1698175906
transform 1 0 22960 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_208
timestamp 1698175906
transform 1 0 24640 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_212
timestamp 1698175906
transform 1 0 25088 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_214
timestamp 1698175906
transform 1 0 25312 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_246
timestamp 1698175906
transform 1 0 28896 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_250
timestamp 1698175906
transform 1 0 29344 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_264
timestamp 1698175906
transform 1 0 30912 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_266
timestamp 1698175906
transform 1 0 31136 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_298
timestamp 1698175906
transform 1 0 34720 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_8
timestamp 1698175906
transform 1 0 2240 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_12
timestamp 1698175906
transform 1 0 2688 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_28
timestamp 1698175906
transform 1 0 4480 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_32
timestamp 1698175906
transform 1 0 4928 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_34
timestamp 1698175906
transform 1 0 5152 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_37
timestamp 1698175906
transform 1 0 5488 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_45
timestamp 1698175906
transform 1 0 6384 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_51
timestamp 1698175906
transform 1 0 7056 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_53
timestamp 1698175906
transform 1 0 7280 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_59
timestamp 1698175906
transform 1 0 7952 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_68
timestamp 1698175906
transform 1 0 8960 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_107
timestamp 1698175906
transform 1 0 13328 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_189
timestamp 1698175906
transform 1 0 22512 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_193
timestamp 1698175906
transform 1 0 22960 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_226
timestamp 1698175906
transform 1 0 26656 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_242
timestamp 1698175906
transform 1 0 28448 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_244
timestamp 1698175906
transform 1 0 28672 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_247
timestamp 1698175906
transform 1 0 29008 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_255
timestamp 1698175906
transform 1 0 29904 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_259
timestamp 1698175906
transform 1 0 30352 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_313
timestamp 1698175906
transform 1 0 36400 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_317
timestamp 1698175906
transform 1 0 36848 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_325
timestamp 1698175906
transform 1 0 37744 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_329
timestamp 1698175906
transform 1 0 38192 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_8
timestamp 1698175906
transform 1 0 2240 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_53_12
timestamp 1698175906
transform 1 0 2688 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_44
timestamp 1698175906
transform 1 0 6272 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_46
timestamp 1698175906
transform 1 0 6496 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_52
timestamp 1698175906
transform 1 0 7168 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_72
timestamp 1698175906
transform 1 0 9408 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_74
timestamp 1698175906
transform 1 0 9632 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_81
timestamp 1698175906
transform 1 0 10416 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_87
timestamp 1698175906
transform 1 0 11088 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_103
timestamp 1698175906
transform 1 0 12880 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_142
timestamp 1698175906
transform 1 0 17248 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_158
timestamp 1698175906
transform 1 0 19040 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_162
timestamp 1698175906
transform 1 0 19488 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_171
timestamp 1698175906
transform 1 0 20496 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_187
timestamp 1698175906
transform 1 0 22288 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_197
timestamp 1698175906
transform 1 0 23408 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_205
timestamp 1698175906
transform 1 0 24304 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_209
timestamp 1698175906
transform 1 0 24752 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_212
timestamp 1698175906
transform 1 0 25088 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_224
timestamp 1698175906
transform 1 0 26432 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_240
timestamp 1698175906
transform 1 0 28224 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_244
timestamp 1698175906
transform 1 0 28672 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_246
timestamp 1698175906
transform 1 0 28896 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_265
timestamp 1698175906
transform 1 0 31024 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_269
timestamp 1698175906
transform 1 0 31472 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_301
timestamp 1698175906
transform 1 0 35056 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_2
timestamp 1698175906
transform 1 0 1568 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_34
timestamp 1698175906
transform 1 0 5152 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_37
timestamp 1698175906
transform 1 0 5488 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_74
timestamp 1698175906
transform 1 0 9632 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_107
timestamp 1698175906
transform 1 0 13328 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_142
timestamp 1698175906
transform 1 0 17248 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_174
timestamp 1698175906
transform 1 0 20832 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_177
timestamp 1698175906
transform 1 0 21168 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_205
timestamp 1698175906
transform 1 0 24304 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_220
timestamp 1698175906
transform 1 0 25984 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_236
timestamp 1698175906
transform 1 0 27776 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_244
timestamp 1698175906
transform 1 0 28672 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_262
timestamp 1698175906
transform 1 0 30688 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_282
timestamp 1698175906
transform 1 0 32928 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_317
timestamp 1698175906
transform 1 0 36848 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_325
timestamp 1698175906
transform 1 0 37744 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_329
timestamp 1698175906
transform 1 0 38192 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_55_2
timestamp 1698175906
transform 1 0 1568 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_34
timestamp 1698175906
transform 1 0 5152 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_50
timestamp 1698175906
transform 1 0 6944 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_58
timestamp 1698175906
transform 1 0 7840 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_77
timestamp 1698175906
transform 1 0 9968 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_86
timestamp 1698175906
transform 1 0 10976 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_55_90
timestamp 1698175906
transform 1 0 11424 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_122
timestamp 1698175906
transform 1 0 15008 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_132
timestamp 1698175906
transform 1 0 16128 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_150
timestamp 1698175906
transform 1 0 18144 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_154
timestamp 1698175906
transform 1 0 18592 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_169
timestamp 1698175906
transform 1 0 20272 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_177
timestamp 1698175906
transform 1 0 21168 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_179
timestamp 1698175906
transform 1 0 21392 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_190
timestamp 1698175906
transform 1 0 22624 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_206
timestamp 1698175906
transform 1 0 24416 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_241
timestamp 1698175906
transform 1 0 28336 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_257
timestamp 1698175906
transform 1 0 30128 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_2
timestamp 1698175906
transform 1 0 1568 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_34
timestamp 1698175906
transform 1 0 5152 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_37
timestamp 1698175906
transform 1 0 5488 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_53
timestamp 1698175906
transform 1 0 7280 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_57
timestamp 1698175906
transform 1 0 7728 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_63
timestamp 1698175906
transform 1 0 8400 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_67
timestamp 1698175906
transform 1 0 8848 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_69
timestamp 1698175906
transform 1 0 9072 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_72
timestamp 1698175906
transform 1 0 9408 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_104
timestamp 1698175906
transform 1 0 12992 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_107
timestamp 1698175906
transform 1 0 13328 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_139
timestamp 1698175906
transform 1 0 16912 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_154
timestamp 1698175906
transform 1 0 18592 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_162
timestamp 1698175906
transform 1 0 19488 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_166
timestamp 1698175906
transform 1 0 19936 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_168
timestamp 1698175906
transform 1 0 20160 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_177
timestamp 1698175906
transform 1 0 21168 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_209
timestamp 1698175906
transform 1 0 24752 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_212
timestamp 1698175906
transform 1 0 25088 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_216
timestamp 1698175906
transform 1 0 25536 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_226
timestamp 1698175906
transform 1 0 26656 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_232
timestamp 1698175906
transform 1 0 27328 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_240
timestamp 1698175906
transform 1 0 28224 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_244
timestamp 1698175906
transform 1 0 28672 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_247
timestamp 1698175906
transform 1 0 29008 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_251
timestamp 1698175906
transform 1 0 29456 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_253
timestamp 1698175906
transform 1 0 29680 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_309
timestamp 1698175906
transform 1 0 35952 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_313
timestamp 1698175906
transform 1 0 36400 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_317
timestamp 1698175906
transform 1 0 36848 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_325
timestamp 1698175906
transform 1 0 37744 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_329
timestamp 1698175906
transform 1 0 38192 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_8
timestamp 1698175906
transform 1 0 2240 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_57_12
timestamp 1698175906
transform 1 0 2688 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_44
timestamp 1698175906
transform 1 0 6272 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_46
timestamp 1698175906
transform 1 0 6496 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_58
timestamp 1698175906
transform 1 0 7840 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_66
timestamp 1698175906
transform 1 0 8736 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_72
timestamp 1698175906
transform 1 0 9408 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_80
timestamp 1698175906
transform 1 0 10304 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_84
timestamp 1698175906
transform 1 0 10752 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_57_96
timestamp 1698175906
transform 1 0 12096 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_128
timestamp 1698175906
transform 1 0 15680 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_136
timestamp 1698175906
transform 1 0 16576 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_142
timestamp 1698175906
transform 1 0 17248 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_146
timestamp 1698175906
transform 1 0 17696 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_148
timestamp 1698175906
transform 1 0 17920 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_158
timestamp 1698175906
transform 1 0 19040 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_166
timestamp 1698175906
transform 1 0 19936 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_198
timestamp 1698175906
transform 1 0 23520 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_218
timestamp 1698175906
transform 1 0 25760 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_240
timestamp 1698175906
transform 1 0 28224 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_256
timestamp 1698175906
transform 1 0 30016 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_279
timestamp 1698175906
transform 1 0 32592 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_304
timestamp 1698175906
transform 1 0 35392 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_8
timestamp 1698175906
transform 1 0 2240 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_12
timestamp 1698175906
transform 1 0 2688 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_28
timestamp 1698175906
transform 1 0 4480 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_32
timestamp 1698175906
transform 1 0 4928 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_34
timestamp 1698175906
transform 1 0 5152 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_37
timestamp 1698175906
transform 1 0 5488 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_45
timestamp 1698175906
transform 1 0 6384 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_56
timestamp 1698175906
transform 1 0 7616 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_60
timestamp 1698175906
transform 1 0 8064 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_69
timestamp 1698175906
transform 1 0 9072 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_73
timestamp 1698175906
transform 1 0 9520 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_75
timestamp 1698175906
transform 1 0 9744 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_78
timestamp 1698175906
transform 1 0 10080 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_94
timestamp 1698175906
transform 1 0 11872 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_102
timestamp 1698175906
transform 1 0 12768 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_104
timestamp 1698175906
transform 1 0 12992 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_107
timestamp 1698175906
transform 1 0 13328 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_123
timestamp 1698175906
transform 1 0 15120 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_136
timestamp 1698175906
transform 1 0 16576 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_168
timestamp 1698175906
transform 1 0 20160 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_172
timestamp 1698175906
transform 1 0 20608 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_174
timestamp 1698175906
transform 1 0 20832 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_177
timestamp 1698175906
transform 1 0 21168 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_202
timestamp 1698175906
transform 1 0 23968 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_232
timestamp 1698175906
transform 1 0 27328 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_240
timestamp 1698175906
transform 1 0 28224 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_244
timestamp 1698175906
transform 1 0 28672 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_292
timestamp 1698175906
transform 1 0 34048 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_312
timestamp 1698175906
transform 1 0 36288 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_314
timestamp 1698175906
transform 1 0 36512 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_317
timestamp 1698175906
transform 1 0 36848 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_325
timestamp 1698175906
transform 1 0 37744 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_329
timestamp 1698175906
transform 1 0 38192 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_8
timestamp 1698175906
transform 1 0 2240 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_12
timestamp 1698175906
transform 1 0 2688 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_16
timestamp 1698175906
transform 1 0 3136 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_32
timestamp 1698175906
transform 1 0 4928 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_64
timestamp 1698175906
transform 1 0 8512 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_68
timestamp 1698175906
transform 1 0 8960 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_77
timestamp 1698175906
transform 1 0 9968 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_84
timestamp 1698175906
transform 1 0 10752 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_86
timestamp 1698175906
transform 1 0 10976 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_135
timestamp 1698175906
transform 1 0 16464 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_139
timestamp 1698175906
transform 1 0 16912 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_142
timestamp 1698175906
transform 1 0 17248 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_144
timestamp 1698175906
transform 1 0 17472 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_160
timestamp 1698175906
transform 1 0 19264 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_168
timestamp 1698175906
transform 1 0 20160 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_172
timestamp 1698175906
transform 1 0 20608 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_205
timestamp 1698175906
transform 1 0 24304 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_209
timestamp 1698175906
transform 1 0 24752 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_212
timestamp 1698175906
transform 1 0 25088 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_228
timestamp 1698175906
transform 1 0 26880 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_236
timestamp 1698175906
transform 1 0 27776 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_269
timestamp 1698175906
transform 1 0 31472 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_277
timestamp 1698175906
transform 1 0 32368 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_279
timestamp 1698175906
transform 1 0 32592 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_282
timestamp 1698175906
transform 1 0 32928 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_327
timestamp 1698175906
transform 1 0 37968 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_14
timestamp 1698175906
transform 1 0 2912 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_18
timestamp 1698175906
transform 1 0 3360 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_34
timestamp 1698175906
transform 1 0 5152 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_37
timestamp 1698175906
transform 1 0 5488 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_53
timestamp 1698175906
transform 1 0 7280 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_59
timestamp 1698175906
transform 1 0 7952 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_67
timestamp 1698175906
transform 1 0 8848 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_85
timestamp 1698175906
transform 1 0 10864 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_107
timestamp 1698175906
transform 1 0 13328 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_115
timestamp 1698175906
transform 1 0 14224 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_119
timestamp 1698175906
transform 1 0 14672 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_121
timestamp 1698175906
transform 1 0 14896 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_126
timestamp 1698175906
transform 1 0 15456 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_154
timestamp 1698175906
transform 1 0 18592 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_227
timestamp 1698175906
transform 1 0 26768 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_231
timestamp 1698175906
transform 1 0 27216 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_239
timestamp 1698175906
transform 1 0 28112 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_243
timestamp 1698175906
transform 1 0 28560 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_60_247
timestamp 1698175906
transform 1 0 29008 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_279
timestamp 1698175906
transform 1 0 32592 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_289
timestamp 1698175906
transform 1 0 33712 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_305
timestamp 1698175906
transform 1 0 35504 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_313
timestamp 1698175906
transform 1 0 36400 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_317
timestamp 1698175906
transform 1 0 36848 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_325
timestamp 1698175906
transform 1 0 37744 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_329
timestamp 1698175906
transform 1 0 38192 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_8
timestamp 1698175906
transform 1 0 2240 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_12
timestamp 1698175906
transform 1 0 2688 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_28
timestamp 1698175906
transform 1 0 4480 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_36
timestamp 1698175906
transform 1 0 5376 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_40
timestamp 1698175906
transform 1 0 5824 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_84
timestamp 1698175906
transform 1 0 10752 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_88
timestamp 1698175906
transform 1 0 11200 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_90
timestamp 1698175906
transform 1 0 11424 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_120
timestamp 1698175906
transform 1 0 14784 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_124
timestamp 1698175906
transform 1 0 15232 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_138
timestamp 1698175906
transform 1 0 16800 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_174
timestamp 1698175906
transform 1 0 20832 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_182
timestamp 1698175906
transform 1 0 21728 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_206
timestamp 1698175906
transform 1 0 24416 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_212
timestamp 1698175906
transform 1 0 25088 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_230
timestamp 1698175906
transform 1 0 27104 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_234
timestamp 1698175906
transform 1 0 27552 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_238
timestamp 1698175906
transform 1 0 28000 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_270
timestamp 1698175906
transform 1 0 31584 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_278
timestamp 1698175906
transform 1 0 32480 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_282
timestamp 1698175906
transform 1 0 32928 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_298
timestamp 1698175906
transform 1 0 34720 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_302
timestamp 1698175906
transform 1 0 35168 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_304
timestamp 1698175906
transform 1 0 35392 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_8
timestamp 1698175906
transform 1 0 2240 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_12
timestamp 1698175906
transform 1 0 2688 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_28
timestamp 1698175906
transform 1 0 4480 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_32
timestamp 1698175906
transform 1 0 4928 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_34
timestamp 1698175906
transform 1 0 5152 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_62_37
timestamp 1698175906
transform 1 0 5488 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_69
timestamp 1698175906
transform 1 0 9072 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_85
timestamp 1698175906
transform 1 0 10864 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_107
timestamp 1698175906
transform 1 0 13328 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_115
timestamp 1698175906
transform 1 0 14224 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_119
timestamp 1698175906
transform 1 0 14672 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_171
timestamp 1698175906
transform 1 0 20496 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_177
timestamp 1698175906
transform 1 0 21168 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_181
timestamp 1698175906
transform 1 0 21616 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_219
timestamp 1698175906
transform 1 0 25872 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_223
timestamp 1698175906
transform 1 0 26320 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_232
timestamp 1698175906
transform 1 0 27328 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_236
timestamp 1698175906
transform 1 0 27776 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_244
timestamp 1698175906
transform 1 0 28672 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_62_247
timestamp 1698175906
transform 1 0 29008 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_279
timestamp 1698175906
transform 1 0 32592 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_287
timestamp 1698175906
transform 1 0 33488 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_294
timestamp 1698175906
transform 1 0 34272 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_310
timestamp 1698175906
transform 1 0 36064 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_314
timestamp 1698175906
transform 1 0 36512 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_317
timestamp 1698175906
transform 1 0 36848 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_325
timestamp 1698175906
transform 1 0 37744 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_329
timestamp 1698175906
transform 1 0 38192 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_2
timestamp 1698175906
transform 1 0 1568 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_66
timestamp 1698175906
transform 1 0 8736 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_72
timestamp 1698175906
transform 1 0 9408 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_76
timestamp 1698175906
transform 1 0 9856 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_63_82
timestamp 1698175906
transform 1 0 10528 0 -1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_114
timestamp 1698175906
transform 1 0 14112 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_118
timestamp 1698175906
transform 1 0 14560 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_158
timestamp 1698175906
transform 1 0 19040 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_195
timestamp 1698175906
transform 1 0 23184 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_199
timestamp 1698175906
transform 1 0 23632 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_212
timestamp 1698175906
transform 1 0 25088 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_216
timestamp 1698175906
transform 1 0 25536 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_63_246
timestamp 1698175906
transform 1 0 28896 0 -1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_278
timestamp 1698175906
transform 1 0 32480 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_311
timestamp 1698175906
transform 1 0 36176 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_327
timestamp 1698175906
transform 1 0 37968 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_8
timestamp 1698175906
transform 1 0 2240 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_12
timestamp 1698175906
transform 1 0 2688 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_28
timestamp 1698175906
transform 1 0 4480 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_32
timestamp 1698175906
transform 1 0 4928 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_34
timestamp 1698175906
transform 1 0 5152 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_37
timestamp 1698175906
transform 1 0 5488 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_101
timestamp 1698175906
transform 1 0 12656 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_107
timestamp 1698175906
transform 1 0 13328 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_115
timestamp 1698175906
transform 1 0 14224 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_119
timestamp 1698175906
transform 1 0 14672 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_121
timestamp 1698175906
transform 1 0 14896 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_166
timestamp 1698175906
transform 1 0 19936 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_174
timestamp 1698175906
transform 1 0 20832 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_185
timestamp 1698175906
transform 1 0 22064 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_236
timestamp 1698175906
transform 1 0 27776 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_244
timestamp 1698175906
transform 1 0 28672 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_247
timestamp 1698175906
transform 1 0 29008 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_311
timestamp 1698175906
transform 1 0 36176 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_317
timestamp 1698175906
transform 1 0 36848 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_325
timestamp 1698175906
transform 1 0 37744 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_329
timestamp 1698175906
transform 1 0 38192 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_65_2
timestamp 1698175906
transform 1 0 1568 0 -1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_34
timestamp 1698175906
transform 1 0 5152 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_50
timestamp 1698175906
transform 1 0 6944 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_54
timestamp 1698175906
transform 1 0 7392 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_61
timestamp 1698175906
transform 1 0 8176 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_72
timestamp 1698175906
transform 1 0 9408 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_80
timestamp 1698175906
transform 1 0 10304 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_88
timestamp 1698175906
transform 1 0 11200 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_92
timestamp 1698175906
transform 1 0 11648 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_138
timestamp 1698175906
transform 1 0 16800 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_65_175
timestamp 1698175906
transform 1 0 20944 0 -1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_207
timestamp 1698175906
transform 1 0 24528 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_209
timestamp 1698175906
transform 1 0 24752 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_218
timestamp 1698175906
transform 1 0 25760 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_226
timestamp 1698175906
transform 1 0 26656 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_257
timestamp 1698175906
transform 1 0 30128 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_273
timestamp 1698175906
transform 1 0 31920 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_277
timestamp 1698175906
transform 1 0 32368 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_279
timestamp 1698175906
transform 1 0 32592 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_282
timestamp 1698175906
transform 1 0 32928 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_298
timestamp 1698175906
transform 1 0 34720 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_302
timestamp 1698175906
transform 1 0 35168 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_304
timestamp 1698175906
transform 1 0 35392 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_8
timestamp 1698175906
transform 1 0 2240 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_12
timestamp 1698175906
transform 1 0 2688 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_28
timestamp 1698175906
transform 1 0 4480 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_32
timestamp 1698175906
transform 1 0 4928 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_34
timestamp 1698175906
transform 1 0 5152 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_37
timestamp 1698175906
transform 1 0 5488 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_41
timestamp 1698175906
transform 1 0 5936 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_76
timestamp 1698175906
transform 1 0 9856 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_78
timestamp 1698175906
transform 1 0 10080 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_107
timestamp 1698175906
transform 1 0 13328 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_115
timestamp 1698175906
transform 1 0 14224 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_119
timestamp 1698175906
transform 1 0 14672 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_162
timestamp 1698175906
transform 1 0 19488 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_170
timestamp 1698175906
transform 1 0 20384 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_174
timestamp 1698175906
transform 1 0 20832 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_177
timestamp 1698175906
transform 1 0 21168 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_179
timestamp 1698175906
transform 1 0 21392 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_193
timestamp 1698175906
transform 1 0 22960 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_201
timestamp 1698175906
transform 1 0 23856 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_205
timestamp 1698175906
transform 1 0 24304 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_207
timestamp 1698175906
transform 1 0 24528 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_255
timestamp 1698175906
transform 1 0 29904 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_287
timestamp 1698175906
transform 1 0 33488 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_303
timestamp 1698175906
transform 1 0 35280 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_311
timestamp 1698175906
transform 1 0 36176 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_317
timestamp 1698175906
transform 1 0 36848 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_325
timestamp 1698175906
transform 1 0 37744 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_329
timestamp 1698175906
transform 1 0 38192 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_8
timestamp 1698175906
transform 1 0 2240 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_12
timestamp 1698175906
transform 1 0 2688 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_28
timestamp 1698175906
transform 1 0 4480 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_36
timestamp 1698175906
transform 1 0 5376 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_38
timestamp 1698175906
transform 1 0 5600 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_80
timestamp 1698175906
transform 1 0 10304 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_88
timestamp 1698175906
transform 1 0 11200 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_159
timestamp 1698175906
transform 1 0 19152 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_187
timestamp 1698175906
transform 1 0 22288 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_203
timestamp 1698175906
transform 1 0 24080 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_212
timestamp 1698175906
transform 1 0 25088 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_221
timestamp 1698175906
transform 1 0 26096 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_225
timestamp 1698175906
transform 1 0 26544 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_227
timestamp 1698175906
transform 1 0 26768 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_257
timestamp 1698175906
transform 1 0 30128 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_273
timestamp 1698175906
transform 1 0 31920 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_277
timestamp 1698175906
transform 1 0 32368 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_279
timestamp 1698175906
transform 1 0 32592 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_282
timestamp 1698175906
transform 1 0 32928 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_314
timestamp 1698175906
transform 1 0 36512 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_330
timestamp 1698175906
transform 1 0 38304 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_8
timestamp 1698175906
transform 1 0 2240 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_68_12
timestamp 1698175906
transform 1 0 2688 0 1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_28
timestamp 1698175906
transform 1 0 4480 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_32
timestamp 1698175906
transform 1 0 4928 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_34
timestamp 1698175906
transform 1 0 5152 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_68_37
timestamp 1698175906
transform 1 0 5488 0 1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_68_66
timestamp 1698175906
transform 1 0 8736 0 1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_68_82
timestamp 1698175906
transform 1 0 10528 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_90
timestamp 1698175906
transform 1 0 11424 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_100
timestamp 1698175906
transform 1 0 12544 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_104
timestamp 1698175906
transform 1 0 12992 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_68_117
timestamp 1698175906
transform 1 0 14448 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_129
timestamp 1698175906
transform 1 0 15792 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_131
timestamp 1698175906
transform 1 0 16016 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_147
timestamp 1698175906
transform 1 0 17808 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_68_151
timestamp 1698175906
transform 1 0 18256 0 1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_68_167
timestamp 1698175906
transform 1 0 20048 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_219
timestamp 1698175906
transform 1 0 25872 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_244
timestamp 1698175906
transform 1 0 28672 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_68_247
timestamp 1698175906
transform 1 0 29008 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_311
timestamp 1698175906
transform 1 0 36176 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_68_317
timestamp 1698175906
transform 1 0 36848 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_325
timestamp 1698175906
transform 1 0 37744 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_329
timestamp 1698175906
transform 1 0 38192 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_8
timestamp 1698175906
transform 1 0 2240 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_69_12
timestamp 1698175906
transform 1 0 2688 0 -1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_69_44
timestamp 1698175906
transform 1 0 6272 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_52
timestamp 1698175906
transform 1 0 7168 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_69_61
timestamp 1698175906
transform 1 0 8176 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_69
timestamp 1698175906
transform 1 0 9072 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_72
timestamp 1698175906
transform 1 0 9408 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_74
timestamp 1698175906
transform 1 0 9632 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_69_81
timestamp 1698175906
transform 1 0 10416 0 -1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_97
timestamp 1698175906
transform 1 0 12208 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_101
timestamp 1698175906
transform 1 0 12656 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_69_109
timestamp 1698175906
transform 1 0 13552 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_69_158
timestamp 1698175906
transform 1 0 19040 0 -1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_174
timestamp 1698175906
transform 1 0 20832 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_178
timestamp 1698175906
transform 1 0 21280 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_208
timestamp 1698175906
transform 1 0 24640 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_212
timestamp 1698175906
transform 1 0 25088 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_216
timestamp 1698175906
transform 1 0 25536 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_69_269
timestamp 1698175906
transform 1 0 31472 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_277
timestamp 1698175906
transform 1 0 32368 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_279
timestamp 1698175906
transform 1 0 32592 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_69_282
timestamp 1698175906
transform 1 0 32928 0 -1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_69_314
timestamp 1698175906
transform 1 0 36512 0 -1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_330
timestamp 1698175906
transform 1 0 38304 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_8
timestamp 1698175906
transform 1 0 2240 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_70_12
timestamp 1698175906
transform 1 0 2688 0 1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_28
timestamp 1698175906
transform 1 0 4480 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_32
timestamp 1698175906
transform 1 0 4928 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_34
timestamp 1698175906
transform 1 0 5152 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_70_37
timestamp 1698175906
transform 1 0 5488 0 1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_69
timestamp 1698175906
transform 1 0 9072 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_73
timestamp 1698175906
transform 1 0 9520 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_70_82
timestamp 1698175906
transform 1 0 10528 0 1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_98
timestamp 1698175906
transform 1 0 12320 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_102
timestamp 1698175906
transform 1 0 12768 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_104
timestamp 1698175906
transform 1 0 12992 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70_117
timestamp 1698175906
transform 1 0 14448 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_125
timestamp 1698175906
transform 1 0 15344 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_129
timestamp 1698175906
transform 1 0 15792 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_139
timestamp 1698175906
transform 1 0 16912 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_155
timestamp 1698175906
transform 1 0 18704 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_70_159
timestamp 1698175906
transform 1 0 19152 0 1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_70_177
timestamp 1698175906
transform 1 0 21168 0 1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70_193
timestamp 1698175906
transform 1 0 22960 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_201
timestamp 1698175906
transform 1 0 23856 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_205
timestamp 1698175906
transform 1 0 24304 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_207
timestamp 1698175906
transform 1 0 24528 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_222
timestamp 1698175906
transform 1 0 26208 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_226
timestamp 1698175906
transform 1 0 26656 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70_236
timestamp 1698175906
transform 1 0 27776 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_244
timestamp 1698175906
transform 1 0 28672 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_247
timestamp 1698175906
transform 1 0 29008 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_311
timestamp 1698175906
transform 1 0 36176 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70_317
timestamp 1698175906
transform 1 0 36848 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_325
timestamp 1698175906
transform 1 0 37744 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_329
timestamp 1698175906
transform 1 0 38192 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_71_2
timestamp 1698175906
transform 1 0 1568 0 -1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_71_34
timestamp 1698175906
transform 1 0 5152 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_50
timestamp 1698175906
transform 1 0 6944 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_54
timestamp 1698175906
transform 1 0 7392 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_56
timestamp 1698175906
transform 1 0 7616 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_65
timestamp 1698175906
transform 1 0 8624 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_69
timestamp 1698175906
transform 1 0 9072 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_71_77
timestamp 1698175906
transform 1 0 9968 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_85
timestamp 1698175906
transform 1 0 10864 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_92
timestamp 1698175906
transform 1 0 11648 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_94
timestamp 1698175906
transform 1 0 11872 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_71_124
timestamp 1698175906
transform 1 0 15232 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_71_158
timestamp 1698175906
transform 1 0 19040 0 -1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_71_190
timestamp 1698175906
transform 1 0 22624 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_206
timestamp 1698175906
transform 1 0 24416 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_212
timestamp 1698175906
transform 1 0 25088 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_216
timestamp 1698175906
transform 1 0 25536 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_218
timestamp 1698175906
transform 1 0 25760 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_71_221
timestamp 1698175906
transform 1 0 26096 0 -1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_71_253
timestamp 1698175906
transform 1 0 29680 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_71_269
timestamp 1698175906
transform 1 0 31472 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_277
timestamp 1698175906
transform 1 0 32368 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_279
timestamp 1698175906
transform 1 0 32592 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_71_282
timestamp 1698175906
transform 1 0 32928 0 -1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_71_314
timestamp 1698175906
transform 1 0 36512 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_330
timestamp 1698175906
transform 1 0 38304 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_8
timestamp 1698175906
transform 1 0 2240 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_72_12
timestamp 1698175906
transform 1 0 2688 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_28
timestamp 1698175906
transform 1 0 4480 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_32
timestamp 1698175906
transform 1 0 4928 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_34
timestamp 1698175906
transform 1 0 5152 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_37
timestamp 1698175906
transform 1 0 5488 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_39
timestamp 1698175906
transform 1 0 5712 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_72_71
timestamp 1698175906
transform 1 0 9296 0 1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_103
timestamp 1698175906
transform 1 0 12880 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_113
timestamp 1698175906
transform 1 0 14000 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_72_167
timestamp 1698175906
transform 1 0 20048 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_72_177
timestamp 1698175906
transform 1 0 21168 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_72_193
timestamp 1698175906
transform 1 0 22960 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_201
timestamp 1698175906
transform 1 0 23856 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_205
timestamp 1698175906
transform 1 0 24304 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_219
timestamp 1698175906
transform 1 0 25872 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_72_227
timestamp 1698175906
transform 1 0 26768 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_243
timestamp 1698175906
transform 1 0 28560 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_72_247
timestamp 1698175906
transform 1 0 29008 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_311
timestamp 1698175906
transform 1 0 36176 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_72_317
timestamp 1698175906
transform 1 0 36848 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_325
timestamp 1698175906
transform 1 0 37744 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_329
timestamp 1698175906
transform 1 0 38192 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_2
timestamp 1698175906
transform 1 0 1568 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_66
timestamp 1698175906
transform 1 0 8736 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_73_72
timestamp 1698175906
transform 1 0 9408 0 -1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_88
timestamp 1698175906
transform 1 0 11200 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_142
timestamp 1698175906
transform 1 0 17248 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_169
timestamp 1698175906
transform 1 0 20272 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_73_193
timestamp 1698175906
transform 1 0 22960 0 -1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_209
timestamp 1698175906
transform 1 0 24752 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_212
timestamp 1698175906
transform 1 0 25088 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_73_245
timestamp 1698175906
transform 1 0 28784 0 -1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_277
timestamp 1698175906
transform 1 0 32368 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_279
timestamp 1698175906
transform 1 0 32592 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_73_282
timestamp 1698175906
transform 1 0 32928 0 -1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_73_314
timestamp 1698175906
transform 1 0 36512 0 -1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_330
timestamp 1698175906
transform 1 0 38304 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_74_2
timestamp 1698175906
transform 1 0 1568 0 1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_34
timestamp 1698175906
transform 1 0 5152 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_74_37
timestamp 1698175906
transform 1 0 5488 0 1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_74_53
timestamp 1698175906
transform 1 0 7280 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_75
timestamp 1698175906
transform 1 0 9744 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_77
timestamp 1698175906
transform 1 0 9968 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_74_83
timestamp 1698175906
transform 1 0 10640 0 1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_99
timestamp 1698175906
transform 1 0 12432 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_103
timestamp 1698175906
transform 1 0 12880 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_74_113
timestamp 1698175906
transform 1 0 14000 0 1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_74_145
timestamp 1698175906
transform 1 0 17584 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_153
timestamp 1698175906
transform 1 0 18480 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_74_177
timestamp 1698175906
transform 1 0 21168 0 1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_193
timestamp 1698175906
transform 1 0 22960 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_198
timestamp 1698175906
transform 1 0 23520 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_244
timestamp 1698175906
transform 1 0 28672 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_74_247
timestamp 1698175906
transform 1 0 29008 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_311
timestamp 1698175906
transform 1 0 36176 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_74_317
timestamp 1698175906
transform 1 0 36848 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_325
timestamp 1698175906
transform 1 0 37744 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_329
timestamp 1698175906
transform 1 0 38192 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_75_2
timestamp 1698175906
transform 1 0 1568 0 -1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_75_34
timestamp 1698175906
transform 1 0 5152 0 -1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_50
timestamp 1698175906
transform 1 0 6944 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_54
timestamp 1698175906
transform 1 0 7392 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_101
timestamp 1698175906
transform 1 0 12656 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_105
timestamp 1698175906
transform 1 0 13104 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_124
timestamp 1698175906
transform 1 0 15232 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_152
timestamp 1698175906
transform 1 0 18368 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_156
timestamp 1698175906
transform 1 0 18816 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_164
timestamp 1698175906
transform 1 0 19712 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_75_188
timestamp 1698175906
transform 1 0 22400 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_196
timestamp 1698175906
transform 1 0 23296 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_200
timestamp 1698175906
transform 1 0 23744 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_202
timestamp 1698175906
transform 1 0 23968 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_75_262
timestamp 1698175906
transform 1 0 30688 0 -1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_278
timestamp 1698175906
transform 1 0 32480 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_75_282
timestamp 1698175906
transform 1 0 32928 0 -1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_75_314
timestamp 1698175906
transform 1 0 36512 0 -1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_330
timestamp 1698175906
transform 1 0 38304 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_8
timestamp 1698175906
transform 1 0 2240 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_76_12
timestamp 1698175906
transform 1 0 2688 0 1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_28
timestamp 1698175906
transform 1 0 4480 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_32
timestamp 1698175906
transform 1 0 4928 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_34
timestamp 1698175906
transform 1 0 5152 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_76_37
timestamp 1698175906
transform 1 0 5488 0 1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_76_53
timestamp 1698175906
transform 1 0 7280 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_61
timestamp 1698175906
transform 1 0 8176 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_65
timestamp 1698175906
transform 1 0 8624 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_71
timestamp 1698175906
transform 1 0 9296 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_76_81
timestamp 1698175906
transform 1 0 10416 0 1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_76_97
timestamp 1698175906
transform 1 0 12208 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_138
timestamp 1698175906
transform 1 0 16800 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_140
timestamp 1698175906
transform 1 0 17024 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_76_177
timestamp 1698175906
transform 1 0 21168 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_185
timestamp 1698175906
transform 1 0 22064 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_189
timestamp 1698175906
transform 1 0 22512 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_215
timestamp 1698175906
transform 1 0 25424 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_217
timestamp 1698175906
transform 1 0 25648 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_236
timestamp 1698175906
transform 1 0 27776 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_240
timestamp 1698175906
transform 1 0 28224 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_244
timestamp 1698175906
transform 1 0 28672 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_76_247
timestamp 1698175906
transform 1 0 29008 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_311
timestamp 1698175906
transform 1 0 36176 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_76_317
timestamp 1698175906
transform 1 0 36848 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_325
timestamp 1698175906
transform 1 0 37744 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_329
timestamp 1698175906
transform 1 0 38192 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_8
timestamp 1698175906
transform 1 0 2240 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_77_12
timestamp 1698175906
transform 1 0 2688 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_77_44
timestamp 1698175906
transform 1 0 6272 0 -1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_77_60
timestamp 1698175906
transform 1 0 8064 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_68
timestamp 1698175906
transform 1 0 8960 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_72
timestamp 1698175906
transform 1 0 9408 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_77_92
timestamp 1698175906
transform 1 0 11648 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_100
timestamp 1698175906
transform 1 0 12544 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_104
timestamp 1698175906
transform 1 0 12992 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_106
timestamp 1698175906
transform 1 0 13216 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_77_121
timestamp 1698175906
transform 1 0 14896 0 -1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_137
timestamp 1698175906
transform 1 0 16688 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_139
timestamp 1698175906
transform 1 0 16912 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_171
timestamp 1698175906
transform 1 0 20496 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_175
timestamp 1698175906
transform 1 0 20944 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_177
timestamp 1698175906
transform 1 0 21168 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_207
timestamp 1698175906
transform 1 0 24528 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_209
timestamp 1698175906
transform 1 0 24752 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_220
timestamp 1698175906
transform 1 0 25984 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_224
timestamp 1698175906
transform 1 0 26432 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_77_256
timestamp 1698175906
transform 1 0 30016 0 -1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_77_272
timestamp 1698175906
transform 1 0 31808 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_77_282
timestamp 1698175906
transform 1 0 32928 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_77_314
timestamp 1698175906
transform 1 0 36512 0 -1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_330
timestamp 1698175906
transform 1 0 38304 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_14
timestamp 1698175906
transform 1 0 2912 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_78_18
timestamp 1698175906
transform 1 0 3360 0 1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_34
timestamp 1698175906
transform 1 0 5152 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_78_37
timestamp 1698175906
transform 1 0 5488 0 1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_78_53
timestamp 1698175906
transform 1 0 7280 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_61
timestamp 1698175906
transform 1 0 8176 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_63
timestamp 1698175906
transform 1 0 8400 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_107
timestamp 1698175906
transform 1 0 13328 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_78_119
timestamp 1698175906
transform 1 0 14672 0 1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_78_151
timestamp 1698175906
transform 1 0 18256 0 1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_78_167
timestamp 1698175906
transform 1 0 20048 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_78_177
timestamp 1698175906
transform 1 0 21168 0 1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_78_209
timestamp 1698175906
transform 1 0 24752 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_78_219
timestamp 1698175906
transform 1 0 25872 0 1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_78_235
timestamp 1698175906
transform 1 0 27664 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_243
timestamp 1698175906
transform 1 0 28560 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_78_247
timestamp 1698175906
transform 1 0 29008 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_311
timestamp 1698175906
transform 1 0 36176 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_78_317
timestamp 1698175906
transform 1 0 36848 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_325
timestamp 1698175906
transform 1 0 37744 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_2
timestamp 1698175906
transform 1 0 1568 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_79_8
timestamp 1698175906
transform 1 0 2240 0 -1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_79_40
timestamp 1698175906
transform 1 0 5824 0 -1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_79_56
timestamp 1698175906
transform 1 0 7616 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_64
timestamp 1698175906
transform 1 0 8512 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_68
timestamp 1698175906
transform 1 0 8960 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_79_72
timestamp 1698175906
transform 1 0 9408 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_136
timestamp 1698175906
transform 1 0 16576 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_79_142
timestamp 1698175906
transform 1 0 17248 0 -1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_79_174
timestamp 1698175906
transform 1 0 20832 0 -1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_79_190
timestamp 1698175906
transform 1 0 22624 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_198
timestamp 1698175906
transform 1 0 23520 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_212
timestamp 1698175906
transform 1 0 25088 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_216
timestamp 1698175906
transform 1 0 25536 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_79_220
timestamp 1698175906
transform 1 0 25984 0 -1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_79_252
timestamp 1698175906
transform 1 0 29568 0 -1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_79_268
timestamp 1698175906
transform 1 0 31360 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_276
timestamp 1698175906
transform 1 0 32256 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_79_282
timestamp 1698175906
transform 1 0 32928 0 -1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_79_314
timestamp 1698175906
transform 1 0 36512 0 -1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_330
timestamp 1698175906
transform 1 0 38304 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_80_2
timestamp 1698175906
transform 1 0 1568 0 1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_34
timestamp 1698175906
transform 1 0 5152 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_80_37
timestamp 1698175906
transform 1 0 5488 0 1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_69
timestamp 1698175906
transform 1 0 9072 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_80_80
timestamp 1698175906
transform 1 0 10304 0 1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_96
timestamp 1698175906
transform 1 0 12096 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_80_107
timestamp 1698175906
transform 1 0 13328 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_171
timestamp 1698175906
transform 1 0 20496 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_80_177
timestamp 1698175906
transform 1 0 21168 0 1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_80_209
timestamp 1698175906
transform 1 0 24752 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_217
timestamp 1698175906
transform 1 0 25648 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_229
timestamp 1698175906
transform 1 0 26992 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_80_233
timestamp 1698175906
transform 1 0 27440 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_241
timestamp 1698175906
transform 1 0 28336 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_80_247
timestamp 1698175906
transform 1 0 29008 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_311
timestamp 1698175906
transform 1 0 36176 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_80_317
timestamp 1698175906
transform 1 0 36848 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_325
timestamp 1698175906
transform 1 0 37744 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_329
timestamp 1698175906
transform 1 0 38192 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_8
timestamp 1698175906
transform 1 0 2240 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_81_12
timestamp 1698175906
transform 1 0 2688 0 -1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_81_44
timestamp 1698175906
transform 1 0 6272 0 -1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_80
timestamp 1698175906
transform 1 0 10304 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_81_115
timestamp 1698175906
transform 1 0 14224 0 -1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_131
timestamp 1698175906
transform 1 0 16016 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_135
timestamp 1698175906
transform 1 0 16464 0 -1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_81_156
timestamp 1698175906
transform 1 0 18816 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_164
timestamp 1698175906
transform 1 0 19712 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_166
timestamp 1698175906
transform 1 0 19936 0 -1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_185
timestamp 1698175906
transform 1 0 22064 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_189
timestamp 1698175906
transform 1 0 22512 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_81_197
timestamp 1698175906
transform 1 0 23408 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_205
timestamp 1698175906
transform 1 0 24304 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_209
timestamp 1698175906
transform 1 0 24752 0 -1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_81_237
timestamp 1698175906
transform 1 0 27888 0 -1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_81_269
timestamp 1698175906
transform 1 0 31472 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_277
timestamp 1698175906
transform 1 0 32368 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_279
timestamp 1698175906
transform 1 0 32592 0 -1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_81_282
timestamp 1698175906
transform 1 0 32928 0 -1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_81_314
timestamp 1698175906
transform 1 0 36512 0 -1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_330
timestamp 1698175906
transform 1 0 38304 0 -1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_8
timestamp 1698175906
transform 1 0 2240 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_82_12
timestamp 1698175906
transform 1 0 2688 0 1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_28
timestamp 1698175906
transform 1 0 4480 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_32
timestamp 1698175906
transform 1 0 4928 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_34
timestamp 1698175906
transform 1 0 5152 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_82_37
timestamp 1698175906
transform 1 0 5488 0 1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_107
timestamp 1698175906
transform 1 0 13328 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_174
timestamp 1698175906
transform 1 0 20832 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_82_177
timestamp 1698175906
transform 1 0 21168 0 1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_193
timestamp 1698175906
transform 1 0 22960 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_215
timestamp 1698175906
transform 1 0 25424 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_82_247
timestamp 1698175906
transform 1 0 29008 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_311
timestamp 1698175906
transform 1 0 36176 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_82_317
timestamp 1698175906
transform 1 0 36848 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_325
timestamp 1698175906
transform 1 0 37744 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_329
timestamp 1698175906
transform 1 0 38192 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_8
timestamp 1698175906
transform 1 0 2240 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_83_12
timestamp 1698175906
transform 1 0 2688 0 -1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_83_44
timestamp 1698175906
transform 1 0 6272 0 -1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_83_60
timestamp 1698175906
transform 1 0 8064 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_68
timestamp 1698175906
transform 1 0 8960 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_83_72
timestamp 1698175906
transform 1 0 9408 0 -1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_138
timestamp 1698175906
transform 1 0 16800 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_172
timestamp 1698175906
transform 1 0 20608 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_83_174
timestamp 1698175906
transform 1 0 20832 0 -1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_83_249
timestamp 1698175906
transform 1 0 29232 0 -1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_83_265
timestamp 1698175906
transform 1 0 31024 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_273
timestamp 1698175906
transform 1 0 31920 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_277
timestamp 1698175906
transform 1 0 32368 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_83_279
timestamp 1698175906
transform 1 0 32592 0 -1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_83_282
timestamp 1698175906
transform 1 0 32928 0 -1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_83_314
timestamp 1698175906
transform 1 0 36512 0 -1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_83_330
timestamp 1698175906
transform 1 0 38304 0 -1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_84_2
timestamp 1698175906
transform 1 0 1568 0 1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_34
timestamp 1698175906
transform 1 0 5152 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_84_37
timestamp 1698175906
transform 1 0 5488 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_101
timestamp 1698175906
transform 1 0 12656 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_84_107
timestamp 1698175906
transform 1 0 13328 0 1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_131
timestamp 1698175906
transform 1 0 16016 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_133
timestamp 1698175906
transform 1 0 16240 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_140
timestamp 1698175906
transform 1 0 17024 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_142
timestamp 1698175906
transform 1 0 17248 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_84_177
timestamp 1698175906
transform 1 0 21168 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_185
timestamp 1698175906
transform 1 0 22064 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_84_225
timestamp 1698175906
transform 1 0 26544 0 1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_241
timestamp 1698175906
transform 1 0 28336 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_84_247
timestamp 1698175906
transform 1 0 29008 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_311
timestamp 1698175906
transform 1 0 36176 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_84_317
timestamp 1698175906
transform 1 0 36848 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_325
timestamp 1698175906
transform 1 0 37744 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_329
timestamp 1698175906
transform 1 0 38192 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_85_2
timestamp 1698175906
transform 1 0 1568 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_66
timestamp 1698175906
transform 1 0 8736 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_85_72
timestamp 1698175906
transform 1 0 9408 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_136
timestamp 1698175906
transform 1 0 16576 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_142
timestamp 1698175906
transform 1 0 17248 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_85_146
timestamp 1698175906
transform 1 0 17696 0 -1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_85_155
timestamp 1698175906
transform 1 0 18704 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_85_163
timestamp 1698175906
transform 1 0 19600 0 -1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_85_174
timestamp 1698175906
transform 1 0 20832 0 -1 70560
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_206
timestamp 1698175906
transform 1 0 24416 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_218
timestamp 1698175906
transform 1 0 25760 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_85_222
timestamp 1698175906
transform 1 0 26208 0 -1 70560
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_85_254
timestamp 1698175906
transform 1 0 29792 0 -1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_85_270
timestamp 1698175906
transform 1 0 31584 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_278
timestamp 1698175906
transform 1 0 32480 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_85_282
timestamp 1698175906
transform 1 0 32928 0 -1 70560
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_85_314
timestamp 1698175906
transform 1 0 36512 0 -1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_85_330
timestamp 1698175906
transform 1 0 38304 0 -1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_86_2
timestamp 1698175906
transform 1 0 1568 0 1 70560
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_34
timestamp 1698175906
transform 1 0 5152 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_37
timestamp 1698175906
transform 1 0 5488 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_101
timestamp 1698175906
transform 1 0 12656 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_107
timestamp 1698175906
transform 1 0 13328 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_171
timestamp 1698175906
transform 1 0 20496 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_177
timestamp 1698175906
transform 1 0 21168 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_241
timestamp 1698175906
transform 1 0 28336 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_247
timestamp 1698175906
transform 1 0 29008 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_311
timestamp 1698175906
transform 1 0 36176 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_86_317
timestamp 1698175906
transform 1 0 36848 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_325
timestamp 1698175906
transform 1 0 37744 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_329
timestamp 1698175906
transform 1 0 38192 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_2
timestamp 1698175906
transform 1 0 1568 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_66
timestamp 1698175906
transform 1 0 8736 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_72
timestamp 1698175906
transform 1 0 9408 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_136
timestamp 1698175906
transform 1 0 16576 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_142
timestamp 1698175906
transform 1 0 17248 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_206
timestamp 1698175906
transform 1 0 24416 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_212
timestamp 1698175906
transform 1 0 25088 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_276
timestamp 1698175906
transform 1 0 32256 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_87_282
timestamp 1698175906
transform 1 0 32928 0 -1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_87_314
timestamp 1698175906
transform 1 0 36512 0 -1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_87_330
timestamp 1698175906
transform 1 0 38304 0 -1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_88_2
timestamp 1698175906
transform 1 0 1568 0 1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_34
timestamp 1698175906
transform 1 0 5152 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_37
timestamp 1698175906
transform 1 0 5488 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_101
timestamp 1698175906
transform 1 0 12656 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_107
timestamp 1698175906
transform 1 0 13328 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_171
timestamp 1698175906
transform 1 0 20496 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_177
timestamp 1698175906
transform 1 0 21168 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_241
timestamp 1698175906
transform 1 0 28336 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_247
timestamp 1698175906
transform 1 0 29008 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_311
timestamp 1698175906
transform 1 0 36176 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_88_317
timestamp 1698175906
transform 1 0 36848 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_325
timestamp 1698175906
transform 1 0 37744 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_329
timestamp 1698175906
transform 1 0 38192 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_2
timestamp 1698175906
transform 1 0 1568 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_66
timestamp 1698175906
transform 1 0 8736 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_72
timestamp 1698175906
transform 1 0 9408 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_136
timestamp 1698175906
transform 1 0 16576 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_142
timestamp 1698175906
transform 1 0 17248 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_206
timestamp 1698175906
transform 1 0 24416 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_212
timestamp 1698175906
transform 1 0 25088 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_276
timestamp 1698175906
transform 1 0 32256 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_89_282
timestamp 1698175906
transform 1 0 32928 0 -1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_89_314
timestamp 1698175906
transform 1 0 36512 0 -1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_89_330
timestamp 1698175906
transform 1 0 38304 0 -1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_90_2
timestamp 1698175906
transform 1 0 1568 0 1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_34
timestamp 1698175906
transform 1 0 5152 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_90_37
timestamp 1698175906
transform 1 0 5488 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_101
timestamp 1698175906
transform 1 0 12656 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_90_107
timestamp 1698175906
transform 1 0 13328 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_171
timestamp 1698175906
transform 1 0 20496 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_90_177
timestamp 1698175906
transform 1 0 21168 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_241
timestamp 1698175906
transform 1 0 28336 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_90_247
timestamp 1698175906
transform 1 0 29008 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_311
timestamp 1698175906
transform 1 0 36176 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_90_317
timestamp 1698175906
transform 1 0 36848 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_325
timestamp 1698175906
transform 1 0 37744 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_329
timestamp 1698175906
transform 1 0 38192 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_91_2
timestamp 1698175906
transform 1 0 1568 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_66
timestamp 1698175906
transform 1 0 8736 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_91_72
timestamp 1698175906
transform 1 0 9408 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_136
timestamp 1698175906
transform 1 0 16576 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_91_142
timestamp 1698175906
transform 1 0 17248 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_206
timestamp 1698175906
transform 1 0 24416 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_91_212
timestamp 1698175906
transform 1 0 25088 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_276
timestamp 1698175906
transform 1 0 32256 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_91_282
timestamp 1698175906
transform 1 0 32928 0 -1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_91_314
timestamp 1698175906
transform 1 0 36512 0 -1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_330
timestamp 1698175906
transform 1 0 38304 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_92_2
timestamp 1698175906
transform 1 0 1568 0 1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_34
timestamp 1698175906
transform 1 0 5152 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_92_37
timestamp 1698175906
transform 1 0 5488 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_101
timestamp 1698175906
transform 1 0 12656 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_92_107
timestamp 1698175906
transform 1 0 13328 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_171
timestamp 1698175906
transform 1 0 20496 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_92_177
timestamp 1698175906
transform 1 0 21168 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_241
timestamp 1698175906
transform 1 0 28336 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_92_247
timestamp 1698175906
transform 1 0 29008 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_311
timestamp 1698175906
transform 1 0 36176 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_92_317
timestamp 1698175906
transform 1 0 36848 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_325
timestamp 1698175906
transform 1 0 37744 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_329
timestamp 1698175906
transform 1 0 38192 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_93_2
timestamp 1698175906
transform 1 0 1568 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_66
timestamp 1698175906
transform 1 0 8736 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_93_72
timestamp 1698175906
transform 1 0 9408 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_136
timestamp 1698175906
transform 1 0 16576 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_93_142
timestamp 1698175906
transform 1 0 17248 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_206
timestamp 1698175906
transform 1 0 24416 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_93_212
timestamp 1698175906
transform 1 0 25088 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_276
timestamp 1698175906
transform 1 0 32256 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_93_282
timestamp 1698175906
transform 1 0 32928 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_93_314
timestamp 1698175906
transform 1 0 36512 0 -1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_330
timestamp 1698175906
transform 1 0 38304 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_94_2
timestamp 1698175906
transform 1 0 1568 0 1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_94_34
timestamp 1698175906
transform 1 0 5152 0 1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_94_37
timestamp 1698175906
transform 1 0 5488 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_94_101
timestamp 1698175906
transform 1 0 12656 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_94_107
timestamp 1698175906
transform 1 0 13328 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_94_171
timestamp 1698175906
transform 1 0 20496 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_94_177
timestamp 1698175906
transform 1 0 21168 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_94_241
timestamp 1698175906
transform 1 0 28336 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_94_247
timestamp 1698175906
transform 1 0 29008 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_94_311
timestamp 1698175906
transform 1 0 36176 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_94_317
timestamp 1698175906
transform 1 0 36848 0 1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_94_325
timestamp 1698175906
transform 1 0 37744 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_94_329
timestamp 1698175906
transform 1 0 38192 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_95_2
timestamp 1698175906
transform 1 0 1568 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_95_66
timestamp 1698175906
transform 1 0 8736 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_95_72
timestamp 1698175906
transform 1 0 9408 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_95_136
timestamp 1698175906
transform 1 0 16576 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_95_142
timestamp 1698175906
transform 1 0 17248 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_95_206
timestamp 1698175906
transform 1 0 24416 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_95_212
timestamp 1698175906
transform 1 0 25088 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_95_276
timestamp 1698175906
transform 1 0 32256 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_95_282
timestamp 1698175906
transform 1 0 32928 0 -1 78400
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_95_314
timestamp 1698175906
transform 1 0 36512 0 -1 78400
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_95_330
timestamp 1698175906
transform 1 0 38304 0 -1 78400
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_96_2
timestamp 1698175906
transform 1 0 1568 0 1 78400
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_96_34
timestamp 1698175906
transform 1 0 5152 0 1 78400
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_96_37
timestamp 1698175906
transform 1 0 5488 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_96_101
timestamp 1698175906
transform 1 0 12656 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_96_107
timestamp 1698175906
transform 1 0 13328 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_96_171
timestamp 1698175906
transform 1 0 20496 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_96_177
timestamp 1698175906
transform 1 0 21168 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_96_241
timestamp 1698175906
transform 1 0 28336 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_96_247
timestamp 1698175906
transform 1 0 29008 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_96_311
timestamp 1698175906
transform 1 0 36176 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_96_317
timestamp 1698175906
transform 1 0 36848 0 1 78400
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_96_325
timestamp 1698175906
transform 1 0 37744 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_96_329
timestamp 1698175906
transform 1 0 38192 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_97_2
timestamp 1698175906
transform 1 0 1568 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_97_66
timestamp 1698175906
transform 1 0 8736 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_97_72
timestamp 1698175906
transform 1 0 9408 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_97_136
timestamp 1698175906
transform 1 0 16576 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_97_142
timestamp 1698175906
transform 1 0 17248 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_97_206
timestamp 1698175906
transform 1 0 24416 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_97_212
timestamp 1698175906
transform 1 0 25088 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_97_276
timestamp 1698175906
transform 1 0 32256 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_97_282
timestamp 1698175906
transform 1 0 32928 0 -1 79968
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_97_314
timestamp 1698175906
transform 1 0 36512 0 -1 79968
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_97_330
timestamp 1698175906
transform 1 0 38304 0 -1 79968
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_98_2
timestamp 1698175906
transform 1 0 1568 0 1 79968
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_98_34
timestamp 1698175906
transform 1 0 5152 0 1 79968
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_98_37
timestamp 1698175906
transform 1 0 5488 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_98_101
timestamp 1698175906
transform 1 0 12656 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_98_107
timestamp 1698175906
transform 1 0 13328 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_98_171
timestamp 1698175906
transform 1 0 20496 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_98_177
timestamp 1698175906
transform 1 0 21168 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_98_241
timestamp 1698175906
transform 1 0 28336 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_98_247
timestamp 1698175906
transform 1 0 29008 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_98_311
timestamp 1698175906
transform 1 0 36176 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_98_317
timestamp 1698175906
transform 1 0 36848 0 1 79968
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_98_325
timestamp 1698175906
transform 1 0 37744 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98_329
timestamp 1698175906
transform 1 0 38192 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_99_2
timestamp 1698175906
transform 1 0 1568 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_99_66
timestamp 1698175906
transform 1 0 8736 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_99_72
timestamp 1698175906
transform 1 0 9408 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_99_136
timestamp 1698175906
transform 1 0 16576 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_99_142
timestamp 1698175906
transform 1 0 17248 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_99_206
timestamp 1698175906
transform 1 0 24416 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_99_212
timestamp 1698175906
transform 1 0 25088 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_99_276
timestamp 1698175906
transform 1 0 32256 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_99_282
timestamp 1698175906
transform 1 0 32928 0 -1 81536
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_99_314
timestamp 1698175906
transform 1 0 36512 0 -1 81536
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_99_330
timestamp 1698175906
transform 1 0 38304 0 -1 81536
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_100_2
timestamp 1698175906
transform 1 0 1568 0 1 81536
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_100_34
timestamp 1698175906
transform 1 0 5152 0 1 81536
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_100_37
timestamp 1698175906
transform 1 0 5488 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_100_101
timestamp 1698175906
transform 1 0 12656 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_100_107
timestamp 1698175906
transform 1 0 13328 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_100_171
timestamp 1698175906
transform 1 0 20496 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_100_177
timestamp 1698175906
transform 1 0 21168 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_100_241
timestamp 1698175906
transform 1 0 28336 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_100_247
timestamp 1698175906
transform 1 0 29008 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_100_311
timestamp 1698175906
transform 1 0 36176 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_100_317
timestamp 1698175906
transform 1 0 36848 0 1 81536
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_100_325
timestamp 1698175906
transform 1 0 37744 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_100_329
timestamp 1698175906
transform 1 0 38192 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_101_2
timestamp 1698175906
transform 1 0 1568 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_101_66
timestamp 1698175906
transform 1 0 8736 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_101_72
timestamp 1698175906
transform 1 0 9408 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_101_136
timestamp 1698175906
transform 1 0 16576 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_101_142
timestamp 1698175906
transform 1 0 17248 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_101_206
timestamp 1698175906
transform 1 0 24416 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_101_212
timestamp 1698175906
transform 1 0 25088 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_101_276
timestamp 1698175906
transform 1 0 32256 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_101_282
timestamp 1698175906
transform 1 0 32928 0 -1 83104
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_101_314
timestamp 1698175906
transform 1 0 36512 0 -1 83104
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_101_330
timestamp 1698175906
transform 1 0 38304 0 -1 83104
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_102_2
timestamp 1698175906
transform 1 0 1568 0 1 83104
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_102_34
timestamp 1698175906
transform 1 0 5152 0 1 83104
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_102_37
timestamp 1698175906
transform 1 0 5488 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_102_101
timestamp 1698175906
transform 1 0 12656 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_102_107
timestamp 1698175906
transform 1 0 13328 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_102_171
timestamp 1698175906
transform 1 0 20496 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_102_177
timestamp 1698175906
transform 1 0 21168 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_102_241
timestamp 1698175906
transform 1 0 28336 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_102_247
timestamp 1698175906
transform 1 0 29008 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_102_311
timestamp 1698175906
transform 1 0 36176 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_102_317
timestamp 1698175906
transform 1 0 36848 0 1 83104
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_102_325
timestamp 1698175906
transform 1 0 37744 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_102_329
timestamp 1698175906
transform 1 0 38192 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_103_2
timestamp 1698175906
transform 1 0 1568 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_103_66
timestamp 1698175906
transform 1 0 8736 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_103_72
timestamp 1698175906
transform 1 0 9408 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_103_136
timestamp 1698175906
transform 1 0 16576 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_103_142
timestamp 1698175906
transform 1 0 17248 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_103_206
timestamp 1698175906
transform 1 0 24416 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_103_212
timestamp 1698175906
transform 1 0 25088 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_103_276
timestamp 1698175906
transform 1 0 32256 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_103_282
timestamp 1698175906
transform 1 0 32928 0 -1 84672
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_103_314
timestamp 1698175906
transform 1 0 36512 0 -1 84672
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_103_330
timestamp 1698175906
transform 1 0 38304 0 -1 84672
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_104_2
timestamp 1698175906
transform 1 0 1568 0 1 84672
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104_34
timestamp 1698175906
transform 1 0 5152 0 1 84672
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_104_37
timestamp 1698175906
transform 1 0 5488 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_104_101
timestamp 1698175906
transform 1 0 12656 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_104_107
timestamp 1698175906
transform 1 0 13328 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_104_171
timestamp 1698175906
transform 1 0 20496 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_104_177
timestamp 1698175906
transform 1 0 21168 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_104_241
timestamp 1698175906
transform 1 0 28336 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_104_247
timestamp 1698175906
transform 1 0 29008 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_104_311
timestamp 1698175906
transform 1 0 36176 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_104_317
timestamp 1698175906
transform 1 0 36848 0 1 84672
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_104_325
timestamp 1698175906
transform 1 0 37744 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_104_329
timestamp 1698175906
transform 1 0 38192 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_105_2
timestamp 1698175906
transform 1 0 1568 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_105_66
timestamp 1698175906
transform 1 0 8736 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_105_72
timestamp 1698175906
transform 1 0 9408 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_105_136
timestamp 1698175906
transform 1 0 16576 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_105_142
timestamp 1698175906
transform 1 0 17248 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_105_206
timestamp 1698175906
transform 1 0 24416 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_105_212
timestamp 1698175906
transform 1 0 25088 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_105_276
timestamp 1698175906
transform 1 0 32256 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_105_282
timestamp 1698175906
transform 1 0 32928 0 -1 86240
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_105_314
timestamp 1698175906
transform 1 0 36512 0 -1 86240
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_105_330
timestamp 1698175906
transform 1 0 38304 0 -1 86240
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_106_2
timestamp 1698175906
transform 1 0 1568 0 1 86240
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_106_34
timestamp 1698175906
transform 1 0 5152 0 1 86240
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_106_37
timestamp 1698175906
transform 1 0 5488 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_106_101
timestamp 1698175906
transform 1 0 12656 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_106_107
timestamp 1698175906
transform 1 0 13328 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_106_171
timestamp 1698175906
transform 1 0 20496 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_106_177
timestamp 1698175906
transform 1 0 21168 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_106_241
timestamp 1698175906
transform 1 0 28336 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_106_247
timestamp 1698175906
transform 1 0 29008 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_106_311
timestamp 1698175906
transform 1 0 36176 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_106_317
timestamp 1698175906
transform 1 0 36848 0 1 86240
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_106_325
timestamp 1698175906
transform 1 0 37744 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_106_329
timestamp 1698175906
transform 1 0 38192 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_107_2
timestamp 1698175906
transform 1 0 1568 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_107_66
timestamp 1698175906
transform 1 0 8736 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_107_72
timestamp 1698175906
transform 1 0 9408 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_107_136
timestamp 1698175906
transform 1 0 16576 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_107_142
timestamp 1698175906
transform 1 0 17248 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_107_206
timestamp 1698175906
transform 1 0 24416 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_107_212
timestamp 1698175906
transform 1 0 25088 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_107_276
timestamp 1698175906
transform 1 0 32256 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_107_282
timestamp 1698175906
transform 1 0 32928 0 -1 87808
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_107_314
timestamp 1698175906
transform 1 0 36512 0 -1 87808
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_107_330
timestamp 1698175906
transform 1 0 38304 0 -1 87808
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_108_2
timestamp 1698175906
transform 1 0 1568 0 1 87808
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_108_34
timestamp 1698175906
transform 1 0 5152 0 1 87808
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_108_37
timestamp 1698175906
transform 1 0 5488 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_108_101
timestamp 1698175906
transform 1 0 12656 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_108_107
timestamp 1698175906
transform 1 0 13328 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_108_171
timestamp 1698175906
transform 1 0 20496 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_108_177
timestamp 1698175906
transform 1 0 21168 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_108_241
timestamp 1698175906
transform 1 0 28336 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_108_247
timestamp 1698175906
transform 1 0 29008 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_108_311
timestamp 1698175906
transform 1 0 36176 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_108_317
timestamp 1698175906
transform 1 0 36848 0 1 87808
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_108_325
timestamp 1698175906
transform 1 0 37744 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_108_329
timestamp 1698175906
transform 1 0 38192 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_109_2
timestamp 1698175906
transform 1 0 1568 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_109_66
timestamp 1698175906
transform 1 0 8736 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_109_72
timestamp 1698175906
transform 1 0 9408 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_109_136
timestamp 1698175906
transform 1 0 16576 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_109_142
timestamp 1698175906
transform 1 0 17248 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_109_206
timestamp 1698175906
transform 1 0 24416 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_109_212
timestamp 1698175906
transform 1 0 25088 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_109_276
timestamp 1698175906
transform 1 0 32256 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_109_282
timestamp 1698175906
transform 1 0 32928 0 -1 89376
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_109_314
timestamp 1698175906
transform 1 0 36512 0 -1 89376
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_109_330
timestamp 1698175906
transform 1 0 38304 0 -1 89376
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_110_2
timestamp 1698175906
transform 1 0 1568 0 1 89376
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_110_34
timestamp 1698175906
transform 1 0 5152 0 1 89376
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_110_37
timestamp 1698175906
transform 1 0 5488 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_110_101
timestamp 1698175906
transform 1 0 12656 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_110_107
timestamp 1698175906
transform 1 0 13328 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_110_171
timestamp 1698175906
transform 1 0 20496 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_110_177
timestamp 1698175906
transform 1 0 21168 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_110_241
timestamp 1698175906
transform 1 0 28336 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_110_247
timestamp 1698175906
transform 1 0 29008 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_110_311
timestamp 1698175906
transform 1 0 36176 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_110_317
timestamp 1698175906
transform 1 0 36848 0 1 89376
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_110_325
timestamp 1698175906
transform 1 0 37744 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_110_329
timestamp 1698175906
transform 1 0 38192 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_111_2
timestamp 1698175906
transform 1 0 1568 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_111_66
timestamp 1698175906
transform 1 0 8736 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_111_72
timestamp 1698175906
transform 1 0 9408 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_111_136
timestamp 1698175906
transform 1 0 16576 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_111_142
timestamp 1698175906
transform 1 0 17248 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_111_206
timestamp 1698175906
transform 1 0 24416 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_111_212
timestamp 1698175906
transform 1 0 25088 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_111_276
timestamp 1698175906
transform 1 0 32256 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_111_282
timestamp 1698175906
transform 1 0 32928 0 -1 90944
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_111_314
timestamp 1698175906
transform 1 0 36512 0 -1 90944
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_111_330
timestamp 1698175906
transform 1 0 38304 0 -1 90944
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_112_2
timestamp 1698175906
transform 1 0 1568 0 1 90944
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_112_34
timestamp 1698175906
transform 1 0 5152 0 1 90944
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_112_37
timestamp 1698175906
transform 1 0 5488 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_112_101
timestamp 1698175906
transform 1 0 12656 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_112_107
timestamp 1698175906
transform 1 0 13328 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_112_171
timestamp 1698175906
transform 1 0 20496 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_112_177
timestamp 1698175906
transform 1 0 21168 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_112_241
timestamp 1698175906
transform 1 0 28336 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_112_247
timestamp 1698175906
transform 1 0 29008 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_112_311
timestamp 1698175906
transform 1 0 36176 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_112_317
timestamp 1698175906
transform 1 0 36848 0 1 90944
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_112_325
timestamp 1698175906
transform 1 0 37744 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_112_329
timestamp 1698175906
transform 1 0 38192 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_113_2
timestamp 1698175906
transform 1 0 1568 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_113_66
timestamp 1698175906
transform 1 0 8736 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_113_72
timestamp 1698175906
transform 1 0 9408 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_113_136
timestamp 1698175906
transform 1 0 16576 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_113_142
timestamp 1698175906
transform 1 0 17248 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_113_206
timestamp 1698175906
transform 1 0 24416 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_113_212
timestamp 1698175906
transform 1 0 25088 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_113_276
timestamp 1698175906
transform 1 0 32256 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_113_282
timestamp 1698175906
transform 1 0 32928 0 -1 92512
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_113_314
timestamp 1698175906
transform 1 0 36512 0 -1 92512
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_113_330
timestamp 1698175906
transform 1 0 38304 0 -1 92512
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_114_2
timestamp 1698175906
transform 1 0 1568 0 1 92512
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_114_34
timestamp 1698175906
transform 1 0 5152 0 1 92512
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_114_37
timestamp 1698175906
transform 1 0 5488 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_114_101
timestamp 1698175906
transform 1 0 12656 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_114_107
timestamp 1698175906
transform 1 0 13328 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_114_171
timestamp 1698175906
transform 1 0 20496 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_114_177
timestamp 1698175906
transform 1 0 21168 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_114_241
timestamp 1698175906
transform 1 0 28336 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_114_247
timestamp 1698175906
transform 1 0 29008 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_114_311
timestamp 1698175906
transform 1 0 36176 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_114_317
timestamp 1698175906
transform 1 0 36848 0 1 92512
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_114_325
timestamp 1698175906
transform 1 0 37744 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_114_329
timestamp 1698175906
transform 1 0 38192 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_115_2
timestamp 1698175906
transform 1 0 1568 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_115_66
timestamp 1698175906
transform 1 0 8736 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_115_72
timestamp 1698175906
transform 1 0 9408 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_115_136
timestamp 1698175906
transform 1 0 16576 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_115_142
timestamp 1698175906
transform 1 0 17248 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_115_206
timestamp 1698175906
transform 1 0 24416 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_115_212
timestamp 1698175906
transform 1 0 25088 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_115_276
timestamp 1698175906
transform 1 0 32256 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_115_282
timestamp 1698175906
transform 1 0 32928 0 -1 94080
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_115_314
timestamp 1698175906
transform 1 0 36512 0 -1 94080
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_115_330
timestamp 1698175906
transform 1 0 38304 0 -1 94080
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_116_2
timestamp 1698175906
transform 1 0 1568 0 1 94080
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_116_34
timestamp 1698175906
transform 1 0 5152 0 1 94080
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_116_37
timestamp 1698175906
transform 1 0 5488 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_116_101
timestamp 1698175906
transform 1 0 12656 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_116_107
timestamp 1698175906
transform 1 0 13328 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_116_171
timestamp 1698175906
transform 1 0 20496 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_116_177
timestamp 1698175906
transform 1 0 21168 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_116_241
timestamp 1698175906
transform 1 0 28336 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_116_247
timestamp 1698175906
transform 1 0 29008 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_116_311
timestamp 1698175906
transform 1 0 36176 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_116_317
timestamp 1698175906
transform 1 0 36848 0 1 94080
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_116_325
timestamp 1698175906
transform 1 0 37744 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_116_329
timestamp 1698175906
transform 1 0 38192 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_117_2
timestamp 1698175906
transform 1 0 1568 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_117_66
timestamp 1698175906
transform 1 0 8736 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_117_72
timestamp 1698175906
transform 1 0 9408 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_117_136
timestamp 1698175906
transform 1 0 16576 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_117_142
timestamp 1698175906
transform 1 0 17248 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_117_206
timestamp 1698175906
transform 1 0 24416 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_117_212
timestamp 1698175906
transform 1 0 25088 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_117_276
timestamp 1698175906
transform 1 0 32256 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_117_282
timestamp 1698175906
transform 1 0 32928 0 -1 95648
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_117_314
timestamp 1698175906
transform 1 0 36512 0 -1 95648
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_117_330
timestamp 1698175906
transform 1 0 38304 0 -1 95648
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_118_2
timestamp 1698175906
transform 1 0 1568 0 1 95648
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_118_18
timestamp 1698175906
transform 1 0 3360 0 1 95648
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_118_23
timestamp 1698175906
transform 1 0 3920 0 1 95648
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_118_31
timestamp 1698175906
transform 1 0 4816 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_118_33
timestamp 1698175906
transform 1 0 5040 0 1 95648
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_118_36
timestamp 1698175906
transform 1 0 5376 0 1 95648
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_118_70
timestamp 1698175906
transform 1 0 9184 0 1 95648
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_118_104
timestamp 1698175906
transform 1 0 12992 0 1 95648
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_118_138
timestamp 1698175906
transform 1 0 16800 0 1 95648
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_118_172
timestamp 1698175906
transform 1 0 20608 0 1 95648
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_118_206
timestamp 1698175906
transform 1 0 24416 0 1 95648
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_118_240
timestamp 1698175906
transform 1 0 28224 0 1 95648
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_118_274
timestamp 1698175906
transform 1 0 32032 0 1 95648
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_118_308
timestamp 1698175906
transform 1 0 35840 0 1 95648
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_118_324
timestamp 1698175906
transform 1 0 37632 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_118_328
timestamp 1698175906
transform 1 0 38080 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_118_330
timestamp 1698175906
transform 1 0 38304 0 1 95648
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698175906
transform 1 0 1568 0 1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698175906
transform 1 0 1568 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698175906
transform 1 0 1568 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698175906
transform 1 0 1568 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698175906
transform 1 0 1568 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698175906
transform 1 0 1568 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698175906
transform 1 0 1568 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1698175906
transform 1 0 1568 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1698175906
transform 1 0 2240 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1698175906
transform 1 0 1568 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1698175906
transform 1 0 1568 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1698175906
transform 1 0 1568 0 -1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1698175906
transform 1 0 1568 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input14
timestamp 1698175906
transform 1 0 1568 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input15
timestamp 1698175906
transform 1 0 1568 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input16
timestamp 1698175906
transform 1 0 1568 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input17
timestamp 1698175906
transform 1 0 1568 0 -1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input18
timestamp 1698175906
transform 1 0 1568 0 1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input19
timestamp 1698175906
transform 1 0 2240 0 1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input20
timestamp 1698175906
transform 1 0 1568 0 1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input21
timestamp 1698175906
transform 1 0 1568 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input22
timestamp 1698175906
transform 1 0 1568 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input23
timestamp 1698175906
transform 1 0 1568 0 -1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input24
timestamp 1698175906
transform 1 0 1568 0 1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input25
timestamp 1698175906
transform 1 0 1568 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input26
timestamp 1698175906
transform 1 0 1568 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output27 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 36624 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output28
timestamp 1698175906
transform 1 0 35504 0 -1 54880
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output29
timestamp 1698175906
transform -1 0 36624 0 1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output30
timestamp 1698175906
transform -1 0 36624 0 1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output31
timestamp 1698175906
transform -1 0 36624 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output32
timestamp 1698175906
transform -1 0 38416 0 -1 48608
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output33
timestamp 1698175906
transform -1 0 38416 0 -1 51744
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_119 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 38640 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_120
timestamp 1698175906
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 38640 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_121
timestamp 1698175906
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 38640 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_122
timestamp 1698175906
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 38640 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_123
timestamp 1698175906
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 38640 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_124
timestamp 1698175906
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 38640 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_125
timestamp 1698175906
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 38640 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_126
timestamp 1698175906
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 38640 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_127
timestamp 1698175906
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 38640 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_128
timestamp 1698175906
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 38640 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_129
timestamp 1698175906
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 38640 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_130
timestamp 1698175906
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 38640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_131
timestamp 1698175906
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 38640 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_132
timestamp 1698175906
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 38640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_133
timestamp 1698175906
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 38640 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_134
timestamp 1698175906
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 38640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_135
timestamp 1698175906
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 38640 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_136
timestamp 1698175906
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 38640 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_137
timestamp 1698175906
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 38640 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_138
timestamp 1698175906
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 38640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_139
timestamp 1698175906
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 38640 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_140
timestamp 1698175906
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 38640 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_141
timestamp 1698175906
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 38640 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_142
timestamp 1698175906
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 38640 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_143
timestamp 1698175906
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 38640 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_144
timestamp 1698175906
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 38640 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_145
timestamp 1698175906
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 38640 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_146
timestamp 1698175906
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 38640 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_147
timestamp 1698175906
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 38640 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_148
timestamp 1698175906
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 38640 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_149
timestamp 1698175906
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 38640 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_150
timestamp 1698175906
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 38640 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_151
timestamp 1698175906
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 38640 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_152
timestamp 1698175906
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 38640 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_153
timestamp 1698175906
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 38640 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_154
timestamp 1698175906
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 38640 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_155
timestamp 1698175906
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 38640 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_156
timestamp 1698175906
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 38640 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_157
timestamp 1698175906
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 38640 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_158
timestamp 1698175906
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 38640 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_159
timestamp 1698175906
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 38640 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_160
timestamp 1698175906
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 38640 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_161
timestamp 1698175906
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 38640 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_162
timestamp 1698175906
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 38640 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_163
timestamp 1698175906
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 38640 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_164
timestamp 1698175906
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698175906
transform -1 0 38640 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_165
timestamp 1698175906
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698175906
transform -1 0 38640 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_166
timestamp 1698175906
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698175906
transform -1 0 38640 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_167
timestamp 1698175906
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698175906
transform -1 0 38640 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_168
timestamp 1698175906
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698175906
transform -1 0 38640 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_169
timestamp 1698175906
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698175906
transform -1 0 38640 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_170
timestamp 1698175906
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698175906
transform -1 0 38640 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_171
timestamp 1698175906
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1698175906
transform -1 0 38640 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_172
timestamp 1698175906
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1698175906
transform -1 0 38640 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_173
timestamp 1698175906
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1698175906
transform -1 0 38640 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Left_174
timestamp 1698175906
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Right_55
timestamp 1698175906
transform -1 0 38640 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Left_175
timestamp 1698175906
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Right_56
timestamp 1698175906
transform -1 0 38640 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Left_176
timestamp 1698175906
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Right_57
timestamp 1698175906
transform -1 0 38640 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Left_177
timestamp 1698175906
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Right_58
timestamp 1698175906
transform -1 0 38640 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Left_178
timestamp 1698175906
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Right_59
timestamp 1698175906
transform -1 0 38640 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Left_179
timestamp 1698175906
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Right_60
timestamp 1698175906
transform -1 0 38640 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Left_180
timestamp 1698175906
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Right_61
timestamp 1698175906
transform -1 0 38640 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Left_181
timestamp 1698175906
transform 1 0 1344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Right_62
timestamp 1698175906
transform -1 0 38640 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Left_182
timestamp 1698175906
transform 1 0 1344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Right_63
timestamp 1698175906
transform -1 0 38640 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Left_183
timestamp 1698175906
transform 1 0 1344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Right_64
timestamp 1698175906
transform -1 0 38640 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Left_184
timestamp 1698175906
transform 1 0 1344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Right_65
timestamp 1698175906
transform -1 0 38640 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Left_185
timestamp 1698175906
transform 1 0 1344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Right_66
timestamp 1698175906
transform -1 0 38640 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Left_186
timestamp 1698175906
transform 1 0 1344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Right_67
timestamp 1698175906
transform -1 0 38640 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_68_Left_187
timestamp 1698175906
transform 1 0 1344 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_68_Right_68
timestamp 1698175906
transform -1 0 38640 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_69_Left_188
timestamp 1698175906
transform 1 0 1344 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_69_Right_69
timestamp 1698175906
transform -1 0 38640 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_70_Left_189
timestamp 1698175906
transform 1 0 1344 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_70_Right_70
timestamp 1698175906
transform -1 0 38640 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_71_Left_190
timestamp 1698175906
transform 1 0 1344 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_71_Right_71
timestamp 1698175906
transform -1 0 38640 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_72_Left_191
timestamp 1698175906
transform 1 0 1344 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_72_Right_72
timestamp 1698175906
transform -1 0 38640 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_73_Left_192
timestamp 1698175906
transform 1 0 1344 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_73_Right_73
timestamp 1698175906
transform -1 0 38640 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_74_Left_193
timestamp 1698175906
transform 1 0 1344 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_74_Right_74
timestamp 1698175906
transform -1 0 38640 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_75_Left_194
timestamp 1698175906
transform 1 0 1344 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_75_Right_75
timestamp 1698175906
transform -1 0 38640 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_76_Left_195
timestamp 1698175906
transform 1 0 1344 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_76_Right_76
timestamp 1698175906
transform -1 0 38640 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_77_Left_196
timestamp 1698175906
transform 1 0 1344 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_77_Right_77
timestamp 1698175906
transform -1 0 38640 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_78_Left_197
timestamp 1698175906
transform 1 0 1344 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_78_Right_78
timestamp 1698175906
transform -1 0 38640 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_79_Left_198
timestamp 1698175906
transform 1 0 1344 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_79_Right_79
timestamp 1698175906
transform -1 0 38640 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_80_Left_199
timestamp 1698175906
transform 1 0 1344 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_80_Right_80
timestamp 1698175906
transform -1 0 38640 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_81_Left_200
timestamp 1698175906
transform 1 0 1344 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_81_Right_81
timestamp 1698175906
transform -1 0 38640 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_82_Left_201
timestamp 1698175906
transform 1 0 1344 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_82_Right_82
timestamp 1698175906
transform -1 0 38640 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_83_Left_202
timestamp 1698175906
transform 1 0 1344 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_83_Right_83
timestamp 1698175906
transform -1 0 38640 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_84_Left_203
timestamp 1698175906
transform 1 0 1344 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_84_Right_84
timestamp 1698175906
transform -1 0 38640 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_85_Left_204
timestamp 1698175906
transform 1 0 1344 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_85_Right_85
timestamp 1698175906
transform -1 0 38640 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_86_Left_205
timestamp 1698175906
transform 1 0 1344 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_86_Right_86
timestamp 1698175906
transform -1 0 38640 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_87_Left_206
timestamp 1698175906
transform 1 0 1344 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_87_Right_87
timestamp 1698175906
transform -1 0 38640 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_88_Left_207
timestamp 1698175906
transform 1 0 1344 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_88_Right_88
timestamp 1698175906
transform -1 0 38640 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_89_Left_208
timestamp 1698175906
transform 1 0 1344 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_89_Right_89
timestamp 1698175906
transform -1 0 38640 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_90_Left_209
timestamp 1698175906
transform 1 0 1344 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_90_Right_90
timestamp 1698175906
transform -1 0 38640 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_91_Left_210
timestamp 1698175906
transform 1 0 1344 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_91_Right_91
timestamp 1698175906
transform -1 0 38640 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_92_Left_211
timestamp 1698175906
transform 1 0 1344 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_92_Right_92
timestamp 1698175906
transform -1 0 38640 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_93_Left_212
timestamp 1698175906
transform 1 0 1344 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_93_Right_93
timestamp 1698175906
transform -1 0 38640 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_94_Left_213
timestamp 1698175906
transform 1 0 1344 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_94_Right_94
timestamp 1698175906
transform -1 0 38640 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_95_Left_214
timestamp 1698175906
transform 1 0 1344 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_95_Right_95
timestamp 1698175906
transform -1 0 38640 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_96_Left_215
timestamp 1698175906
transform 1 0 1344 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_96_Right_96
timestamp 1698175906
transform -1 0 38640 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_97_Left_216
timestamp 1698175906
transform 1 0 1344 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_97_Right_97
timestamp 1698175906
transform -1 0 38640 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_98_Left_217
timestamp 1698175906
transform 1 0 1344 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_98_Right_98
timestamp 1698175906
transform -1 0 38640 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_99_Left_218
timestamp 1698175906
transform 1 0 1344 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_99_Right_99
timestamp 1698175906
transform -1 0 38640 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_100_Left_219
timestamp 1698175906
transform 1 0 1344 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_100_Right_100
timestamp 1698175906
transform -1 0 38640 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_101_Left_220
timestamp 1698175906
transform 1 0 1344 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_101_Right_101
timestamp 1698175906
transform -1 0 38640 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_102_Left_221
timestamp 1698175906
transform 1 0 1344 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_102_Right_102
timestamp 1698175906
transform -1 0 38640 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_103_Left_222
timestamp 1698175906
transform 1 0 1344 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_103_Right_103
timestamp 1698175906
transform -1 0 38640 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_104_Left_223
timestamp 1698175906
transform 1 0 1344 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_104_Right_104
timestamp 1698175906
transform -1 0 38640 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_105_Left_224
timestamp 1698175906
transform 1 0 1344 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_105_Right_105
timestamp 1698175906
transform -1 0 38640 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_106_Left_225
timestamp 1698175906
transform 1 0 1344 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_106_Right_106
timestamp 1698175906
transform -1 0 38640 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_107_Left_226
timestamp 1698175906
transform 1 0 1344 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_107_Right_107
timestamp 1698175906
transform -1 0 38640 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_108_Left_227
timestamp 1698175906
transform 1 0 1344 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_108_Right_108
timestamp 1698175906
transform -1 0 38640 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_109_Left_228
timestamp 1698175906
transform 1 0 1344 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_109_Right_109
timestamp 1698175906
transform -1 0 38640 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_110_Left_229
timestamp 1698175906
transform 1 0 1344 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_110_Right_110
timestamp 1698175906
transform -1 0 38640 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_111_Left_230
timestamp 1698175906
transform 1 0 1344 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_111_Right_111
timestamp 1698175906
transform -1 0 38640 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_112_Left_231
timestamp 1698175906
transform 1 0 1344 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_112_Right_112
timestamp 1698175906
transform -1 0 38640 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_113_Left_232
timestamp 1698175906
transform 1 0 1344 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_113_Right_113
timestamp 1698175906
transform -1 0 38640 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_114_Left_233
timestamp 1698175906
transform 1 0 1344 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_114_Right_114
timestamp 1698175906
transform -1 0 38640 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_115_Left_234
timestamp 1698175906
transform 1 0 1344 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_115_Right_115
timestamp 1698175906
transform -1 0 38640 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_116_Left_235
timestamp 1698175906
transform 1 0 1344 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_116_Right_116
timestamp 1698175906
transform -1 0 38640 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_117_Left_236
timestamp 1698175906
transform 1 0 1344 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_117_Right_117
timestamp 1698175906
transform -1 0 38640 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_118_Left_237
timestamp 1698175906
transform 1 0 1344 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_118_Right_118
timestamp 1698175906
transform -1 0 38640 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer1
timestamp 1698175906
transform 1 0 14784 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  rebuffer2
timestamp 1698175906
transform 1 0 22064 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  rebuffer3
timestamp 1698175906
transform 1 0 14896 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  rebuffer4
timestamp 1698175906
transform 1 0 16016 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  rebuffer5
timestamp 1698175906
transform 1 0 22736 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  rebuffer6 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15904 0 -1 62720
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  rebuffer7
timestamp 1698175906
transform -1 0 26992 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  riscv_top_34 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 37968 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  riscv_top_35
timestamp 1698175906
transform -1 0 3248 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  riscv_top_36
timestamp 1698175906
transform 1 0 37968 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  riscv_top_37
timestamp 1698175906
transform 1 0 37968 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  riscv_top_38
timestamp 1698175906
transform 1 0 37968 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  riscv_top_39
timestamp 1698175906
transform -1 0 3920 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  riscv_top_40
timestamp 1698175906
transform -1 0 2016 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_238 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_239
timestamp 1698175906
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_240
timestamp 1698175906
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_241
timestamp 1698175906
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_242
timestamp 1698175906
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_243
timestamp 1698175906
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_244
timestamp 1698175906
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_245
timestamp 1698175906
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_246
timestamp 1698175906
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_247
timestamp 1698175906
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_248
timestamp 1698175906
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_249
timestamp 1698175906
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_250
timestamp 1698175906
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_251
timestamp 1698175906
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_252
timestamp 1698175906
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_253
timestamp 1698175906
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_254
timestamp 1698175906
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_255
timestamp 1698175906
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_256
timestamp 1698175906
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_257
timestamp 1698175906
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_258
timestamp 1698175906
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_259
timestamp 1698175906
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_260
timestamp 1698175906
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_261
timestamp 1698175906
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_262
timestamp 1698175906
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_263
timestamp 1698175906
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_264
timestamp 1698175906
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_265
timestamp 1698175906
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_266
timestamp 1698175906
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_267
timestamp 1698175906
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_268
timestamp 1698175906
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_269
timestamp 1698175906
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_270
timestamp 1698175906
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_271
timestamp 1698175906
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_272
timestamp 1698175906
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_273
timestamp 1698175906
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_274
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_275
timestamp 1698175906
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_276
timestamp 1698175906
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_277
timestamp 1698175906
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_278
timestamp 1698175906
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_279
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_280
timestamp 1698175906
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_281
timestamp 1698175906
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_282
timestamp 1698175906
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_283
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_284
timestamp 1698175906
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_285
timestamp 1698175906
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_286
timestamp 1698175906
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_287
timestamp 1698175906
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_288
timestamp 1698175906
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_289
timestamp 1698175906
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_290
timestamp 1698175906
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_291
timestamp 1698175906
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_292
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_293
timestamp 1698175906
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_294
timestamp 1698175906
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_295
timestamp 1698175906
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_296
timestamp 1698175906
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_297
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_298
timestamp 1698175906
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_299
timestamp 1698175906
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_300
timestamp 1698175906
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_301
timestamp 1698175906
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_302
timestamp 1698175906
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_303
timestamp 1698175906
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_304
timestamp 1698175906
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_305
timestamp 1698175906
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_306
timestamp 1698175906
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_307
timestamp 1698175906
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_308
timestamp 1698175906
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_309
timestamp 1698175906
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_310
timestamp 1698175906
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_311
timestamp 1698175906
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_312
timestamp 1698175906
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_313
timestamp 1698175906
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_314
timestamp 1698175906
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_315
timestamp 1698175906
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_316
timestamp 1698175906
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_317
timestamp 1698175906
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_318
timestamp 1698175906
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_319
timestamp 1698175906
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_320
timestamp 1698175906
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_321
timestamp 1698175906
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_322
timestamp 1698175906
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_323
timestamp 1698175906
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_324
timestamp 1698175906
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_325
timestamp 1698175906
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_326
timestamp 1698175906
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_327
timestamp 1698175906
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_328
timestamp 1698175906
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_329
timestamp 1698175906
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_330
timestamp 1698175906
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_331
timestamp 1698175906
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_332
timestamp 1698175906
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_333
timestamp 1698175906
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_334
timestamp 1698175906
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_335
timestamp 1698175906
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_336
timestamp 1698175906
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_337
timestamp 1698175906
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_338
timestamp 1698175906
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_339
timestamp 1698175906
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_340
timestamp 1698175906
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_341
timestamp 1698175906
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_342
timestamp 1698175906
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_343
timestamp 1698175906
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_344
timestamp 1698175906
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_345
timestamp 1698175906
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_346
timestamp 1698175906
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_347
timestamp 1698175906
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_348
timestamp 1698175906
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_349
timestamp 1698175906
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_350
timestamp 1698175906
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_351
timestamp 1698175906
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_352
timestamp 1698175906
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_353
timestamp 1698175906
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_354
timestamp 1698175906
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_355
timestamp 1698175906
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_356
timestamp 1698175906
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_357
timestamp 1698175906
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_358
timestamp 1698175906
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_359
timestamp 1698175906
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_360
timestamp 1698175906
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_361
timestamp 1698175906
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_362
timestamp 1698175906
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_363
timestamp 1698175906
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_364
timestamp 1698175906
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_365
timestamp 1698175906
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_366
timestamp 1698175906
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_367
timestamp 1698175906
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_368
timestamp 1698175906
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_369
timestamp 1698175906
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_370
timestamp 1698175906
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_371
timestamp 1698175906
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_372
timestamp 1698175906
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_373
timestamp 1698175906
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_374
timestamp 1698175906
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_375
timestamp 1698175906
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_376
timestamp 1698175906
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_377
timestamp 1698175906
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_378
timestamp 1698175906
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_379
timestamp 1698175906
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_380
timestamp 1698175906
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_381
timestamp 1698175906
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_382
timestamp 1698175906
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_383
timestamp 1698175906
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_384
timestamp 1698175906
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_385
timestamp 1698175906
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_386
timestamp 1698175906
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_387
timestamp 1698175906
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_388
timestamp 1698175906
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_389
timestamp 1698175906
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_390
timestamp 1698175906
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_391
timestamp 1698175906
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_392
timestamp 1698175906
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_393
timestamp 1698175906
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_394
timestamp 1698175906
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_395
timestamp 1698175906
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_396
timestamp 1698175906
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_397
timestamp 1698175906
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_398
timestamp 1698175906
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_399
timestamp 1698175906
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_400
timestamp 1698175906
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_401
timestamp 1698175906
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_402
timestamp 1698175906
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_403
timestamp 1698175906
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_404
timestamp 1698175906
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_405
timestamp 1698175906
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_406
timestamp 1698175906
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_407
timestamp 1698175906
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_408
timestamp 1698175906
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_409
timestamp 1698175906
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_410
timestamp 1698175906
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_411
timestamp 1698175906
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_412
timestamp 1698175906
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_413
timestamp 1698175906
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_414
timestamp 1698175906
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_415
timestamp 1698175906
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_416
timestamp 1698175906
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_417
timestamp 1698175906
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_418
timestamp 1698175906
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_419
timestamp 1698175906
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_420
timestamp 1698175906
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_421
timestamp 1698175906
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_422
timestamp 1698175906
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_423
timestamp 1698175906
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_424
timestamp 1698175906
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_425
timestamp 1698175906
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_426
timestamp 1698175906
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_427
timestamp 1698175906
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_428
timestamp 1698175906
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_429
timestamp 1698175906
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_430
timestamp 1698175906
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_431
timestamp 1698175906
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_432
timestamp 1698175906
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_433
timestamp 1698175906
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_434
timestamp 1698175906
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_435
timestamp 1698175906
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_436
timestamp 1698175906
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_437
timestamp 1698175906
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_438
timestamp 1698175906
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_439
timestamp 1698175906
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_440
timestamp 1698175906
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_441
timestamp 1698175906
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_442
timestamp 1698175906
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_443
timestamp 1698175906
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_444
timestamp 1698175906
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_445
timestamp 1698175906
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_446
timestamp 1698175906
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_447
timestamp 1698175906
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_448
timestamp 1698175906
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_449
timestamp 1698175906
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_450
timestamp 1698175906
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_451
timestamp 1698175906
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_452
timestamp 1698175906
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_453
timestamp 1698175906
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_454
timestamp 1698175906
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_455
timestamp 1698175906
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_456
timestamp 1698175906
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_457
timestamp 1698175906
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_458
timestamp 1698175906
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_459
timestamp 1698175906
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_460
timestamp 1698175906
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_461
timestamp 1698175906
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_462
timestamp 1698175906
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_463
timestamp 1698175906
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_464
timestamp 1698175906
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_465
timestamp 1698175906
transform 1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_466
timestamp 1698175906
transform 1 0 32704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_467
timestamp 1698175906
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_468
timestamp 1698175906
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_469
timestamp 1698175906
transform 1 0 20944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_470
timestamp 1698175906
transform 1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_471
timestamp 1698175906
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_472
timestamp 1698175906
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_473
timestamp 1698175906
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_474
timestamp 1698175906
transform 1 0 24864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_475
timestamp 1698175906
transform 1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_476
timestamp 1698175906
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_477
timestamp 1698175906
transform 1 0 13104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_478
timestamp 1698175906
transform 1 0 20944 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_479
timestamp 1698175906
transform 1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_480
timestamp 1698175906
transform 1 0 36624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_481
timestamp 1698175906
transform 1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_482
timestamp 1698175906
transform 1 0 17024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_483
timestamp 1698175906
transform 1 0 24864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_484
timestamp 1698175906
transform 1 0 32704 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_485
timestamp 1698175906
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_486
timestamp 1698175906
transform 1 0 13104 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_487
timestamp 1698175906
transform 1 0 20944 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_488
timestamp 1698175906
transform 1 0 28784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_489
timestamp 1698175906
transform 1 0 36624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_490
timestamp 1698175906
transform 1 0 9184 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_491
timestamp 1698175906
transform 1 0 17024 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_492
timestamp 1698175906
transform 1 0 24864 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_493
timestamp 1698175906
transform 1 0 32704 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_494
timestamp 1698175906
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_495
timestamp 1698175906
transform 1 0 13104 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_496
timestamp 1698175906
transform 1 0 20944 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_497
timestamp 1698175906
transform 1 0 28784 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_498
timestamp 1698175906
transform 1 0 36624 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_499
timestamp 1698175906
transform 1 0 9184 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_500
timestamp 1698175906
transform 1 0 17024 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_501
timestamp 1698175906
transform 1 0 24864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_502
timestamp 1698175906
transform 1 0 32704 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_503
timestamp 1698175906
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_504
timestamp 1698175906
transform 1 0 13104 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_505
timestamp 1698175906
transform 1 0 20944 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_506
timestamp 1698175906
transform 1 0 28784 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_507
timestamp 1698175906
transform 1 0 36624 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_508
timestamp 1698175906
transform 1 0 9184 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_509
timestamp 1698175906
transform 1 0 17024 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_510
timestamp 1698175906
transform 1 0 24864 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_511
timestamp 1698175906
transform 1 0 32704 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_512
timestamp 1698175906
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_513
timestamp 1698175906
transform 1 0 13104 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_514
timestamp 1698175906
transform 1 0 20944 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_515
timestamp 1698175906
transform 1 0 28784 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_516
timestamp 1698175906
transform 1 0 36624 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_517
timestamp 1698175906
transform 1 0 9184 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_518
timestamp 1698175906
transform 1 0 17024 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_519
timestamp 1698175906
transform 1 0 24864 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_520
timestamp 1698175906
transform 1 0 32704 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_521
timestamp 1698175906
transform 1 0 5264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_522
timestamp 1698175906
transform 1 0 13104 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_523
timestamp 1698175906
transform 1 0 20944 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_524
timestamp 1698175906
transform 1 0 28784 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_525
timestamp 1698175906
transform 1 0 36624 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_526
timestamp 1698175906
transform 1 0 9184 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_527
timestamp 1698175906
transform 1 0 17024 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_528
timestamp 1698175906
transform 1 0 24864 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_529
timestamp 1698175906
transform 1 0 32704 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_530
timestamp 1698175906
transform 1 0 5264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_531
timestamp 1698175906
transform 1 0 13104 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_532
timestamp 1698175906
transform 1 0 20944 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_533
timestamp 1698175906
transform 1 0 28784 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_534
timestamp 1698175906
transform 1 0 36624 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_535
timestamp 1698175906
transform 1 0 9184 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_536
timestamp 1698175906
transform 1 0 17024 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_537
timestamp 1698175906
transform 1 0 24864 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_538
timestamp 1698175906
transform 1 0 32704 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_539
timestamp 1698175906
transform 1 0 5264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_540
timestamp 1698175906
transform 1 0 13104 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_541
timestamp 1698175906
transform 1 0 20944 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_542
timestamp 1698175906
transform 1 0 28784 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_543
timestamp 1698175906
transform 1 0 36624 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_544
timestamp 1698175906
transform 1 0 9184 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_545
timestamp 1698175906
transform 1 0 17024 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_546
timestamp 1698175906
transform 1 0 24864 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_547
timestamp 1698175906
transform 1 0 32704 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_548
timestamp 1698175906
transform 1 0 5264 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_549
timestamp 1698175906
transform 1 0 13104 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_550
timestamp 1698175906
transform 1 0 20944 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_551
timestamp 1698175906
transform 1 0 28784 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_552
timestamp 1698175906
transform 1 0 36624 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_553
timestamp 1698175906
transform 1 0 9184 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_554
timestamp 1698175906
transform 1 0 17024 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_555
timestamp 1698175906
transform 1 0 24864 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_556
timestamp 1698175906
transform 1 0 32704 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_557
timestamp 1698175906
transform 1 0 5264 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_558
timestamp 1698175906
transform 1 0 13104 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_559
timestamp 1698175906
transform 1 0 20944 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_560
timestamp 1698175906
transform 1 0 28784 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_561
timestamp 1698175906
transform 1 0 36624 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_562
timestamp 1698175906
transform 1 0 9184 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_563
timestamp 1698175906
transform 1 0 17024 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_564
timestamp 1698175906
transform 1 0 24864 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_565
timestamp 1698175906
transform 1 0 32704 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_566
timestamp 1698175906
transform 1 0 5264 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_567
timestamp 1698175906
transform 1 0 13104 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_568
timestamp 1698175906
transform 1 0 20944 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_569
timestamp 1698175906
transform 1 0 28784 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_570
timestamp 1698175906
transform 1 0 36624 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_571
timestamp 1698175906
transform 1 0 9184 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_572
timestamp 1698175906
transform 1 0 17024 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_573
timestamp 1698175906
transform 1 0 24864 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_574
timestamp 1698175906
transform 1 0 32704 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_575
timestamp 1698175906
transform 1 0 5264 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_576
timestamp 1698175906
transform 1 0 13104 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_577
timestamp 1698175906
transform 1 0 20944 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_578
timestamp 1698175906
transform 1 0 28784 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_579
timestamp 1698175906
transform 1 0 36624 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_580
timestamp 1698175906
transform 1 0 9184 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_581
timestamp 1698175906
transform 1 0 17024 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_582
timestamp 1698175906
transform 1 0 24864 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_583
timestamp 1698175906
transform 1 0 32704 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_584
timestamp 1698175906
transform 1 0 5264 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_585
timestamp 1698175906
transform 1 0 13104 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_586
timestamp 1698175906
transform 1 0 20944 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_587
timestamp 1698175906
transform 1 0 28784 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_588
timestamp 1698175906
transform 1 0 36624 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_589
timestamp 1698175906
transform 1 0 9184 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_590
timestamp 1698175906
transform 1 0 17024 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_591
timestamp 1698175906
transform 1 0 24864 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_592
timestamp 1698175906
transform 1 0 32704 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_593
timestamp 1698175906
transform 1 0 5264 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_594
timestamp 1698175906
transform 1 0 13104 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_595
timestamp 1698175906
transform 1 0 20944 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_596
timestamp 1698175906
transform 1 0 28784 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_597
timestamp 1698175906
transform 1 0 36624 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_598
timestamp 1698175906
transform 1 0 9184 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_599
timestamp 1698175906
transform 1 0 17024 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_600
timestamp 1698175906
transform 1 0 24864 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_601
timestamp 1698175906
transform 1 0 32704 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_602
timestamp 1698175906
transform 1 0 5264 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_603
timestamp 1698175906
transform 1 0 13104 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_604
timestamp 1698175906
transform 1 0 20944 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_605
timestamp 1698175906
transform 1 0 28784 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_606
timestamp 1698175906
transform 1 0 36624 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_607
timestamp 1698175906
transform 1 0 9184 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_608
timestamp 1698175906
transform 1 0 17024 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_609
timestamp 1698175906
transform 1 0 24864 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_610
timestamp 1698175906
transform 1 0 32704 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_611
timestamp 1698175906
transform 1 0 5264 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_612
timestamp 1698175906
transform 1 0 13104 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_613
timestamp 1698175906
transform 1 0 20944 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_614
timestamp 1698175906
transform 1 0 28784 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_615
timestamp 1698175906
transform 1 0 36624 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_616
timestamp 1698175906
transform 1 0 9184 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_617
timestamp 1698175906
transform 1 0 17024 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_618
timestamp 1698175906
transform 1 0 24864 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_619
timestamp 1698175906
transform 1 0 32704 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_620
timestamp 1698175906
transform 1 0 5264 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_621
timestamp 1698175906
transform 1 0 13104 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_622
timestamp 1698175906
transform 1 0 20944 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_623
timestamp 1698175906
transform 1 0 28784 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_624
timestamp 1698175906
transform 1 0 36624 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_625
timestamp 1698175906
transform 1 0 9184 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_626
timestamp 1698175906
transform 1 0 17024 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_627
timestamp 1698175906
transform 1 0 24864 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_628
timestamp 1698175906
transform 1 0 32704 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_629
timestamp 1698175906
transform 1 0 5264 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_630
timestamp 1698175906
transform 1 0 13104 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_631
timestamp 1698175906
transform 1 0 20944 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_632
timestamp 1698175906
transform 1 0 28784 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_633
timestamp 1698175906
transform 1 0 36624 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_634
timestamp 1698175906
transform 1 0 9184 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_635
timestamp 1698175906
transform 1 0 17024 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_636
timestamp 1698175906
transform 1 0 24864 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_637
timestamp 1698175906
transform 1 0 32704 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_638
timestamp 1698175906
transform 1 0 5264 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_639
timestamp 1698175906
transform 1 0 13104 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_640
timestamp 1698175906
transform 1 0 20944 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_641
timestamp 1698175906
transform 1 0 28784 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_642
timestamp 1698175906
transform 1 0 36624 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_643
timestamp 1698175906
transform 1 0 9184 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_644
timestamp 1698175906
transform 1 0 17024 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_645
timestamp 1698175906
transform 1 0 24864 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_646
timestamp 1698175906
transform 1 0 32704 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_647
timestamp 1698175906
transform 1 0 5264 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_648
timestamp 1698175906
transform 1 0 13104 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_649
timestamp 1698175906
transform 1 0 20944 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_650
timestamp 1698175906
transform 1 0 28784 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_651
timestamp 1698175906
transform 1 0 36624 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_652
timestamp 1698175906
transform 1 0 9184 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_653
timestamp 1698175906
transform 1 0 17024 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_654
timestamp 1698175906
transform 1 0 24864 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_655
timestamp 1698175906
transform 1 0 32704 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_656
timestamp 1698175906
transform 1 0 5264 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_657
timestamp 1698175906
transform 1 0 13104 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_658
timestamp 1698175906
transform 1 0 20944 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_659
timestamp 1698175906
transform 1 0 28784 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_660
timestamp 1698175906
transform 1 0 36624 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_661
timestamp 1698175906
transform 1 0 9184 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_662
timestamp 1698175906
transform 1 0 17024 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_663
timestamp 1698175906
transform 1 0 24864 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_664
timestamp 1698175906
transform 1 0 32704 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_94_665
timestamp 1698175906
transform 1 0 5264 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_94_666
timestamp 1698175906
transform 1 0 13104 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_94_667
timestamp 1698175906
transform 1 0 20944 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_94_668
timestamp 1698175906
transform 1 0 28784 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_94_669
timestamp 1698175906
transform 1 0 36624 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_95_670
timestamp 1698175906
transform 1 0 9184 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_95_671
timestamp 1698175906
transform 1 0 17024 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_95_672
timestamp 1698175906
transform 1 0 24864 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_95_673
timestamp 1698175906
transform 1 0 32704 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_96_674
timestamp 1698175906
transform 1 0 5264 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_96_675
timestamp 1698175906
transform 1 0 13104 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_96_676
timestamp 1698175906
transform 1 0 20944 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_96_677
timestamp 1698175906
transform 1 0 28784 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_96_678
timestamp 1698175906
transform 1 0 36624 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_97_679
timestamp 1698175906
transform 1 0 9184 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_97_680
timestamp 1698175906
transform 1 0 17024 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_97_681
timestamp 1698175906
transform 1 0 24864 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_97_682
timestamp 1698175906
transform 1 0 32704 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_98_683
timestamp 1698175906
transform 1 0 5264 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_98_684
timestamp 1698175906
transform 1 0 13104 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_98_685
timestamp 1698175906
transform 1 0 20944 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_98_686
timestamp 1698175906
transform 1 0 28784 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_98_687
timestamp 1698175906
transform 1 0 36624 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_99_688
timestamp 1698175906
transform 1 0 9184 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_99_689
timestamp 1698175906
transform 1 0 17024 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_99_690
timestamp 1698175906
transform 1 0 24864 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_99_691
timestamp 1698175906
transform 1 0 32704 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_100_692
timestamp 1698175906
transform 1 0 5264 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_100_693
timestamp 1698175906
transform 1 0 13104 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_100_694
timestamp 1698175906
transform 1 0 20944 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_100_695
timestamp 1698175906
transform 1 0 28784 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_100_696
timestamp 1698175906
transform 1 0 36624 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_101_697
timestamp 1698175906
transform 1 0 9184 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_101_698
timestamp 1698175906
transform 1 0 17024 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_101_699
timestamp 1698175906
transform 1 0 24864 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_101_700
timestamp 1698175906
transform 1 0 32704 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_102_701
timestamp 1698175906
transform 1 0 5264 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_102_702
timestamp 1698175906
transform 1 0 13104 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_102_703
timestamp 1698175906
transform 1 0 20944 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_102_704
timestamp 1698175906
transform 1 0 28784 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_102_705
timestamp 1698175906
transform 1 0 36624 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_103_706
timestamp 1698175906
transform 1 0 9184 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_103_707
timestamp 1698175906
transform 1 0 17024 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_103_708
timestamp 1698175906
transform 1 0 24864 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_103_709
timestamp 1698175906
transform 1 0 32704 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_104_710
timestamp 1698175906
transform 1 0 5264 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_104_711
timestamp 1698175906
transform 1 0 13104 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_104_712
timestamp 1698175906
transform 1 0 20944 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_104_713
timestamp 1698175906
transform 1 0 28784 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_104_714
timestamp 1698175906
transform 1 0 36624 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_105_715
timestamp 1698175906
transform 1 0 9184 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_105_716
timestamp 1698175906
transform 1 0 17024 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_105_717
timestamp 1698175906
transform 1 0 24864 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_105_718
timestamp 1698175906
transform 1 0 32704 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_106_719
timestamp 1698175906
transform 1 0 5264 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_106_720
timestamp 1698175906
transform 1 0 13104 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_106_721
timestamp 1698175906
transform 1 0 20944 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_106_722
timestamp 1698175906
transform 1 0 28784 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_106_723
timestamp 1698175906
transform 1 0 36624 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_107_724
timestamp 1698175906
transform 1 0 9184 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_107_725
timestamp 1698175906
transform 1 0 17024 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_107_726
timestamp 1698175906
transform 1 0 24864 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_107_727
timestamp 1698175906
transform 1 0 32704 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_108_728
timestamp 1698175906
transform 1 0 5264 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_108_729
timestamp 1698175906
transform 1 0 13104 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_108_730
timestamp 1698175906
transform 1 0 20944 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_108_731
timestamp 1698175906
transform 1 0 28784 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_108_732
timestamp 1698175906
transform 1 0 36624 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_109_733
timestamp 1698175906
transform 1 0 9184 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_109_734
timestamp 1698175906
transform 1 0 17024 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_109_735
timestamp 1698175906
transform 1 0 24864 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_109_736
timestamp 1698175906
transform 1 0 32704 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_110_737
timestamp 1698175906
transform 1 0 5264 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_110_738
timestamp 1698175906
transform 1 0 13104 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_110_739
timestamp 1698175906
transform 1 0 20944 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_110_740
timestamp 1698175906
transform 1 0 28784 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_110_741
timestamp 1698175906
transform 1 0 36624 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_111_742
timestamp 1698175906
transform 1 0 9184 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_111_743
timestamp 1698175906
transform 1 0 17024 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_111_744
timestamp 1698175906
transform 1 0 24864 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_111_745
timestamp 1698175906
transform 1 0 32704 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_112_746
timestamp 1698175906
transform 1 0 5264 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_112_747
timestamp 1698175906
transform 1 0 13104 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_112_748
timestamp 1698175906
transform 1 0 20944 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_112_749
timestamp 1698175906
transform 1 0 28784 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_112_750
timestamp 1698175906
transform 1 0 36624 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_113_751
timestamp 1698175906
transform 1 0 9184 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_113_752
timestamp 1698175906
transform 1 0 17024 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_113_753
timestamp 1698175906
transform 1 0 24864 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_113_754
timestamp 1698175906
transform 1 0 32704 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_114_755
timestamp 1698175906
transform 1 0 5264 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_114_756
timestamp 1698175906
transform 1 0 13104 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_114_757
timestamp 1698175906
transform 1 0 20944 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_114_758
timestamp 1698175906
transform 1 0 28784 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_114_759
timestamp 1698175906
transform 1 0 36624 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_115_760
timestamp 1698175906
transform 1 0 9184 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_115_761
timestamp 1698175906
transform 1 0 17024 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_115_762
timestamp 1698175906
transform 1 0 24864 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_115_763
timestamp 1698175906
transform 1 0 32704 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_116_764
timestamp 1698175906
transform 1 0 5264 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_116_765
timestamp 1698175906
transform 1 0 13104 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_116_766
timestamp 1698175906
transform 1 0 20944 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_116_767
timestamp 1698175906
transform 1 0 28784 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_116_768
timestamp 1698175906
transform 1 0 36624 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_117_769
timestamp 1698175906
transform 1 0 9184 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_117_770
timestamp 1698175906
transform 1 0 17024 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_117_771
timestamp 1698175906
transform 1 0 24864 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_117_772
timestamp 1698175906
transform 1 0 32704 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_118_773
timestamp 1698175906
transform 1 0 5152 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_118_774
timestamp 1698175906
transform 1 0 8960 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_118_775
timestamp 1698175906
transform 1 0 12768 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_118_776
timestamp 1698175906
transform 1 0 16576 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_118_777
timestamp 1698175906
transform 1 0 20384 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_118_778
timestamp 1698175906
transform 1 0 24192 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_118_779
timestamp 1698175906
transform 1 0 28000 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_118_780
timestamp 1698175906
transform 1 0 31808 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_118_781
timestamp 1698175906
transform 1 0 35616 0 1 95648
box -86 -86 310 870
<< labels >>
flabel metal3 s 39200 30912 40000 31024 0 FreeSans 448 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 0 63840 800 63952 0 FreeSans 448 0 0 0 compare_in[0]
port 1 nsew signal input
flabel metal3 s 0 49056 800 49168 0 FreeSans 448 0 0 0 compare_in[10]
port 2 nsew signal input
flabel metal3 s 0 56448 800 56560 0 FreeSans 448 0 0 0 compare_in[11]
port 3 nsew signal input
flabel metal3 s 0 51744 800 51856 0 FreeSans 448 0 0 0 compare_in[12]
port 4 nsew signal input
flabel metal3 s 0 48384 800 48496 0 FreeSans 448 0 0 0 compare_in[13]
port 5 nsew signal input
flabel metal3 s 0 55776 800 55888 0 FreeSans 448 0 0 0 compare_in[14]
port 6 nsew signal input
flabel metal3 s 0 51072 800 51184 0 FreeSans 448 0 0 0 compare_in[15]
port 7 nsew signal input
flabel metal3 s 0 50400 800 50512 0 FreeSans 448 0 0 0 compare_in[16]
port 8 nsew signal input
flabel metal3 s 0 49728 800 49840 0 FreeSans 448 0 0 0 compare_in[17]
port 9 nsew signal input
flabel metal3 s 0 44352 800 44464 0 FreeSans 448 0 0 0 compare_in[18]
port 10 nsew signal input
flabel metal3 s 0 47712 800 47824 0 FreeSans 448 0 0 0 compare_in[19]
port 11 nsew signal input
flabel metal3 s 0 66528 800 66640 0 FreeSans 448 0 0 0 compare_in[1]
port 12 nsew signal input
flabel metal3 s 0 38976 800 39088 0 FreeSans 448 0 0 0 compare_in[20]
port 13 nsew signal input
flabel metal3 s 0 39648 800 39760 0 FreeSans 448 0 0 0 compare_in[21]
port 14 nsew signal input
flabel metal3 s 0 40320 800 40432 0 FreeSans 448 0 0 0 compare_in[22]
port 15 nsew signal input
flabel metal3 s 0 43680 800 43792 0 FreeSans 448 0 0 0 compare_in[23]
port 16 nsew signal input
flabel metal3 s 0 67872 800 67984 0 FreeSans 448 0 0 0 compare_in[2]
port 17 nsew signal input
flabel metal3 s 0 67200 800 67312 0 FreeSans 448 0 0 0 compare_in[3]
port 18 nsew signal input
flabel metal3 s 0 64512 800 64624 0 FreeSans 448 0 0 0 compare_in[4]
port 19 nsew signal input
flabel metal3 s 0 62496 800 62608 0 FreeSans 448 0 0 0 compare_in[5]
port 20 nsew signal input
flabel metal3 s 0 63168 800 63280 0 FreeSans 448 0 0 0 compare_in[6]
port 21 nsew signal input
flabel metal3 s 0 59136 800 59248 0 FreeSans 448 0 0 0 compare_in[7]
port 22 nsew signal input
flabel metal3 s 0 57120 800 57232 0 FreeSans 448 0 0 0 compare_in[8]
port 23 nsew signal input
flabel metal3 s 0 57792 800 57904 0 FreeSans 448 0 0 0 compare_in[9]
port 24 nsew signal input
flabel metal3 s 39200 30240 40000 30352 0 FreeSans 448 0 0 0 io_oeb[0]
port 25 nsew signal tristate
flabel metal2 s 2688 0 2800 800 0 FreeSans 448 90 0 0 io_oeb[1]
port 26 nsew signal tristate
flabel metal3 s 39200 63840 40000 63952 0 FreeSans 448 0 0 0 io_oeb[2]
port 27 nsew signal tristate
flabel metal3 s 39200 36288 40000 36400 0 FreeSans 448 0 0 0 io_oeb[3]
port 28 nsew signal tristate
flabel metal3 s 39200 22848 40000 22960 0 FreeSans 448 0 0 0 io_oeb[4]
port 29 nsew signal tristate
flabel metal2 s 3360 99200 3472 100000 0 FreeSans 448 90 0 0 io_oeb[5]
port 30 nsew signal tristate
flabel metal3 s 0 32928 800 33040 0 FreeSans 448 0 0 0 io_oeb[6]
port 31 nsew signal tristate
flabel metal3 s 39200 38976 40000 39088 0 FreeSans 448 0 0 0 led_out[0]
port 32 nsew signal tristate
flabel metal3 s 39200 53088 40000 53200 0 FreeSans 448 0 0 0 led_out[1]
port 33 nsew signal tristate
flabel metal3 s 39200 41664 40000 41776 0 FreeSans 448 0 0 0 led_out[2]
port 34 nsew signal tristate
flabel metal3 s 39200 42336 40000 42448 0 FreeSans 448 0 0 0 led_out[3]
port 35 nsew signal tristate
flabel metal3 s 39200 46368 40000 46480 0 FreeSans 448 0 0 0 led_out[4]
port 36 nsew signal tristate
flabel metal3 s 39200 47040 40000 47152 0 FreeSans 448 0 0 0 led_out[5]
port 37 nsew signal tristate
flabel metal3 s 39200 49728 40000 49840 0 FreeSans 448 0 0 0 led_out[6]
port 38 nsew signal tristate
flabel metal3 s 0 55104 800 55216 0 FreeSans 448 0 0 0 reset
port 39 nsew signal input
flabel metal3 s 0 53088 800 53200 0 FreeSans 448 0 0 0 update_compare
port 40 nsew signal input
flabel metal4 s 4448 3076 4768 96492 0 FreeSans 1280 90 0 0 vdd
port 41 nsew power bidirectional
flabel metal4 s 35168 3076 35488 96492 0 FreeSans 1280 90 0 0 vdd
port 41 nsew power bidirectional
flabel metal4 s 19808 3076 20128 96492 0 FreeSans 1280 90 0 0 vss
port 42 nsew ground bidirectional
rlabel metal1 19992 96432 19992 96432 0 vdd
rlabel via1 19992 95648 19992 95648 0 vss
rlabel metal2 34160 38920 34160 38920 0 _000_
rlabel metal2 34104 52416 34104 52416 0 _001_
rlabel metal2 34552 42056 34552 42056 0 _002_
rlabel metal3 34944 41832 34944 41832 0 _003_
rlabel metal2 36120 44912 36120 44912 0 _004_
rlabel metal2 36120 47208 36120 47208 0 _005_
rlabel metal2 35672 49392 35672 49392 0 _006_
rlabel metal2 31920 38136 31920 38136 0 _007_
rlabel metal2 32424 49392 32424 49392 0 _008_
rlabel metal2 33600 48328 33600 48328 0 _009_
rlabel metal2 33320 43120 33320 43120 0 _010_
rlabel metal2 14224 64456 14224 64456 0 _011_
rlabel metal2 11032 68208 11032 68208 0 _012_
rlabel metal2 11704 67200 11704 67200 0 _013_
rlabel metal2 9800 67480 9800 67480 0 _014_
rlabel metal2 10472 64344 10472 64344 0 _015_
rlabel metal3 9632 62216 9632 62216 0 _016_
rlabel metal2 14280 62776 14280 62776 0 _017_
rlabel metal2 12936 58632 12936 58632 0 _018_
rlabel metal2 12712 55608 12712 55608 0 _019_
rlabel metal2 8008 59640 8008 59640 0 _020_
rlabel metal2 7448 50904 7448 50904 0 _021_
rlabel metal3 8176 55944 8176 55944 0 _022_
rlabel metal2 12488 51688 12488 51688 0 _023_
rlabel metal3 6328 48440 6328 48440 0 _024_
rlabel metal3 7560 55160 7560 55160 0 _025_
rlabel metal2 12768 49896 12768 49896 0 _026_
rlabel metal2 10864 45976 10864 45976 0 _027_
rlabel metal2 10752 44408 10752 44408 0 _028_
rlabel metal3 6440 44856 6440 44856 0 _029_
rlabel metal2 7336 46256 7336 46256 0 _030_
rlabel metal2 9072 38136 9072 38136 0 _031_
rlabel metal2 8792 37016 8792 37016 0 _032_
rlabel metal2 11144 39256 11144 39256 0 _033_
rlabel metal2 8008 42392 8008 42392 0 _034_
rlabel metal2 24472 69720 24472 69720 0 _035_
rlabel metal2 23240 67872 23240 67872 0 _036_
rlabel metal3 27496 68488 27496 68488 0 _037_
rlabel metal2 26488 67424 26488 67424 0 _038_
rlabel metal2 23632 63000 23632 63000 0 _039_
rlabel metal2 27496 63504 27496 63504 0 _040_
rlabel metal2 26600 60256 26600 60256 0 _041_
rlabel metal2 23688 57960 23688 57960 0 _042_
rlabel metal2 27832 57344 27832 57344 0 _043_
rlabel metal2 27888 54600 27888 54600 0 _044_
rlabel metal2 26600 52584 26600 52584 0 _045_
rlabel metal2 25816 36120 25816 36120 0 _046_
rlabel metal2 26152 45920 26152 45920 0 _047_
rlabel metal2 27720 36008 27720 36008 0 _048_
rlabel metal2 27496 32872 27496 32872 0 _049_
rlabel metal2 21112 32928 21112 32928 0 _050_
rlabel metal2 25592 48272 25592 48272 0 _051_
rlabel metal2 18424 33208 18424 33208 0 _052_
rlabel metal2 17528 34440 17528 34440 0 _053_
rlabel metal3 12880 35112 12880 35112 0 _054_
rlabel metal2 12600 33768 12600 33768 0 _055_
rlabel metal2 12152 31360 12152 31360 0 _056_
rlabel metal2 22120 30520 22120 30520 0 _057_
rlabel metal2 25592 31248 25592 31248 0 _058_
rlabel metal2 10584 49000 10584 49000 0 _059_
rlabel metal3 30744 43512 30744 43512 0 _060_
rlabel metal2 29288 40880 29288 40880 0 _061_
rlabel metal2 29624 41888 29624 41888 0 _062_
rlabel metal2 16296 58912 16296 58912 0 _063_
rlabel metal2 15848 58744 15848 58744 0 _064_
rlabel metal2 17864 55944 17864 55944 0 _065_
rlabel metal2 18704 48440 18704 48440 0 _066_
rlabel metal2 15400 49952 15400 49952 0 _067_
rlabel metal2 15904 49896 15904 49896 0 _068_
rlabel metal2 16016 49000 16016 49000 0 _069_
rlabel metal2 17584 46648 17584 46648 0 _070_
rlabel metal2 14840 42336 14840 42336 0 _071_
rlabel metal2 14280 41384 14280 41384 0 _072_
rlabel metal2 21840 44408 21840 44408 0 _073_
rlabel metal2 22848 38024 22848 38024 0 _074_
rlabel metal3 14392 38920 14392 38920 0 _075_
rlabel metal2 16632 52976 16632 52976 0 _076_
rlabel metal2 17528 41776 17528 41776 0 _077_
rlabel metal2 14728 43148 14728 43148 0 _078_
rlabel metal2 14952 40600 14952 40600 0 _079_
rlabel metal2 15176 39088 15176 39088 0 _080_
rlabel metal2 13160 38304 13160 38304 0 _081_
rlabel metal2 22624 38584 22624 38584 0 _082_
rlabel metal2 22848 31192 22848 31192 0 _083_
rlabel metal2 24248 38304 24248 38304 0 _084_
rlabel metal2 24472 38472 24472 38472 0 _085_
rlabel metal4 24808 39648 24808 39648 0 _086_
rlabel metal2 18200 54040 18200 54040 0 _087_
rlabel metal3 16352 56616 16352 56616 0 _088_
rlabel metal2 17416 55944 17416 55944 0 _089_
rlabel metal2 17584 56280 17584 56280 0 _090_
rlabel metal3 19880 55384 19880 55384 0 _091_
rlabel metal2 22344 52472 22344 52472 0 _092_
rlabel metal2 17640 62272 17640 62272 0 _093_
rlabel metal2 21560 62832 21560 62832 0 _094_
rlabel metal2 18536 68096 18536 68096 0 _095_
rlabel metal2 17416 69440 17416 69440 0 _096_
rlabel metal2 18984 65408 18984 65408 0 _097_
rlabel metal2 20328 63392 20328 63392 0 _098_
rlabel metal2 20384 62888 20384 62888 0 _099_
rlabel metal3 17192 62440 17192 62440 0 _100_
rlabel metal2 18928 61432 18928 61432 0 _101_
rlabel metal2 17640 62552 17640 62552 0 _102_
rlabel metal3 20048 62104 20048 62104 0 _103_
rlabel metal3 19208 61544 19208 61544 0 _104_
rlabel metal2 20888 60872 20888 60872 0 _105_
rlabel metal2 19880 69888 19880 69888 0 _106_
rlabel metal2 17640 69104 17640 69104 0 _107_
rlabel metal2 20216 69104 20216 69104 0 _108_
rlabel metal2 20776 68236 20776 68236 0 _109_
rlabel metal2 21056 69944 21056 69944 0 _110_
rlabel metal2 19656 68544 19656 68544 0 _111_
rlabel metal2 20216 67760 20216 67760 0 _112_
rlabel metal2 19096 69664 19096 69664 0 _113_
rlabel metal2 20440 67928 20440 67928 0 _114_
rlabel metal2 21168 66808 21168 66808 0 _115_
rlabel metal3 23856 61320 23856 61320 0 _116_
rlabel metal2 18200 59696 18200 59696 0 _117_
rlabel metal2 19096 60760 19096 60760 0 _118_
rlabel metal2 19880 60424 19880 60424 0 _119_
rlabel metal2 19768 60088 19768 60088 0 _120_
rlabel metal2 21728 60536 21728 60536 0 _121_
rlabel metal2 17696 47320 17696 47320 0 _122_
rlabel metal2 18032 46648 18032 46648 0 _123_
rlabel metal2 14784 45640 14784 45640 0 _124_
rlabel metal2 15064 45528 15064 45528 0 _125_
rlabel metal3 14980 45304 14980 45304 0 _126_
rlabel via2 18760 44072 18760 44072 0 _127_
rlabel metal2 16184 42840 16184 42840 0 _128_
rlabel metal2 14168 43176 14168 43176 0 _129_
rlabel metal2 17528 45528 17528 45528 0 _130_
rlabel metal2 17080 45080 17080 45080 0 _131_
rlabel metal2 19768 43344 19768 43344 0 _132_
rlabel metal2 19992 45192 19992 45192 0 _133_
rlabel metal2 19992 53480 19992 53480 0 _134_
rlabel metal3 18984 53480 18984 53480 0 _135_
rlabel metal2 17976 51968 17976 51968 0 _136_
rlabel metal2 15512 52416 15512 52416 0 _137_
rlabel metal2 20776 51184 20776 51184 0 _138_
rlabel metal2 25704 46200 25704 46200 0 _139_
rlabel metal2 21952 46872 21952 46872 0 _140_
rlabel metal2 23576 50148 23576 50148 0 _141_
rlabel metal2 26936 54600 26936 54600 0 _142_
rlabel metal2 19320 54712 19320 54712 0 _143_
rlabel metal2 19432 53368 19432 53368 0 _144_
rlabel metal2 24248 52136 24248 52136 0 _145_
rlabel metal2 15512 47544 15512 47544 0 _146_
rlabel metal2 20328 48328 20328 48328 0 _147_
rlabel metal3 18592 47992 18592 47992 0 _148_
rlabel metal2 21448 48664 21448 48664 0 _149_
rlabel metal2 23128 35112 23128 35112 0 _150_
rlabel metal3 22120 51464 22120 51464 0 _151_
rlabel metal2 23352 50736 23352 50736 0 _152_
rlabel metal3 23632 49896 23632 49896 0 _153_
rlabel metal2 20776 53928 20776 53928 0 _154_
rlabel metal3 22232 49784 22232 49784 0 _155_
rlabel metal2 14280 59080 14280 59080 0 _156_
rlabel metal2 21448 57008 21448 57008 0 _157_
rlabel metal2 22344 55888 22344 55888 0 _158_
rlabel metal2 24024 51632 24024 51632 0 _159_
rlabel metal2 24136 42728 24136 42728 0 _160_
rlabel metal2 21448 41328 21448 41328 0 _161_
rlabel metal2 18256 36344 18256 36344 0 _162_
rlabel metal2 20664 42336 20664 42336 0 _163_
rlabel metal2 19880 42056 19880 42056 0 _164_
rlabel metal2 19992 41888 19992 41888 0 _165_
rlabel metal2 20440 43008 20440 43008 0 _166_
rlabel metal2 20216 43008 20216 43008 0 _167_
rlabel metal2 20104 37296 20104 37296 0 _168_
rlabel metal2 19320 47320 19320 47320 0 _169_
rlabel metal2 19544 44576 19544 44576 0 _170_
rlabel metal2 21056 42616 21056 42616 0 _171_
rlabel metal3 23744 41832 23744 41832 0 _172_
rlabel metal2 17752 37492 17752 37492 0 _173_
rlabel metal2 16016 46424 16016 46424 0 _174_
rlabel metal2 14056 41328 14056 41328 0 _175_
rlabel metal3 17304 38808 17304 38808 0 _176_
rlabel metal2 20664 38920 20664 38920 0 _177_
rlabel metal3 20048 38808 20048 38808 0 _178_
rlabel metal2 19264 38472 19264 38472 0 _179_
rlabel metal2 19656 39816 19656 39816 0 _180_
rlabel metal2 23072 41160 23072 41160 0 _181_
rlabel metal2 15624 51800 15624 51800 0 _182_
rlabel metal2 19096 49000 19096 49000 0 _183_
rlabel metal2 19264 49896 19264 49896 0 _184_
rlabel metal2 21896 40824 21896 40824 0 _185_
rlabel metal2 21560 40320 21560 40320 0 _186_
rlabel metal2 20664 45752 20664 45752 0 _187_
rlabel metal2 20216 39760 20216 39760 0 _188_
rlabel metal3 21392 40264 21392 40264 0 _189_
rlabel metal3 24472 38808 24472 38808 0 _190_
rlabel metal2 21672 47152 21672 47152 0 _191_
rlabel metal3 23240 42056 23240 42056 0 _192_
rlabel metal2 17528 53312 17528 53312 0 _193_
rlabel metal3 20272 40488 20272 40488 0 _194_
rlabel metal2 23744 40264 23744 40264 0 _195_
rlabel metal2 22792 39536 22792 39536 0 _196_
rlabel metal2 25928 41160 25928 41160 0 _197_
rlabel metal2 29400 41552 29400 41552 0 _198_
rlabel metal2 31528 40768 31528 40768 0 _199_
rlabel metal2 30632 41328 30632 41328 0 _200_
rlabel metal2 30632 42224 30632 42224 0 _201_
rlabel metal2 30632 43008 30632 43008 0 _202_
rlabel metal2 30240 42056 30240 42056 0 _203_
rlabel metal2 30072 40992 30072 40992 0 _204_
rlabel metal2 31976 41496 31976 41496 0 _205_
rlabel metal3 33152 46648 33152 46648 0 _206_
rlabel metal2 29960 47824 29960 47824 0 _207_
rlabel metal2 32648 42504 32648 42504 0 _208_
rlabel metal2 19544 60816 19544 60816 0 _209_
rlabel metal3 19768 45080 19768 45080 0 _210_
rlabel metal3 20888 43624 20888 43624 0 _211_
rlabel metal2 21560 44016 21560 44016 0 _212_
rlabel metal2 23072 53032 23072 53032 0 _213_
rlabel metal3 25816 62440 25816 62440 0 _214_
rlabel metal2 19936 62216 19936 62216 0 _215_
rlabel metal2 21896 43568 21896 43568 0 _216_
rlabel metal2 23240 43792 23240 43792 0 _217_
rlabel metal2 22792 56336 22792 56336 0 _218_
rlabel metal2 21448 43288 21448 43288 0 _219_
rlabel metal3 22288 39592 22288 39592 0 _220_
rlabel metal2 26824 43344 26824 43344 0 _221_
rlabel metal2 21672 41272 21672 41272 0 _222_
rlabel metal2 21896 36008 21896 36008 0 _223_
rlabel metal2 21336 37688 21336 37688 0 _224_
rlabel metal2 21672 38332 21672 38332 0 _225_
rlabel metal2 23688 43904 23688 43904 0 _226_
rlabel metal2 22232 49000 22232 49000 0 _227_
rlabel metal3 21952 48216 21952 48216 0 _228_
rlabel metal2 22568 48664 22568 48664 0 _229_
rlabel metal3 21784 47656 21784 47656 0 _230_
rlabel metal2 23800 46088 23800 46088 0 _231_
rlabel metal2 24920 45080 24920 45080 0 _232_
rlabel metal2 32312 42392 32312 42392 0 _233_
rlabel metal2 32200 45808 32200 45808 0 _234_
rlabel metal2 30296 43176 30296 43176 0 _235_
rlabel metal2 27832 41608 27832 41608 0 _236_
rlabel metal2 28280 42056 28280 42056 0 _237_
rlabel metal2 24360 43680 24360 43680 0 _238_
rlabel metal2 30912 45976 30912 45976 0 _239_
rlabel metal2 32424 45360 32424 45360 0 _240_
rlabel metal3 35280 49000 35280 49000 0 _241_
rlabel metal2 33208 45472 33208 45472 0 _242_
rlabel metal2 30688 47320 30688 47320 0 _243_
rlabel metal2 33096 42784 33096 42784 0 _244_
rlabel metal2 28728 41720 28728 41720 0 _245_
rlabel metal2 28728 42840 28728 42840 0 _246_
rlabel metal2 32984 41888 32984 41888 0 _247_
rlabel metal2 33432 42168 33432 42168 0 _248_
rlabel metal2 32648 47824 32648 47824 0 _249_
rlabel metal2 34328 47600 34328 47600 0 _250_
rlabel metal2 34664 45864 34664 45864 0 _251_
rlabel metal2 33376 50568 33376 50568 0 _252_
rlabel metal3 32480 46760 32480 46760 0 _253_
rlabel metal2 33544 50736 33544 50736 0 _254_
rlabel metal2 32984 51464 32984 51464 0 _255_
rlabel metal2 34384 42168 34384 42168 0 _256_
rlabel metal3 32536 40936 32536 40936 0 _257_
rlabel metal2 34888 44296 34888 44296 0 _258_
rlabel metal3 33264 48888 33264 48888 0 _259_
rlabel metal3 34216 48440 34216 48440 0 _260_
rlabel metal2 10584 54208 10584 54208 0 _261_
rlabel metal2 11648 49784 11648 49784 0 _262_
rlabel metal2 14168 63056 14168 63056 0 _263_
rlabel metal2 9912 63504 9912 63504 0 _264_
rlabel metal3 11088 46872 11088 46872 0 _265_
rlabel metal2 12376 57120 12376 57120 0 _266_
rlabel metal2 14504 64400 14504 64400 0 _267_
rlabel metal2 11200 49672 11200 49672 0 _268_
rlabel metal2 12600 66360 12600 66360 0 _269_
rlabel metal2 7672 48664 7672 48664 0 _270_
rlabel metal2 8232 39088 8232 39088 0 _271_
rlabel metal2 10248 66696 10248 66696 0 _272_
rlabel metal3 11928 67704 11928 67704 0 _273_
rlabel metal2 12152 67872 12152 67872 0 _274_
rlabel metal2 8344 67872 8344 67872 0 _275_
rlabel metal2 11816 68096 11816 68096 0 _276_
rlabel metal2 10360 56392 10360 56392 0 _277_
rlabel metal2 11368 64456 11368 64456 0 _278_
rlabel metal2 9128 66920 9128 66920 0 _279_
rlabel metal2 8624 67144 8624 67144 0 _280_
rlabel metal2 10976 64120 10976 64120 0 _281_
rlabel metal2 10248 63952 10248 63952 0 _282_
rlabel metal2 10136 61656 10136 61656 0 _283_
rlabel metal2 9128 62608 9128 62608 0 _284_
rlabel metal2 8568 56448 8568 56448 0 _285_
rlabel metal2 13720 62776 13720 62776 0 _286_
rlabel metal3 12600 58632 12600 58632 0 _287_
rlabel metal2 13608 59080 13608 59080 0 _288_
rlabel metal2 13440 56840 13440 56840 0 _289_
rlabel metal3 8848 59192 8848 59192 0 _290_
rlabel metal2 9744 49896 9744 49896 0 _291_
rlabel metal2 8120 58072 8120 58072 0 _292_
rlabel metal2 7168 44184 7168 44184 0 _293_
rlabel metal2 7616 49000 7616 49000 0 _294_
rlabel metal2 11536 48216 11536 48216 0 _295_
rlabel metal3 9520 45192 9520 45192 0 _296_
rlabel metal3 8680 50456 8680 50456 0 _297_
rlabel metal2 9688 46256 9688 46256 0 _298_
rlabel metal2 9072 54712 9072 54712 0 _299_
rlabel metal2 8176 54712 8176 54712 0 _300_
rlabel metal2 11816 52192 11816 52192 0 _301_
rlabel metal2 6888 48608 6888 48608 0 _302_
rlabel metal2 8680 49616 8680 49616 0 _303_
rlabel metal2 7056 48328 7056 48328 0 _304_
rlabel metal2 9352 55328 9352 55328 0 _305_
rlabel metal2 7896 56728 7896 56728 0 _306_
rlabel metal2 11704 50624 11704 50624 0 _307_
rlabel metal2 11368 48944 11368 48944 0 _308_
rlabel metal2 10584 45976 10584 45976 0 _309_
rlabel metal2 10136 47040 10136 47040 0 _310_
rlabel metal2 6776 44856 6776 44856 0 _311_
rlabel metal2 8344 44576 8344 44576 0 _312_
rlabel metal3 9128 46760 9128 46760 0 _313_
rlabel metal2 8344 46984 8344 46984 0 _314_
rlabel metal3 8624 38808 8624 38808 0 _315_
rlabel metal2 10416 42728 10416 42728 0 _316_
rlabel metal2 8456 39312 8456 39312 0 _317_
rlabel metal3 8792 38920 8792 38920 0 _318_
rlabel metal2 7560 38976 7560 38976 0 _319_
rlabel metal2 11312 38920 11312 38920 0 _320_
rlabel metal2 11480 39032 11480 39032 0 _321_
rlabel metal2 7896 43876 7896 43876 0 _322_
rlabel metal2 8344 42280 8344 42280 0 _323_
rlabel metal2 24696 67760 24696 67760 0 _324_
rlabel metal2 28056 43568 28056 43568 0 _325_
rlabel metal3 26040 36904 26040 36904 0 _326_
rlabel metal3 26936 70056 26936 70056 0 _327_
rlabel metal2 25256 62832 25256 62832 0 _328_
rlabel metal3 25536 64456 25536 64456 0 _329_
rlabel metal2 25816 68992 25816 68992 0 _330_
rlabel metal2 24248 67452 24248 67452 0 _331_
rlabel metal3 23464 65464 23464 65464 0 _332_
rlabel metal2 27160 51464 27160 51464 0 _333_
rlabel metal2 26208 31192 26208 31192 0 _334_
rlabel metal2 26488 66640 26488 66640 0 _335_
rlabel metal2 25872 68376 25872 68376 0 _336_
rlabel metal2 26600 64484 26600 64484 0 _337_
rlabel metal3 26544 67032 26544 67032 0 _338_
rlabel metal2 27272 67032 27272 67032 0 _339_
rlabel metal3 25480 63112 25480 63112 0 _340_
rlabel metal2 24696 63392 24696 63392 0 _341_
rlabel metal2 24136 63000 24136 63000 0 _342_
rlabel metal2 27104 63000 27104 63000 0 _343_
rlabel metal2 27160 60200 27160 60200 0 _344_
rlabel metal2 24808 58352 24808 58352 0 _345_
rlabel metal2 24360 61544 24360 61544 0 _346_
rlabel metal2 25368 60200 25368 60200 0 _347_
rlabel metal2 26040 59864 26040 59864 0 _348_
rlabel metal2 27384 55496 27384 55496 0 _349_
rlabel metal2 27384 56784 27384 56784 0 _350_
rlabel metal3 25648 56616 25648 56616 0 _351_
rlabel metal2 27272 57680 27272 57680 0 _352_
rlabel metal2 25368 55608 25368 55608 0 _353_
rlabel metal3 27944 56840 27944 56840 0 _354_
rlabel metal3 28840 55384 28840 55384 0 _355_
rlabel metal2 26936 52584 26936 52584 0 _356_
rlabel metal2 27664 52248 27664 52248 0 _357_
rlabel metal3 25088 34328 25088 34328 0 _358_
rlabel metal2 25704 36176 25704 36176 0 _359_
rlabel metal2 26096 38920 26096 38920 0 _360_
rlabel metal2 26264 43904 26264 43904 0 _361_
rlabel metal3 26824 38584 26824 38584 0 _362_
rlabel metal2 28000 37352 28000 37352 0 _363_
rlabel metal2 25368 35728 25368 35728 0 _364_
rlabel metal2 26040 33768 26040 33768 0 _365_
rlabel metal2 22344 34272 22344 34272 0 _366_
rlabel metal2 21728 33544 21728 33544 0 _367_
rlabel metal3 21448 34328 21448 34328 0 _368_
rlabel metal3 23856 35000 23856 35000 0 _369_
rlabel metal3 25032 48216 25032 48216 0 _370_
rlabel metal3 19656 33320 19656 33320 0 _371_
rlabel metal2 17192 33768 17192 33768 0 _372_
rlabel metal2 17640 34832 17640 34832 0 _373_
rlabel metal2 17360 34104 17360 34104 0 _374_
rlabel metal2 15288 35056 15288 35056 0 _375_
rlabel metal2 14840 34944 14840 34944 0 _376_
rlabel metal3 13944 34776 13944 34776 0 _377_
rlabel metal3 14616 33208 14616 33208 0 _378_
rlabel metal2 14392 33712 14392 33712 0 _379_
rlabel metal2 14728 32088 14728 32088 0 _380_
rlabel metal2 23240 32256 23240 32256 0 _381_
rlabel metal2 23296 31752 23296 31752 0 _382_
rlabel metal2 21896 31304 21896 31304 0 _383_
rlabel metal2 24248 31584 24248 31584 0 _384_
rlabel metal3 24976 30968 24976 30968 0 _385_
rlabel metal3 33138 30968 33138 30968 0 clk
rlabel metal3 21448 38136 21448 38136 0 clknet_0_clk
rlabel metal2 20776 31528 20776 31528 0 clknet_3_0__leaf_clk
rlabel metal3 6832 42728 6832 42728 0 clknet_3_1__leaf_clk
rlabel metal2 27664 36456 27664 36456 0 clknet_3_2__leaf_clk
rlabel metal2 28000 46648 28000 46648 0 clknet_3_3__leaf_clk
rlabel metal2 5600 49784 5600 49784 0 clknet_3_4__leaf_clk
rlabel metal2 9520 62328 9520 62328 0 clknet_3_5__leaf_clk
rlabel metal3 27832 53704 27832 53704 0 clknet_3_6__leaf_clk
rlabel metal2 25816 67984 25816 67984 0 clknet_3_7__leaf_clk
rlabel metal2 16632 68096 16632 68096 0 compare\[0\]
rlabel metal2 16968 53648 16968 53648 0 compare\[10\]
rlabel metal2 16408 53256 16408 53256 0 compare\[11\]
rlabel metal2 15736 50904 15736 50904 0 compare\[12\]
rlabel metal2 8232 49728 8232 49728 0 compare\[13\]
rlabel metal2 17752 50904 17752 50904 0 compare\[14\]
rlabel metal2 14840 49504 14840 49504 0 compare\[15\]
rlabel metal2 13888 45640 13888 45640 0 compare\[16\]
rlabel metal2 12936 44352 12936 44352 0 compare\[17\]
rlabel metal2 8232 43960 8232 43960 0 compare\[18\]
rlabel metal2 9464 45080 9464 45080 0 compare\[19\]
rlabel via2 15848 68488 15848 68488 0 compare\[1\]
rlabel metal2 13720 39872 13720 39872 0 compare\[20\]
rlabel metal2 12600 38976 12600 38976 0 compare\[21\]
rlabel metal2 13496 40432 13496 40432 0 compare\[22\]
rlabel metal2 10584 42784 10584 42784 0 compare\[23\]
rlabel metal2 13944 67536 13944 67536 0 compare\[2\]
rlabel metal2 16744 67816 16744 67816 0 compare\[3\]
rlabel metal2 16072 62664 16072 62664 0 compare\[4\]
rlabel metal2 13608 61432 13608 61432 0 compare\[5\]
rlabel metal3 17864 63000 17864 63000 0 compare\[6\]
rlabel metal2 15064 59472 15064 59472 0 compare\[7\]
rlabel metal2 15512 55048 15512 55048 0 compare\[8\]
rlabel metal2 17640 54096 17640 54096 0 compare\[9\]
rlabel metal2 1848 64288 1848 64288 0 compare_in[0]
rlabel metal2 1736 49448 1736 49448 0 compare_in[10]
rlabel metal2 1736 56616 1736 56616 0 compare_in[11]
rlabel metal2 1736 51968 1736 51968 0 compare_in[12]
rlabel metal2 1736 48664 1736 48664 0 compare_in[13]
rlabel metal2 1736 55944 1736 55944 0 compare_in[14]
rlabel metal2 1736 51240 1736 51240 0 compare_in[15]
rlabel metal3 1246 50456 1246 50456 0 compare_in[16]
rlabel metal2 2408 50120 2408 50120 0 compare_in[17]
rlabel metal2 1736 44744 1736 44744 0 compare_in[18]
rlabel metal2 1736 47992 1736 47992 0 compare_in[19]
rlabel metal2 1736 66808 1736 66808 0 compare_in[1]
rlabel metal2 1736 39256 1736 39256 0 compare_in[20]
rlabel metal2 1736 40040 1736 40040 0 compare_in[21]
rlabel metal2 1848 40768 1848 40768 0 compare_in[22]
rlabel metal2 1736 43960 1736 43960 0 compare_in[23]
rlabel metal2 1736 68264 1736 68264 0 compare_in[2]
rlabel metal2 1736 67480 1736 67480 0 compare_in[3]
rlabel metal3 1582 64568 1582 64568 0 compare_in[4]
rlabel metal2 1736 62776 1736 62776 0 compare_in[5]
rlabel metal2 1736 63560 1736 63560 0 compare_in[6]
rlabel metal2 1736 59528 1736 59528 0 compare_in[7]
rlabel metal2 1736 57400 1736 57400 0 compare_in[8]
rlabel metal2 1736 58072 1736 58072 0 compare_in[9]
rlabel metal3 37114 39032 37114 39032 0 led_out[0]
rlabel metal2 38024 53704 38024 53704 0 led_out[1]
rlabel metal3 37114 41720 37114 41720 0 led_out[2]
rlabel metal3 37338 42392 37338 42392 0 led_out[3]
rlabel metal3 37002 46424 37002 46424 0 led_out[4]
rlabel metal2 36904 47600 36904 47600 0 led_out[5]
rlabel metal3 38010 49784 38010 49784 0 led_out[6]
rlabel metal2 2184 63896 2184 63896 0 net1
rlabel metal2 6664 44744 6664 44744 0 net10
rlabel metal2 8008 47880 8008 47880 0 net11
rlabel metal2 9912 66696 9912 66696 0 net12
rlabel metal2 8120 39144 8120 39144 0 net13
rlabel metal2 2072 40040 2072 40040 0 net14
rlabel metal2 9688 40712 9688 40712 0 net15
rlabel metal3 4872 44072 4872 44072 0 net16
rlabel metal3 5880 68712 5880 68712 0 net17
rlabel metal2 2072 67480 2072 67480 0 net18
rlabel metal3 5712 64568 5712 64568 0 net19
rlabel metal2 7224 49448 7224 49448 0 net2
rlabel metal3 5488 63000 5488 63000 0 net20
rlabel metal2 2072 63896 2072 63896 0 net21
rlabel metal3 2716 59752 2716 59752 0 net22
rlabel metal3 7560 57736 7560 57736 0 net23
rlabel metal2 7784 57960 7784 57960 0 net24
rlabel metal2 2072 55216 2072 55216 0 net25
rlabel metal2 2184 52752 2184 52752 0 net26
rlabel metal2 36344 38360 36344 38360 0 net27
rlabel metal2 36008 53648 36008 53648 0 net28
rlabel metal2 38248 42840 38248 42840 0 net29
rlabel metal2 2184 56392 2184 56392 0 net3
rlabel metal2 36456 42280 36456 42280 0 net30
rlabel metal2 36456 45416 36456 45416 0 net31
rlabel metal2 38248 47376 38248 47376 0 net32
rlabel metal2 37800 50512 37800 50512 0 net33
rlabel metal2 38248 30688 38248 30688 0 net34
rlabel metal2 2744 2030 2744 2030 0 net35
rlabel metal2 38248 64176 38248 64176 0 net36
rlabel metal3 38738 36344 38738 36344 0 net37
rlabel metal2 38248 23072 38248 23072 0 net38
rlabel metal2 3528 95928 3528 95928 0 net39
rlabel metal2 2072 52080 2072 52080 0 net4
rlabel metal3 1246 32984 1246 32984 0 net40
rlabel metal2 15288 54152 15288 54152 0 net41
rlabel metal2 21896 54768 21896 54768 0 net42
rlabel metal2 15400 42672 15400 42672 0 net43
rlabel metal2 16744 57960 16744 57960 0 net44
rlabel metal2 23296 45192 23296 45192 0 net45
rlabel metal2 17976 63168 17976 63168 0 net46
rlabel metal2 26488 44016 26488 44016 0 net47
rlabel metal3 4368 48888 4368 48888 0 net5
rlabel metal2 7448 56504 7448 56504 0 net6
rlabel metal2 11480 51128 11480 51128 0 net7
rlabel metal2 11256 50120 11256 50120 0 net8
rlabel metal2 2744 50512 2744 50512 0 net9
rlabel metal3 1246 55160 1246 55160 0 reset
rlabel metal3 21392 69496 21392 69496 0 second_counter\[0\]
rlabel metal2 27384 53144 27384 53144 0 second_counter\[10\]
rlabel metal2 24696 37296 24696 37296 0 second_counter\[11\]
rlabel metal2 25256 46200 25256 46200 0 second_counter\[12\]
rlabel metal2 26488 37856 26488 37856 0 second_counter\[13\]
rlabel metal2 22680 36008 22680 36008 0 second_counter\[14\]
rlabel metal3 21168 34104 21168 34104 0 second_counter\[15\]
rlabel metal3 21504 48776 21504 48776 0 second_counter\[16\]
rlabel metal2 20216 33936 20216 33936 0 second_counter\[17\]
rlabel metal2 19208 35728 19208 35728 0 second_counter\[18\]
rlabel metal3 15736 35784 15736 35784 0 second_counter\[19\]
rlabel metal3 22736 68488 22736 68488 0 second_counter\[1\]
rlabel metal2 16296 35336 16296 35336 0 second_counter\[20\]
rlabel metal2 13776 38696 13776 38696 0 second_counter\[21\]
rlabel metal2 23240 30632 23240 30632 0 second_counter\[22\]
rlabel metal2 23464 31416 23464 31416 0 second_counter\[23\]
rlabel metal2 25256 68768 25256 68768 0 second_counter\[2\]
rlabel metal2 25816 66976 25816 66976 0 second_counter\[3\]
rlabel metal2 21448 63448 21448 63448 0 second_counter\[4\]
rlabel metal2 26264 63056 26264 63056 0 second_counter\[5\]
rlabel metal3 22064 61432 22064 61432 0 second_counter\[6\]
rlabel metal3 22288 56840 22288 56840 0 second_counter\[7\]
rlabel metal2 26936 56504 26936 56504 0 second_counter\[8\]
rlabel metal2 29960 54824 29960 54824 0 second_counter\[9\]
rlabel metal2 31864 41272 31864 41272 0 seg7.counter\[0\]
rlabel metal2 29288 46424 29288 46424 0 seg7.counter\[1\]
rlabel metal2 30744 43792 30744 43792 0 seg7.counter\[2\]
rlabel metal3 34048 40376 34048 40376 0 seg7.counter\[3\]
rlabel metal2 1736 53312 1736 53312 0 update_compare
<< properties >>
string FIXED_BBOX 0 0 40000 100000
<< end >>
