magic
tech gf180mcuD
magscale 1 5
timestamp 1700152634
<< obsm1 >>
rect 672 1538 9376 8262
<< metal2 >>
rect 3024 9600 3080 10000
rect 3360 9600 3416 10000
rect 3696 9600 3752 10000
rect 4032 9600 4088 10000
rect 4368 9600 4424 10000
rect 4704 9600 4760 10000
rect 5376 9600 5432 10000
rect 5712 9600 5768 10000
rect 6720 9600 6776 10000
rect 7056 9600 7112 10000
rect 7392 9600 7448 10000
rect 0 0 56 400
rect 336 0 392 400
rect 672 0 728 400
rect 1008 0 1064 400
rect 1344 0 1400 400
rect 1680 0 1736 400
rect 2016 0 2072 400
rect 2352 0 2408 400
rect 2688 0 2744 400
rect 3024 0 3080 400
rect 3360 0 3416 400
rect 3696 0 3752 400
rect 4032 0 4088 400
rect 4368 0 4424 400
rect 4704 0 4760 400
rect 5040 0 5096 400
rect 5376 0 5432 400
rect 5712 0 5768 400
rect 6048 0 6104 400
rect 6384 0 6440 400
rect 6720 0 6776 400
rect 7056 0 7112 400
rect 7392 0 7448 400
rect 7728 0 7784 400
rect 8064 0 8120 400
rect 8400 0 8456 400
rect 8736 0 8792 400
rect 9072 0 9128 400
rect 9408 0 9464 400
<< obsm2 >>
rect 14 9570 2994 9600
rect 3110 9570 3330 9600
rect 3446 9570 3666 9600
rect 3782 9570 4002 9600
rect 4118 9570 4338 9600
rect 4454 9570 4674 9600
rect 4790 9570 5346 9600
rect 5462 9570 5682 9600
rect 5798 9570 6690 9600
rect 6806 9570 7026 9600
rect 7142 9570 7362 9600
rect 7478 9570 9450 9600
rect 14 430 9450 9570
rect 86 400 306 430
rect 422 400 642 430
rect 758 400 978 430
rect 1094 400 1314 430
rect 1430 400 1650 430
rect 1766 400 1986 430
rect 2102 400 2322 430
rect 2438 400 2658 430
rect 2774 400 2994 430
rect 3110 400 3330 430
rect 3446 400 3666 430
rect 3782 400 4002 430
rect 4118 400 4338 430
rect 4454 400 4674 430
rect 4790 400 5010 430
rect 5126 400 5346 430
rect 5462 400 5682 430
rect 5798 400 6018 430
rect 6134 400 6354 430
rect 6470 400 6690 430
rect 6806 400 7026 430
rect 7142 400 7362 430
rect 7478 400 7698 430
rect 7814 400 8034 430
rect 8150 400 8370 430
rect 8486 400 8706 430
rect 8822 400 9042 430
rect 9158 400 9378 430
<< metal3 >>
rect 0 8400 400 8456
rect 0 8064 400 8120
rect 0 7728 400 7784
rect 9600 7728 10000 7784
rect 0 7392 400 7448
rect 9600 7392 10000 7448
rect 0 7056 400 7112
rect 9600 7056 10000 7112
rect 0 6720 400 6776
rect 0 6384 400 6440
rect 9600 6384 10000 6440
rect 0 6048 400 6104
rect 9600 6048 10000 6104
rect 0 5712 400 5768
rect 9600 5712 10000 5768
rect 0 5376 400 5432
rect 9600 5376 10000 5432
rect 0 5040 400 5096
rect 9600 5040 10000 5096
rect 0 4704 400 4760
rect 9600 4704 10000 4760
rect 0 4368 400 4424
rect 9600 4368 10000 4424
rect 0 4032 400 4088
rect 9600 4032 10000 4088
rect 0 3696 400 3752
rect 9600 3696 10000 3752
rect 0 3360 400 3416
rect 0 3024 400 3080
rect 9600 3024 10000 3080
rect 0 2688 400 2744
rect 0 2352 400 2408
rect 0 2016 400 2072
rect 9600 2016 10000 2072
rect 0 1680 400 1736
rect 0 1344 400 1400
rect 0 1008 400 1064
<< obsm3 >>
rect 430 8370 9600 8442
rect 9 8150 9600 8370
rect 430 8034 9600 8150
rect 9 7814 9600 8034
rect 430 7698 9570 7814
rect 9 7478 9600 7698
rect 430 7362 9570 7478
rect 9 7142 9600 7362
rect 430 7026 9570 7142
rect 9 6806 9600 7026
rect 430 6690 9600 6806
rect 9 6470 9600 6690
rect 430 6354 9570 6470
rect 9 6134 9600 6354
rect 430 6018 9570 6134
rect 9 5798 9600 6018
rect 430 5682 9570 5798
rect 9 5462 9600 5682
rect 430 5346 9570 5462
rect 9 5126 9600 5346
rect 430 5010 9570 5126
rect 9 4790 9600 5010
rect 430 4674 9570 4790
rect 9 4454 9600 4674
rect 430 4338 9570 4454
rect 9 4118 9600 4338
rect 430 4002 9570 4118
rect 9 3782 9600 4002
rect 430 3666 9570 3782
rect 9 3446 9600 3666
rect 430 3330 9600 3446
rect 9 3110 9600 3330
rect 430 2994 9570 3110
rect 9 2774 9600 2994
rect 430 2658 9600 2774
rect 9 2438 9600 2658
rect 430 2322 9600 2438
rect 9 2102 9600 2322
rect 430 1986 9570 2102
rect 9 1766 9600 1986
rect 430 1650 9600 1766
rect 9 1430 9600 1650
rect 430 1314 9600 1430
rect 9 1094 9600 1314
rect 430 1022 9600 1094
<< metal4 >>
rect 1670 1538 1830 8262
rect 2748 1538 2908 8262
rect 3826 1538 3986 8262
rect 4904 1538 5064 8262
rect 5982 1538 6142 8262
rect 7060 1538 7220 8262
rect 8138 1538 8298 8262
rect 9216 1538 9376 8262
<< labels >>
rlabel metal4 s 1670 1538 1830 8262 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 3826 1538 3986 8262 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 5982 1538 6142 8262 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 8138 1538 8298 8262 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 2748 1538 2908 8262 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 4904 1538 5064 8262 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 7060 1538 7220 8262 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 9216 1538 9376 8262 6 VSS
port 2 nsew ground bidirectional
rlabel metal3 s 9600 5712 10000 5768 6 buttons[0]
port 3 nsew signal input
rlabel metal3 s 9600 4704 10000 4760 6 buttons[1]
port 4 nsew signal input
rlabel metal3 s 0 6720 400 6776 6 clk
port 5 nsew signal input
rlabel metal2 s 0 0 56 400 6 i_wb_addr[0]
port 6 nsew signal input
rlabel metal2 s 336 0 392 400 6 i_wb_addr[10]
port 7 nsew signal input
rlabel metal2 s 9408 0 9464 400 6 i_wb_addr[11]
port 8 nsew signal input
rlabel metal2 s 9072 0 9128 400 6 i_wb_addr[12]
port 9 nsew signal input
rlabel metal2 s 5376 0 5432 400 6 i_wb_addr[13]
port 10 nsew signal input
rlabel metal2 s 4368 0 4424 400 6 i_wb_addr[14]
port 11 nsew signal input
rlabel metal2 s 8400 0 8456 400 6 i_wb_addr[15]
port 12 nsew signal input
rlabel metal2 s 8736 0 8792 400 6 i_wb_addr[16]
port 13 nsew signal input
rlabel metal2 s 7728 0 7784 400 6 i_wb_addr[17]
port 14 nsew signal input
rlabel metal2 s 6720 0 6776 400 6 i_wb_addr[18]
port 15 nsew signal input
rlabel metal2 s 6384 0 6440 400 6 i_wb_addr[19]
port 16 nsew signal input
rlabel metal2 s 1344 0 1400 400 6 i_wb_addr[1]
port 17 nsew signal input
rlabel metal2 s 7392 0 7448 400 6 i_wb_addr[20]
port 18 nsew signal input
rlabel metal2 s 7056 0 7112 400 6 i_wb_addr[21]
port 19 nsew signal input
rlabel metal2 s 8064 0 8120 400 6 i_wb_addr[22]
port 20 nsew signal input
rlabel metal2 s 6048 0 6104 400 6 i_wb_addr[23]
port 21 nsew signal input
rlabel metal3 s 0 4368 400 4424 6 i_wb_addr[24]
port 22 nsew signal input
rlabel metal3 s 0 4032 400 4088 6 i_wb_addr[25]
port 23 nsew signal input
rlabel metal3 s 0 2352 400 2408 6 i_wb_addr[26]
port 24 nsew signal input
rlabel metal3 s 0 4704 400 4760 6 i_wb_addr[27]
port 25 nsew signal input
rlabel metal3 s 0 2688 400 2744 6 i_wb_addr[28]
port 26 nsew signal input
rlabel metal3 s 0 3696 400 3752 6 i_wb_addr[29]
port 27 nsew signal input
rlabel metal2 s 1680 0 1736 400 6 i_wb_addr[2]
port 28 nsew signal input
rlabel metal3 s 0 3360 400 3416 6 i_wb_addr[30]
port 29 nsew signal input
rlabel metal3 s 0 3024 400 3080 6 i_wb_addr[31]
port 30 nsew signal input
rlabel metal2 s 3360 0 3416 400 6 i_wb_addr[3]
port 31 nsew signal input
rlabel metal2 s 672 0 728 400 6 i_wb_addr[4]
port 32 nsew signal input
rlabel metal2 s 4032 0 4088 400 6 i_wb_addr[5]
port 33 nsew signal input
rlabel metal2 s 1008 0 1064 400 6 i_wb_addr[6]
port 34 nsew signal input
rlabel metal2 s 3696 0 3752 400 6 i_wb_addr[7]
port 35 nsew signal input
rlabel metal2 s 4704 0 4760 400 6 i_wb_addr[8]
port 36 nsew signal input
rlabel metal2 s 5040 0 5096 400 6 i_wb_addr[9]
port 37 nsew signal input
rlabel metal3 s 9600 3696 10000 3752 6 i_wb_cyc
port 38 nsew signal input
rlabel metal3 s 0 6384 400 6440 6 i_wb_data[0]
port 39 nsew signal input
rlabel metal3 s 0 5040 400 5096 6 i_wb_data[1]
port 40 nsew signal input
rlabel metal3 s 9600 4032 10000 4088 6 i_wb_stb
port 41 nsew signal input
rlabel metal3 s 9600 4368 10000 4424 6 i_wb_we
port 42 nsew signal input
rlabel metal2 s 4032 9600 4088 10000 6 leds[0]
port 43 nsew signal output
rlabel metal3 s 0 5376 400 5432 6 leds[1]
port 44 nsew signal output
rlabel metal3 s 9600 5376 10000 5432 6 o_wb_ack
port 45 nsew signal output
rlabel metal3 s 9600 6384 10000 6440 6 o_wb_data[0]
port 46 nsew signal output
rlabel metal2 s 2016 0 2072 400 6 o_wb_data[10]
port 47 nsew signal output
rlabel metal3 s 0 6048 400 6104 6 o_wb_data[11]
port 48 nsew signal output
rlabel metal3 s 0 1008 400 1064 6 o_wb_data[12]
port 49 nsew signal output
rlabel metal3 s 9600 2016 10000 2072 6 o_wb_data[13]
port 50 nsew signal output
rlabel metal2 s 4704 9600 4760 10000 6 o_wb_data[14]
port 51 nsew signal output
rlabel metal3 s 0 8400 400 8456 6 o_wb_data[15]
port 52 nsew signal output
rlabel metal2 s 3024 9600 3080 10000 6 o_wb_data[16]
port 53 nsew signal output
rlabel metal2 s 3696 9600 3752 10000 6 o_wb_data[17]
port 54 nsew signal output
rlabel metal3 s 0 7392 400 7448 6 o_wb_data[18]
port 55 nsew signal output
rlabel metal2 s 3024 0 3080 400 6 o_wb_data[19]
port 56 nsew signal output
rlabel metal3 s 9600 6048 10000 6104 6 o_wb_data[1]
port 57 nsew signal output
rlabel metal3 s 9600 3024 10000 3080 6 o_wb_data[20]
port 58 nsew signal output
rlabel metal2 s 2352 0 2408 400 6 o_wb_data[21]
port 59 nsew signal output
rlabel metal3 s 9600 7728 10000 7784 6 o_wb_data[22]
port 60 nsew signal output
rlabel metal2 s 7392 9600 7448 10000 6 o_wb_data[23]
port 61 nsew signal output
rlabel metal3 s 0 7728 400 7784 6 o_wb_data[24]
port 62 nsew signal output
rlabel metal2 s 3360 9600 3416 10000 6 o_wb_data[25]
port 63 nsew signal output
rlabel metal3 s 9600 7392 10000 7448 6 o_wb_data[26]
port 64 nsew signal output
rlabel metal3 s 0 1344 400 1400 6 o_wb_data[27]
port 65 nsew signal output
rlabel metal2 s 5712 0 5768 400 6 o_wb_data[28]
port 66 nsew signal output
rlabel metal3 s 0 1680 400 1736 6 o_wb_data[29]
port 67 nsew signal output
rlabel metal2 s 2688 0 2744 400 6 o_wb_data[2]
port 68 nsew signal output
rlabel metal3 s 9600 7056 10000 7112 6 o_wb_data[30]
port 69 nsew signal output
rlabel metal3 s 0 2016 400 2072 6 o_wb_data[31]
port 70 nsew signal output
rlabel metal2 s 5376 9600 5432 10000 6 o_wb_data[3]
port 71 nsew signal output
rlabel metal2 s 6720 9600 6776 10000 6 o_wb_data[4]
port 72 nsew signal output
rlabel metal2 s 7056 9600 7112 10000 6 o_wb_data[5]
port 73 nsew signal output
rlabel metal3 s 0 5712 400 5768 6 o_wb_data[6]
port 74 nsew signal output
rlabel metal3 s 0 8064 400 8120 6 o_wb_data[7]
port 75 nsew signal output
rlabel metal3 s 0 7056 400 7112 6 o_wb_data[8]
port 76 nsew signal output
rlabel metal2 s 5712 9600 5768 10000 6 o_wb_data[9]
port 77 nsew signal output
rlabel metal2 s 4368 9600 4424 10000 6 o_wb_stall
port 78 nsew signal output
rlabel metal3 s 9600 5040 10000 5096 6 reset
port 79 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 10000 10000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 367704
string GDS_FILE /home/farag/carvel_riscv_soc/gf180mcu_riscv_soc/openlane/wb_buttons_leds/runs/23_11_16_18_34/results/signoff/wb_buttons_leds.magic.gds
string GDS_START 139434
<< end >>

