VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DSM_core
  CLASS BLOCK ;
  FOREIGN DSM_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 200.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 198.000 49.280 200.000 49.840 ;
    END
  END clk
  PIN i_wb_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 21.280 2.000 21.840 ;
    END
  END i_wb_addr[0]
  PIN i_wb_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 97.440 2.000 98.000 ;
    END
  END i_wb_addr[10]
  PIN i_wb_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 101.920 2.000 102.480 ;
    END
  END i_wb_addr[11]
  PIN i_wb_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 106.400 2.000 106.960 ;
    END
  END i_wb_addr[12]
  PIN i_wb_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 110.880 2.000 111.440 ;
    END
  END i_wb_addr[13]
  PIN i_wb_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 115.360 2.000 115.920 ;
    END
  END i_wb_addr[14]
  PIN i_wb_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 119.840 2.000 120.400 ;
    END
  END i_wb_addr[15]
  PIN i_wb_addr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 124.320 2.000 124.880 ;
    END
  END i_wb_addr[16]
  PIN i_wb_addr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 128.800 2.000 129.360 ;
    END
  END i_wb_addr[17]
  PIN i_wb_addr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 133.280 2.000 133.840 ;
    END
  END i_wb_addr[18]
  PIN i_wb_addr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 137.760 2.000 138.320 ;
    END
  END i_wb_addr[19]
  PIN i_wb_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 30.240 2.000 30.800 ;
    END
  END i_wb_addr[1]
  PIN i_wb_addr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 142.240 2.000 142.800 ;
    END
  END i_wb_addr[20]
  PIN i_wb_addr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 146.720 2.000 147.280 ;
    END
  END i_wb_addr[21]
  PIN i_wb_addr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 151.200 2.000 151.760 ;
    END
  END i_wb_addr[22]
  PIN i_wb_addr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 155.680 2.000 156.240 ;
    END
  END i_wb_addr[23]
  PIN i_wb_addr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 160.160 2.000 160.720 ;
    END
  END i_wb_addr[24]
  PIN i_wb_addr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 164.640 2.000 165.200 ;
    END
  END i_wb_addr[25]
  PIN i_wb_addr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 169.120 2.000 169.680 ;
    END
  END i_wb_addr[26]
  PIN i_wb_addr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 173.600 2.000 174.160 ;
    END
  END i_wb_addr[27]
  PIN i_wb_addr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 178.080 2.000 178.640 ;
    END
  END i_wb_addr[28]
  PIN i_wb_addr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 182.560 2.000 183.120 ;
    END
  END i_wb_addr[29]
  PIN i_wb_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 39.200 2.000 39.760 ;
    END
  END i_wb_addr[2]
  PIN i_wb_addr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 187.040 2.000 187.600 ;
    END
  END i_wb_addr[30]
  PIN i_wb_addr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 191.520 2.000 192.080 ;
    END
  END i_wb_addr[31]
  PIN i_wb_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 48.160 2.000 48.720 ;
    END
  END i_wb_addr[3]
  PIN i_wb_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 57.120 2.000 57.680 ;
    END
  END i_wb_addr[4]
  PIN i_wb_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 66.080 2.000 66.640 ;
    END
  END i_wb_addr[5]
  PIN i_wb_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 75.040 2.000 75.600 ;
    END
  END i_wb_addr[6]
  PIN i_wb_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 84.000 2.000 84.560 ;
    END
  END i_wb_addr[7]
  PIN i_wb_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 88.480 2.000 89.040 ;
    END
  END i_wb_addr[8]
  PIN i_wb_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 92.960 2.000 93.520 ;
    END
  END i_wb_addr[9]
  PIN i_wb_cyc
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 7.840 2.000 8.400 ;
    END
  END i_wb_cyc
  PIN i_wb_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 25.760 2.000 26.320 ;
    END
  END i_wb_data[0]
  PIN i_wb_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 34.720 2.000 35.280 ;
    END
  END i_wb_data[1]
  PIN i_wb_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 43.680 2.000 44.240 ;
    END
  END i_wb_data[2]
  PIN i_wb_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 52.640 2.000 53.200 ;
    END
  END i_wb_data[3]
  PIN i_wb_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 61.600 2.000 62.160 ;
    END
  END i_wb_data[4]
  PIN i_wb_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 70.560 2.000 71.120 ;
    END
  END i_wb_data[5]
  PIN i_wb_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 79.520 2.000 80.080 ;
    END
  END i_wb_data[6]
  PIN i_wb_stb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 12.320 2.000 12.880 ;
    END
  END i_wb_stb
  PIN i_wb_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 16.800 2.000 17.360 ;
    END
  END i_wb_we
  PIN o_wb_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.604400 ;
    PORT
      LAYER Metal2 ;
        RECT 15.680 0.000 16.240 2.000 ;
    END
  END o_wb_ack
  PIN o_wb_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 2.604400 ;
    PORT
      LAYER Metal2 ;
        RECT 71.680 0.000 72.240 2.000 ;
    END
  END o_wb_data[0]
  PIN o_wb_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 2.604400 ;
    PORT
      LAYER Metal2 ;
        RECT 99.680 0.000 100.240 2.000 ;
    END
  END o_wb_data[1]
  PIN o_wb_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 2.604400 ;
    PORT
      LAYER Metal2 ;
        RECT 127.680 0.000 128.240 2.000 ;
    END
  END o_wb_data[2]
  PIN o_wb_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 2.604400 ;
    PORT
      LAYER Metal2 ;
        RECT 155.680 0.000 156.240 2.000 ;
    END
  END o_wb_data[3]
  PIN o_wb_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 2.604400 ;
    PORT
      LAYER Metal2 ;
        RECT 183.680 0.000 184.240 2.000 ;
    END
  END o_wb_data[4]
  PIN o_wb_stall
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 43.680 0.000 44.240 2.000 ;
    END
  END o_wb_stall
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 198.000 148.960 200.000 149.520 ;
    END
  END reset
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 7.540 23.840 192.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 7.540 177.440 192.380 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 7.540 100.640 192.380 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 7.540 193.200 192.380 ;
      LAYER Metal2 ;
        RECT 7.980 2.300 191.940 192.270 ;
        RECT 7.980 1.260 15.380 2.300 ;
        RECT 16.540 1.260 43.380 2.300 ;
        RECT 44.540 1.260 71.380 2.300 ;
        RECT 72.540 1.260 99.380 2.300 ;
        RECT 100.540 1.260 127.380 2.300 ;
        RECT 128.540 1.260 155.380 2.300 ;
        RECT 156.540 1.260 183.380 2.300 ;
        RECT 184.540 1.260 191.940 2.300 ;
      LAYER Metal3 ;
        RECT 2.300 191.220 198.000 192.220 ;
        RECT 2.000 187.900 198.000 191.220 ;
        RECT 2.300 186.740 198.000 187.900 ;
        RECT 2.000 183.420 198.000 186.740 ;
        RECT 2.300 182.260 198.000 183.420 ;
        RECT 2.000 178.940 198.000 182.260 ;
        RECT 2.300 177.780 198.000 178.940 ;
        RECT 2.000 174.460 198.000 177.780 ;
        RECT 2.300 173.300 198.000 174.460 ;
        RECT 2.000 169.980 198.000 173.300 ;
        RECT 2.300 168.820 198.000 169.980 ;
        RECT 2.000 165.500 198.000 168.820 ;
        RECT 2.300 164.340 198.000 165.500 ;
        RECT 2.000 161.020 198.000 164.340 ;
        RECT 2.300 159.860 198.000 161.020 ;
        RECT 2.000 156.540 198.000 159.860 ;
        RECT 2.300 155.380 198.000 156.540 ;
        RECT 2.000 152.060 198.000 155.380 ;
        RECT 2.300 150.900 198.000 152.060 ;
        RECT 2.000 149.820 198.000 150.900 ;
        RECT 2.000 148.660 197.700 149.820 ;
        RECT 2.000 147.580 198.000 148.660 ;
        RECT 2.300 146.420 198.000 147.580 ;
        RECT 2.000 143.100 198.000 146.420 ;
        RECT 2.300 141.940 198.000 143.100 ;
        RECT 2.000 138.620 198.000 141.940 ;
        RECT 2.300 137.460 198.000 138.620 ;
        RECT 2.000 134.140 198.000 137.460 ;
        RECT 2.300 132.980 198.000 134.140 ;
        RECT 2.000 129.660 198.000 132.980 ;
        RECT 2.300 128.500 198.000 129.660 ;
        RECT 2.000 125.180 198.000 128.500 ;
        RECT 2.300 124.020 198.000 125.180 ;
        RECT 2.000 120.700 198.000 124.020 ;
        RECT 2.300 119.540 198.000 120.700 ;
        RECT 2.000 116.220 198.000 119.540 ;
        RECT 2.300 115.060 198.000 116.220 ;
        RECT 2.000 111.740 198.000 115.060 ;
        RECT 2.300 110.580 198.000 111.740 ;
        RECT 2.000 107.260 198.000 110.580 ;
        RECT 2.300 106.100 198.000 107.260 ;
        RECT 2.000 102.780 198.000 106.100 ;
        RECT 2.300 101.620 198.000 102.780 ;
        RECT 2.000 98.300 198.000 101.620 ;
        RECT 2.300 97.140 198.000 98.300 ;
        RECT 2.000 93.820 198.000 97.140 ;
        RECT 2.300 92.660 198.000 93.820 ;
        RECT 2.000 89.340 198.000 92.660 ;
        RECT 2.300 88.180 198.000 89.340 ;
        RECT 2.000 84.860 198.000 88.180 ;
        RECT 2.300 83.700 198.000 84.860 ;
        RECT 2.000 80.380 198.000 83.700 ;
        RECT 2.300 79.220 198.000 80.380 ;
        RECT 2.000 75.900 198.000 79.220 ;
        RECT 2.300 74.740 198.000 75.900 ;
        RECT 2.000 71.420 198.000 74.740 ;
        RECT 2.300 70.260 198.000 71.420 ;
        RECT 2.000 66.940 198.000 70.260 ;
        RECT 2.300 65.780 198.000 66.940 ;
        RECT 2.000 62.460 198.000 65.780 ;
        RECT 2.300 61.300 198.000 62.460 ;
        RECT 2.000 57.980 198.000 61.300 ;
        RECT 2.300 56.820 198.000 57.980 ;
        RECT 2.000 53.500 198.000 56.820 ;
        RECT 2.300 52.340 198.000 53.500 ;
        RECT 2.000 50.140 198.000 52.340 ;
        RECT 2.000 49.020 197.700 50.140 ;
        RECT 2.300 48.980 197.700 49.020 ;
        RECT 2.300 47.860 198.000 48.980 ;
        RECT 2.000 44.540 198.000 47.860 ;
        RECT 2.300 43.380 198.000 44.540 ;
        RECT 2.000 40.060 198.000 43.380 ;
        RECT 2.300 38.900 198.000 40.060 ;
        RECT 2.000 35.580 198.000 38.900 ;
        RECT 2.300 34.420 198.000 35.580 ;
        RECT 2.000 31.100 198.000 34.420 ;
        RECT 2.300 29.940 198.000 31.100 ;
        RECT 2.000 26.620 198.000 29.940 ;
        RECT 2.300 25.460 198.000 26.620 ;
        RECT 2.000 22.140 198.000 25.460 ;
        RECT 2.300 20.980 198.000 22.140 ;
        RECT 2.000 17.660 198.000 20.980 ;
        RECT 2.300 16.500 198.000 17.660 ;
        RECT 2.000 13.180 198.000 16.500 ;
        RECT 2.300 12.020 198.000 13.180 ;
        RECT 2.000 8.700 198.000 12.020 ;
        RECT 2.300 7.700 198.000 8.700 ;
      LAYER Metal4 ;
        RECT 21.420 81.290 21.700 87.830 ;
  END
END DSM_core
END LIBRARY

