VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO riscv_top
  CLASS BLOCK ;
  FOREIGN riscv_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 500.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 154.560 200.000 155.120 ;
    END
  END clk
  PIN compare_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 319.200 4.000 319.760 ;
    END
  END compare_in[0]
  PIN compare_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 245.280 4.000 245.840 ;
    END
  END compare_in[10]
  PIN compare_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 282.240 4.000 282.800 ;
    END
  END compare_in[11]
  PIN compare_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 258.720 4.000 259.280 ;
    END
  END compare_in[12]
  PIN compare_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 241.920 4.000 242.480 ;
    END
  END compare_in[13]
  PIN compare_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 278.880 4.000 279.440 ;
    END
  END compare_in[14]
  PIN compare_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 255.360 4.000 255.920 ;
    END
  END compare_in[15]
  PIN compare_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 252.000 4.000 252.560 ;
    END
  END compare_in[16]
  PIN compare_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 248.640 4.000 249.200 ;
    END
  END compare_in[17]
  PIN compare_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 221.760 4.000 222.320 ;
    END
  END compare_in[18]
  PIN compare_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 238.560 4.000 239.120 ;
    END
  END compare_in[19]
  PIN compare_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 332.640 4.000 333.200 ;
    END
  END compare_in[1]
  PIN compare_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 194.880 4.000 195.440 ;
    END
  END compare_in[20]
  PIN compare_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 198.240 4.000 198.800 ;
    END
  END compare_in[21]
  PIN compare_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 201.600 4.000 202.160 ;
    END
  END compare_in[22]
  PIN compare_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 218.400 4.000 218.960 ;
    END
  END compare_in[23]
  PIN compare_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 339.360 4.000 339.920 ;
    END
  END compare_in[2]
  PIN compare_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 336.000 4.000 336.560 ;
    END
  END compare_in[3]
  PIN compare_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 322.560 4.000 323.120 ;
    END
  END compare_in[4]
  PIN compare_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 312.480 4.000 313.040 ;
    END
  END compare_in[5]
  PIN compare_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 315.840 4.000 316.400 ;
    END
  END compare_in[6]
  PIN compare_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 295.680 4.000 296.240 ;
    END
  END compare_in[7]
  PIN compare_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 285.600 4.000 286.160 ;
    END
  END compare_in[8]
  PIN compare_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 288.960 4.000 289.520 ;
    END
  END compare_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 151.200 200.000 151.760 ;
    END
  END io_oeb[0]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 13.440 0.000 14.000 4.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 319.200 200.000 319.760 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 181.440 200.000 182.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 114.240 200.000 114.800 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 16.800 496.000 17.360 500.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 164.640 4.000 165.200 ;
    END
  END io_oeb[6]
  PIN led_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 194.880 200.000 195.440 ;
    END
  END led_out[0]
  PIN led_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 265.440 200.000 266.000 ;
    END
  END led_out[1]
  PIN led_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 208.320 200.000 208.880 ;
    END
  END led_out[2]
  PIN led_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 211.680 200.000 212.240 ;
    END
  END led_out[3]
  PIN led_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 231.840 200.000 232.400 ;
    END
  END led_out[4]
  PIN led_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 235.200 200.000 235.760 ;
    END
  END led_out[5]
  PIN led_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 196.000 248.640 200.000 249.200 ;
    END
  END led_out[6]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 275.520 4.000 276.080 ;
    END
  END reset
  PIN update_compare
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 265.440 4.000 266.000 ;
    END
  END update_compare
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 482.460 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 482.460 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 482.460 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 193.200 482.460 ;
      LAYER Metal2 ;
        RECT 8.540 495.700 16.500 496.000 ;
        RECT 17.660 495.700 191.380 496.000 ;
        RECT 8.540 4.300 191.380 495.700 ;
        RECT 8.540 4.000 13.140 4.300 ;
        RECT 14.300 4.000 191.380 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 340.220 196.000 482.300 ;
        RECT 4.300 339.060 196.000 340.220 ;
        RECT 4.000 336.860 196.000 339.060 ;
        RECT 4.300 335.700 196.000 336.860 ;
        RECT 4.000 333.500 196.000 335.700 ;
        RECT 4.300 332.340 196.000 333.500 ;
        RECT 4.000 323.420 196.000 332.340 ;
        RECT 4.300 322.260 196.000 323.420 ;
        RECT 4.000 320.060 196.000 322.260 ;
        RECT 4.300 318.900 195.700 320.060 ;
        RECT 4.000 316.700 196.000 318.900 ;
        RECT 4.300 315.540 196.000 316.700 ;
        RECT 4.000 313.340 196.000 315.540 ;
        RECT 4.300 312.180 196.000 313.340 ;
        RECT 4.000 296.540 196.000 312.180 ;
        RECT 4.300 295.380 196.000 296.540 ;
        RECT 4.000 289.820 196.000 295.380 ;
        RECT 4.300 288.660 196.000 289.820 ;
        RECT 4.000 286.460 196.000 288.660 ;
        RECT 4.300 285.300 196.000 286.460 ;
        RECT 4.000 283.100 196.000 285.300 ;
        RECT 4.300 281.940 196.000 283.100 ;
        RECT 4.000 279.740 196.000 281.940 ;
        RECT 4.300 278.580 196.000 279.740 ;
        RECT 4.000 276.380 196.000 278.580 ;
        RECT 4.300 275.220 196.000 276.380 ;
        RECT 4.000 266.300 196.000 275.220 ;
        RECT 4.300 265.140 195.700 266.300 ;
        RECT 4.000 259.580 196.000 265.140 ;
        RECT 4.300 258.420 196.000 259.580 ;
        RECT 4.000 256.220 196.000 258.420 ;
        RECT 4.300 255.060 196.000 256.220 ;
        RECT 4.000 252.860 196.000 255.060 ;
        RECT 4.300 251.700 196.000 252.860 ;
        RECT 4.000 249.500 196.000 251.700 ;
        RECT 4.300 248.340 195.700 249.500 ;
        RECT 4.000 246.140 196.000 248.340 ;
        RECT 4.300 244.980 196.000 246.140 ;
        RECT 4.000 242.780 196.000 244.980 ;
        RECT 4.300 241.620 196.000 242.780 ;
        RECT 4.000 239.420 196.000 241.620 ;
        RECT 4.300 238.260 196.000 239.420 ;
        RECT 4.000 236.060 196.000 238.260 ;
        RECT 4.000 234.900 195.700 236.060 ;
        RECT 4.000 232.700 196.000 234.900 ;
        RECT 4.000 231.540 195.700 232.700 ;
        RECT 4.000 222.620 196.000 231.540 ;
        RECT 4.300 221.460 196.000 222.620 ;
        RECT 4.000 219.260 196.000 221.460 ;
        RECT 4.300 218.100 196.000 219.260 ;
        RECT 4.000 212.540 196.000 218.100 ;
        RECT 4.000 211.380 195.700 212.540 ;
        RECT 4.000 209.180 196.000 211.380 ;
        RECT 4.000 208.020 195.700 209.180 ;
        RECT 4.000 202.460 196.000 208.020 ;
        RECT 4.300 201.300 196.000 202.460 ;
        RECT 4.000 199.100 196.000 201.300 ;
        RECT 4.300 197.940 196.000 199.100 ;
        RECT 4.000 195.740 196.000 197.940 ;
        RECT 4.300 194.580 195.700 195.740 ;
        RECT 4.000 182.300 196.000 194.580 ;
        RECT 4.000 181.140 195.700 182.300 ;
        RECT 4.000 165.500 196.000 181.140 ;
        RECT 4.300 164.340 196.000 165.500 ;
        RECT 4.000 155.420 196.000 164.340 ;
        RECT 4.000 154.260 195.700 155.420 ;
        RECT 4.000 152.060 196.000 154.260 ;
        RECT 4.000 150.900 195.700 152.060 ;
        RECT 4.000 115.100 196.000 150.900 ;
        RECT 4.000 113.940 195.700 115.100 ;
        RECT 4.000 15.540 196.000 113.940 ;
      LAYER Metal4 ;
        RECT 93.100 169.770 98.740 311.830 ;
        RECT 100.940 169.770 174.580 311.830 ;
  END
END riscv_top
END LIBRARY

