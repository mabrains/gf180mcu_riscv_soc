magic
tech gf180mcuD
magscale 1 5
timestamp 1700067814
<< obsm1 >>
rect 672 1538 89320 98489
<< metal2 >>
rect 2352 99600 2408 100000
rect 2912 99600 2968 100000
rect 3472 99600 3528 100000
rect 4032 99600 4088 100000
rect 4592 99600 4648 100000
rect 5152 99600 5208 100000
rect 5712 99600 5768 100000
rect 6272 99600 6328 100000
rect 6832 99600 6888 100000
rect 7392 99600 7448 100000
rect 7952 99600 8008 100000
rect 8512 99600 8568 100000
rect 9072 99600 9128 100000
rect 9632 99600 9688 100000
rect 10192 99600 10248 100000
rect 10752 99600 10808 100000
rect 11312 99600 11368 100000
rect 11872 99600 11928 100000
rect 12432 99600 12488 100000
rect 12992 99600 13048 100000
rect 13552 99600 13608 100000
rect 14112 99600 14168 100000
rect 14672 99600 14728 100000
rect 15232 99600 15288 100000
rect 15792 99600 15848 100000
rect 16352 99600 16408 100000
rect 16912 99600 16968 100000
rect 17472 99600 17528 100000
rect 18032 99600 18088 100000
rect 18592 99600 18648 100000
rect 19152 99600 19208 100000
rect 19712 99600 19768 100000
rect 20272 99600 20328 100000
rect 20832 99600 20888 100000
rect 21392 99600 21448 100000
rect 21952 99600 22008 100000
rect 22512 99600 22568 100000
rect 23072 99600 23128 100000
rect 23632 99600 23688 100000
rect 24192 99600 24248 100000
rect 24752 99600 24808 100000
rect 25312 99600 25368 100000
rect 25872 99600 25928 100000
rect 26432 99600 26488 100000
rect 26992 99600 27048 100000
rect 27552 99600 27608 100000
rect 28112 99600 28168 100000
rect 28672 99600 28728 100000
rect 29232 99600 29288 100000
rect 29792 99600 29848 100000
rect 30352 99600 30408 100000
rect 30912 99600 30968 100000
rect 31472 99600 31528 100000
rect 32032 99600 32088 100000
rect 32592 99600 32648 100000
rect 33152 99600 33208 100000
rect 33712 99600 33768 100000
rect 34272 99600 34328 100000
rect 34832 99600 34888 100000
rect 35392 99600 35448 100000
rect 35952 99600 36008 100000
rect 36512 99600 36568 100000
rect 37072 99600 37128 100000
rect 37632 99600 37688 100000
rect 38192 99600 38248 100000
rect 38752 99600 38808 100000
rect 39312 99600 39368 100000
rect 39872 99600 39928 100000
rect 40432 99600 40488 100000
rect 40992 99600 41048 100000
rect 41552 99600 41608 100000
rect 42112 99600 42168 100000
rect 42672 99600 42728 100000
rect 43232 99600 43288 100000
rect 43792 99600 43848 100000
rect 44352 99600 44408 100000
rect 44912 99600 44968 100000
rect 45472 99600 45528 100000
rect 46032 99600 46088 100000
rect 46592 99600 46648 100000
rect 47152 99600 47208 100000
rect 47712 99600 47768 100000
rect 48272 99600 48328 100000
rect 48832 99600 48888 100000
rect 49392 99600 49448 100000
rect 49952 99600 50008 100000
rect 50512 99600 50568 100000
rect 51072 99600 51128 100000
rect 51632 99600 51688 100000
rect 52192 99600 52248 100000
rect 52752 99600 52808 100000
rect 53312 99600 53368 100000
rect 53872 99600 53928 100000
rect 54432 99600 54488 100000
rect 54992 99600 55048 100000
rect 55552 99600 55608 100000
rect 56112 99600 56168 100000
rect 56672 99600 56728 100000
rect 57232 99600 57288 100000
rect 57792 99600 57848 100000
rect 58352 99600 58408 100000
rect 58912 99600 58968 100000
rect 59472 99600 59528 100000
rect 60032 99600 60088 100000
rect 60592 99600 60648 100000
rect 61152 99600 61208 100000
rect 61712 99600 61768 100000
rect 62272 99600 62328 100000
rect 62832 99600 62888 100000
rect 63392 99600 63448 100000
rect 63952 99600 64008 100000
rect 64512 99600 64568 100000
rect 65072 99600 65128 100000
rect 65632 99600 65688 100000
rect 66192 99600 66248 100000
rect 66752 99600 66808 100000
rect 67312 99600 67368 100000
rect 67872 99600 67928 100000
rect 68432 99600 68488 100000
rect 68992 99600 69048 100000
rect 69552 99600 69608 100000
rect 70112 99600 70168 100000
rect 70672 99600 70728 100000
rect 71232 99600 71288 100000
rect 71792 99600 71848 100000
rect 72352 99600 72408 100000
rect 72912 99600 72968 100000
rect 73472 99600 73528 100000
rect 74032 99600 74088 100000
rect 74592 99600 74648 100000
rect 75152 99600 75208 100000
rect 75712 99600 75768 100000
rect 76272 99600 76328 100000
rect 76832 99600 76888 100000
rect 77392 99600 77448 100000
rect 77952 99600 78008 100000
rect 78512 99600 78568 100000
rect 79072 99600 79128 100000
rect 79632 99600 79688 100000
rect 80192 99600 80248 100000
rect 80752 99600 80808 100000
rect 81312 99600 81368 100000
rect 81872 99600 81928 100000
rect 82432 99600 82488 100000
rect 82992 99600 83048 100000
rect 83552 99600 83608 100000
rect 84112 99600 84168 100000
rect 84672 99600 84728 100000
rect 85232 99600 85288 100000
rect 85792 99600 85848 100000
rect 86352 99600 86408 100000
rect 86912 99600 86968 100000
rect 87472 99600 87528 100000
rect 2576 0 2632 400
rect 4928 0 4984 400
rect 7280 0 7336 400
rect 9632 0 9688 400
rect 11984 0 12040 400
rect 14336 0 14392 400
rect 16688 0 16744 400
rect 19040 0 19096 400
rect 21392 0 21448 400
rect 23744 0 23800 400
rect 26096 0 26152 400
rect 28448 0 28504 400
rect 30800 0 30856 400
rect 33152 0 33208 400
rect 35504 0 35560 400
rect 37856 0 37912 400
rect 40208 0 40264 400
rect 42560 0 42616 400
rect 44912 0 44968 400
rect 47264 0 47320 400
rect 49616 0 49672 400
rect 51968 0 52024 400
rect 54320 0 54376 400
rect 56672 0 56728 400
rect 59024 0 59080 400
rect 61376 0 61432 400
rect 63728 0 63784 400
rect 66080 0 66136 400
rect 68432 0 68488 400
rect 70784 0 70840 400
rect 73136 0 73192 400
rect 75488 0 75544 400
rect 77840 0 77896 400
rect 80192 0 80248 400
rect 82544 0 82600 400
rect 84896 0 84952 400
rect 87248 0 87304 400
<< obsm2 >>
rect 798 99570 2322 99666
rect 2438 99570 2882 99666
rect 2998 99570 3442 99666
rect 3558 99570 4002 99666
rect 4118 99570 4562 99666
rect 4678 99570 5122 99666
rect 5238 99570 5682 99666
rect 5798 99570 6242 99666
rect 6358 99570 6802 99666
rect 6918 99570 7362 99666
rect 7478 99570 7922 99666
rect 8038 99570 8482 99666
rect 8598 99570 9042 99666
rect 9158 99570 9602 99666
rect 9718 99570 10162 99666
rect 10278 99570 10722 99666
rect 10838 99570 11282 99666
rect 11398 99570 11842 99666
rect 11958 99570 12402 99666
rect 12518 99570 12962 99666
rect 13078 99570 13522 99666
rect 13638 99570 14082 99666
rect 14198 99570 14642 99666
rect 14758 99570 15202 99666
rect 15318 99570 15762 99666
rect 15878 99570 16322 99666
rect 16438 99570 16882 99666
rect 16998 99570 17442 99666
rect 17558 99570 18002 99666
rect 18118 99570 18562 99666
rect 18678 99570 19122 99666
rect 19238 99570 19682 99666
rect 19798 99570 20242 99666
rect 20358 99570 20802 99666
rect 20918 99570 21362 99666
rect 21478 99570 21922 99666
rect 22038 99570 22482 99666
rect 22598 99570 23042 99666
rect 23158 99570 23602 99666
rect 23718 99570 24162 99666
rect 24278 99570 24722 99666
rect 24838 99570 25282 99666
rect 25398 99570 25842 99666
rect 25958 99570 26402 99666
rect 26518 99570 26962 99666
rect 27078 99570 27522 99666
rect 27638 99570 28082 99666
rect 28198 99570 28642 99666
rect 28758 99570 29202 99666
rect 29318 99570 29762 99666
rect 29878 99570 30322 99666
rect 30438 99570 30882 99666
rect 30998 99570 31442 99666
rect 31558 99570 32002 99666
rect 32118 99570 32562 99666
rect 32678 99570 33122 99666
rect 33238 99570 33682 99666
rect 33798 99570 34242 99666
rect 34358 99570 34802 99666
rect 34918 99570 35362 99666
rect 35478 99570 35922 99666
rect 36038 99570 36482 99666
rect 36598 99570 37042 99666
rect 37158 99570 37602 99666
rect 37718 99570 38162 99666
rect 38278 99570 38722 99666
rect 38838 99570 39282 99666
rect 39398 99570 39842 99666
rect 39958 99570 40402 99666
rect 40518 99570 40962 99666
rect 41078 99570 41522 99666
rect 41638 99570 42082 99666
rect 42198 99570 42642 99666
rect 42758 99570 43202 99666
rect 43318 99570 43762 99666
rect 43878 99570 44322 99666
rect 44438 99570 44882 99666
rect 44998 99570 45442 99666
rect 45558 99570 46002 99666
rect 46118 99570 46562 99666
rect 46678 99570 47122 99666
rect 47238 99570 47682 99666
rect 47798 99570 48242 99666
rect 48358 99570 48802 99666
rect 48918 99570 49362 99666
rect 49478 99570 49922 99666
rect 50038 99570 50482 99666
rect 50598 99570 51042 99666
rect 51158 99570 51602 99666
rect 51718 99570 52162 99666
rect 52278 99570 52722 99666
rect 52838 99570 53282 99666
rect 53398 99570 53842 99666
rect 53958 99570 54402 99666
rect 54518 99570 54962 99666
rect 55078 99570 55522 99666
rect 55638 99570 56082 99666
rect 56198 99570 56642 99666
rect 56758 99570 57202 99666
rect 57318 99570 57762 99666
rect 57878 99570 58322 99666
rect 58438 99570 58882 99666
rect 58998 99570 59442 99666
rect 59558 99570 60002 99666
rect 60118 99570 60562 99666
rect 60678 99570 61122 99666
rect 61238 99570 61682 99666
rect 61798 99570 62242 99666
rect 62358 99570 62802 99666
rect 62918 99570 63362 99666
rect 63478 99570 63922 99666
rect 64038 99570 64482 99666
rect 64598 99570 65042 99666
rect 65158 99570 65602 99666
rect 65718 99570 66162 99666
rect 66278 99570 66722 99666
rect 66838 99570 67282 99666
rect 67398 99570 67842 99666
rect 67958 99570 68402 99666
rect 68518 99570 68962 99666
rect 69078 99570 69522 99666
rect 69638 99570 70082 99666
rect 70198 99570 70642 99666
rect 70758 99570 71202 99666
rect 71318 99570 71762 99666
rect 71878 99570 72322 99666
rect 72438 99570 72882 99666
rect 72998 99570 73442 99666
rect 73558 99570 74002 99666
rect 74118 99570 74562 99666
rect 74678 99570 75122 99666
rect 75238 99570 75682 99666
rect 75798 99570 76242 99666
rect 76358 99570 76802 99666
rect 76918 99570 77362 99666
rect 77478 99570 77922 99666
rect 78038 99570 78482 99666
rect 78598 99570 79042 99666
rect 79158 99570 79602 99666
rect 79718 99570 80162 99666
rect 80278 99570 80722 99666
rect 80838 99570 81282 99666
rect 81398 99570 81842 99666
rect 81958 99570 82402 99666
rect 82518 99570 82962 99666
rect 83078 99570 83522 99666
rect 83638 99570 84082 99666
rect 84198 99570 84642 99666
rect 84758 99570 85202 99666
rect 85318 99570 85762 99666
rect 85878 99570 86322 99666
rect 86438 99570 86882 99666
rect 86998 99570 87442 99666
rect 87558 99570 89194 99666
rect 798 430 89194 99570
rect 798 350 2546 430
rect 2662 350 4898 430
rect 5014 350 7250 430
rect 7366 350 9602 430
rect 9718 350 11954 430
rect 12070 350 14306 430
rect 14422 350 16658 430
rect 16774 350 19010 430
rect 19126 350 21362 430
rect 21478 350 23714 430
rect 23830 350 26066 430
rect 26182 350 28418 430
rect 28534 350 30770 430
rect 30886 350 33122 430
rect 33238 350 35474 430
rect 35590 350 37826 430
rect 37942 350 40178 430
rect 40294 350 42530 430
rect 42646 350 44882 430
rect 44998 350 47234 430
rect 47350 350 49586 430
rect 49702 350 51938 430
rect 52054 350 54290 430
rect 54406 350 56642 430
rect 56758 350 58994 430
rect 59110 350 61346 430
rect 61462 350 63698 430
rect 63814 350 66050 430
rect 66166 350 68402 430
rect 68518 350 70754 430
rect 70870 350 73106 430
rect 73222 350 75458 430
rect 75574 350 77810 430
rect 77926 350 80162 430
rect 80278 350 82514 430
rect 82630 350 84866 430
rect 84982 350 87218 430
rect 87334 350 89194 430
<< metal3 >>
rect 0 97552 400 97608
rect 89600 96768 90000 96824
rect 0 96432 400 96488
rect 0 95312 400 95368
rect 89600 94640 90000 94696
rect 0 94192 400 94248
rect 0 93072 400 93128
rect 89600 92512 90000 92568
rect 0 91952 400 92008
rect 0 90832 400 90888
rect 89600 90384 90000 90440
rect 0 89712 400 89768
rect 0 88592 400 88648
rect 89600 88256 90000 88312
rect 0 87472 400 87528
rect 0 86352 400 86408
rect 89600 86128 90000 86184
rect 0 85232 400 85288
rect 0 84112 400 84168
rect 89600 84000 90000 84056
rect 0 82992 400 83048
rect 0 81872 400 81928
rect 89600 81872 90000 81928
rect 0 80752 400 80808
rect 89600 79744 90000 79800
rect 0 79632 400 79688
rect 0 78512 400 78568
rect 89600 77616 90000 77672
rect 0 77392 400 77448
rect 0 76272 400 76328
rect 89600 75488 90000 75544
rect 0 75152 400 75208
rect 0 74032 400 74088
rect 89600 73360 90000 73416
rect 0 72912 400 72968
rect 0 71792 400 71848
rect 89600 71232 90000 71288
rect 0 70672 400 70728
rect 0 69552 400 69608
rect 89600 69104 90000 69160
rect 0 68432 400 68488
rect 0 67312 400 67368
rect 89600 66976 90000 67032
rect 0 66192 400 66248
rect 0 65072 400 65128
rect 89600 64848 90000 64904
rect 0 63952 400 64008
rect 0 62832 400 62888
rect 89600 62720 90000 62776
rect 0 61712 400 61768
rect 0 60592 400 60648
rect 89600 60592 90000 60648
rect 0 59472 400 59528
rect 89600 58464 90000 58520
rect 0 58352 400 58408
rect 0 57232 400 57288
rect 89600 56336 90000 56392
rect 0 56112 400 56168
rect 0 54992 400 55048
rect 89600 54208 90000 54264
rect 0 53872 400 53928
rect 0 52752 400 52808
rect 89600 52080 90000 52136
rect 0 51632 400 51688
rect 0 50512 400 50568
rect 89600 49952 90000 50008
rect 0 49392 400 49448
rect 0 48272 400 48328
rect 89600 47824 90000 47880
rect 0 47152 400 47208
rect 0 46032 400 46088
rect 89600 45696 90000 45752
rect 0 44912 400 44968
rect 0 43792 400 43848
rect 89600 43568 90000 43624
rect 0 42672 400 42728
rect 0 41552 400 41608
rect 89600 41440 90000 41496
rect 0 40432 400 40488
rect 0 39312 400 39368
rect 89600 39312 90000 39368
rect 0 38192 400 38248
rect 89600 37184 90000 37240
rect 0 37072 400 37128
rect 0 35952 400 36008
rect 89600 35056 90000 35112
rect 0 34832 400 34888
rect 0 33712 400 33768
rect 89600 32928 90000 32984
rect 0 32592 400 32648
rect 0 31472 400 31528
rect 89600 30800 90000 30856
rect 0 30352 400 30408
rect 0 29232 400 29288
rect 89600 28672 90000 28728
rect 0 28112 400 28168
rect 0 26992 400 27048
rect 89600 26544 90000 26600
rect 0 25872 400 25928
rect 0 24752 400 24808
rect 89600 24416 90000 24472
rect 0 23632 400 23688
rect 0 22512 400 22568
rect 89600 22288 90000 22344
rect 0 21392 400 21448
rect 0 20272 400 20328
rect 89600 20160 90000 20216
rect 0 19152 400 19208
rect 0 18032 400 18088
rect 89600 18032 90000 18088
rect 0 16912 400 16968
rect 89600 15904 90000 15960
rect 0 15792 400 15848
rect 0 14672 400 14728
rect 89600 13776 90000 13832
rect 0 13552 400 13608
rect 0 12432 400 12488
rect 89600 11648 90000 11704
rect 0 11312 400 11368
rect 0 10192 400 10248
rect 89600 9520 90000 9576
rect 0 9072 400 9128
rect 0 7952 400 8008
rect 89600 7392 90000 7448
rect 0 6832 400 6888
rect 0 5712 400 5768
rect 89600 5264 90000 5320
rect 0 4592 400 4648
rect 0 3472 400 3528
rect 89600 3136 90000 3192
rect 0 2352 400 2408
<< obsm3 >>
rect 350 97638 89600 98406
rect 430 97522 89600 97638
rect 350 96854 89600 97522
rect 350 96738 89570 96854
rect 350 96518 89600 96738
rect 430 96402 89600 96518
rect 350 95398 89600 96402
rect 430 95282 89600 95398
rect 350 94726 89600 95282
rect 350 94610 89570 94726
rect 350 94278 89600 94610
rect 430 94162 89600 94278
rect 350 93158 89600 94162
rect 430 93042 89600 93158
rect 350 92598 89600 93042
rect 350 92482 89570 92598
rect 350 92038 89600 92482
rect 430 91922 89600 92038
rect 350 90918 89600 91922
rect 430 90802 89600 90918
rect 350 90470 89600 90802
rect 350 90354 89570 90470
rect 350 89798 89600 90354
rect 430 89682 89600 89798
rect 350 88678 89600 89682
rect 430 88562 89600 88678
rect 350 88342 89600 88562
rect 350 88226 89570 88342
rect 350 87558 89600 88226
rect 430 87442 89600 87558
rect 350 86438 89600 87442
rect 430 86322 89600 86438
rect 350 86214 89600 86322
rect 350 86098 89570 86214
rect 350 85318 89600 86098
rect 430 85202 89600 85318
rect 350 84198 89600 85202
rect 430 84086 89600 84198
rect 430 84082 89570 84086
rect 350 83970 89570 84082
rect 350 83078 89600 83970
rect 430 82962 89600 83078
rect 350 81958 89600 82962
rect 430 81842 89570 81958
rect 350 80838 89600 81842
rect 430 80722 89600 80838
rect 350 79830 89600 80722
rect 350 79718 89570 79830
rect 430 79714 89570 79718
rect 430 79602 89600 79714
rect 350 78598 89600 79602
rect 430 78482 89600 78598
rect 350 77702 89600 78482
rect 350 77586 89570 77702
rect 350 77478 89600 77586
rect 430 77362 89600 77478
rect 350 76358 89600 77362
rect 430 76242 89600 76358
rect 350 75574 89600 76242
rect 350 75458 89570 75574
rect 350 75238 89600 75458
rect 430 75122 89600 75238
rect 350 74118 89600 75122
rect 430 74002 89600 74118
rect 350 73446 89600 74002
rect 350 73330 89570 73446
rect 350 72998 89600 73330
rect 430 72882 89600 72998
rect 350 71878 89600 72882
rect 430 71762 89600 71878
rect 350 71318 89600 71762
rect 350 71202 89570 71318
rect 350 70758 89600 71202
rect 430 70642 89600 70758
rect 350 69638 89600 70642
rect 430 69522 89600 69638
rect 350 69190 89600 69522
rect 350 69074 89570 69190
rect 350 68518 89600 69074
rect 430 68402 89600 68518
rect 350 67398 89600 68402
rect 430 67282 89600 67398
rect 350 67062 89600 67282
rect 350 66946 89570 67062
rect 350 66278 89600 66946
rect 430 66162 89600 66278
rect 350 65158 89600 66162
rect 430 65042 89600 65158
rect 350 64934 89600 65042
rect 350 64818 89570 64934
rect 350 64038 89600 64818
rect 430 63922 89600 64038
rect 350 62918 89600 63922
rect 430 62806 89600 62918
rect 430 62802 89570 62806
rect 350 62690 89570 62802
rect 350 61798 89600 62690
rect 430 61682 89600 61798
rect 350 60678 89600 61682
rect 430 60562 89570 60678
rect 350 59558 89600 60562
rect 430 59442 89600 59558
rect 350 58550 89600 59442
rect 350 58438 89570 58550
rect 430 58434 89570 58438
rect 430 58322 89600 58434
rect 350 57318 89600 58322
rect 430 57202 89600 57318
rect 350 56422 89600 57202
rect 350 56306 89570 56422
rect 350 56198 89600 56306
rect 430 56082 89600 56198
rect 350 55078 89600 56082
rect 430 54962 89600 55078
rect 350 54294 89600 54962
rect 350 54178 89570 54294
rect 350 53958 89600 54178
rect 430 53842 89600 53958
rect 350 52838 89600 53842
rect 430 52722 89600 52838
rect 350 52166 89600 52722
rect 350 52050 89570 52166
rect 350 51718 89600 52050
rect 430 51602 89600 51718
rect 350 50598 89600 51602
rect 430 50482 89600 50598
rect 350 50038 89600 50482
rect 350 49922 89570 50038
rect 350 49478 89600 49922
rect 430 49362 89600 49478
rect 350 48358 89600 49362
rect 430 48242 89600 48358
rect 350 47910 89600 48242
rect 350 47794 89570 47910
rect 350 47238 89600 47794
rect 430 47122 89600 47238
rect 350 46118 89600 47122
rect 430 46002 89600 46118
rect 350 45782 89600 46002
rect 350 45666 89570 45782
rect 350 44998 89600 45666
rect 430 44882 89600 44998
rect 350 43878 89600 44882
rect 430 43762 89600 43878
rect 350 43654 89600 43762
rect 350 43538 89570 43654
rect 350 42758 89600 43538
rect 430 42642 89600 42758
rect 350 41638 89600 42642
rect 430 41526 89600 41638
rect 430 41522 89570 41526
rect 350 41410 89570 41522
rect 350 40518 89600 41410
rect 430 40402 89600 40518
rect 350 39398 89600 40402
rect 430 39282 89570 39398
rect 350 38278 89600 39282
rect 430 38162 89600 38278
rect 350 37270 89600 38162
rect 350 37158 89570 37270
rect 430 37154 89570 37158
rect 430 37042 89600 37154
rect 350 36038 89600 37042
rect 430 35922 89600 36038
rect 350 35142 89600 35922
rect 350 35026 89570 35142
rect 350 34918 89600 35026
rect 430 34802 89600 34918
rect 350 33798 89600 34802
rect 430 33682 89600 33798
rect 350 33014 89600 33682
rect 350 32898 89570 33014
rect 350 32678 89600 32898
rect 430 32562 89600 32678
rect 350 31558 89600 32562
rect 430 31442 89600 31558
rect 350 30886 89600 31442
rect 350 30770 89570 30886
rect 350 30438 89600 30770
rect 430 30322 89600 30438
rect 350 29318 89600 30322
rect 430 29202 89600 29318
rect 350 28758 89600 29202
rect 350 28642 89570 28758
rect 350 28198 89600 28642
rect 430 28082 89600 28198
rect 350 27078 89600 28082
rect 430 26962 89600 27078
rect 350 26630 89600 26962
rect 350 26514 89570 26630
rect 350 25958 89600 26514
rect 430 25842 89600 25958
rect 350 24838 89600 25842
rect 430 24722 89600 24838
rect 350 24502 89600 24722
rect 350 24386 89570 24502
rect 350 23718 89600 24386
rect 430 23602 89600 23718
rect 350 22598 89600 23602
rect 430 22482 89600 22598
rect 350 22374 89600 22482
rect 350 22258 89570 22374
rect 350 21478 89600 22258
rect 430 21362 89600 21478
rect 350 20358 89600 21362
rect 430 20246 89600 20358
rect 430 20242 89570 20246
rect 350 20130 89570 20242
rect 350 19238 89600 20130
rect 430 19122 89600 19238
rect 350 18118 89600 19122
rect 430 18002 89570 18118
rect 350 16998 89600 18002
rect 430 16882 89600 16998
rect 350 15990 89600 16882
rect 350 15878 89570 15990
rect 430 15874 89570 15878
rect 430 15762 89600 15874
rect 350 14758 89600 15762
rect 430 14642 89600 14758
rect 350 13862 89600 14642
rect 350 13746 89570 13862
rect 350 13638 89600 13746
rect 430 13522 89600 13638
rect 350 12518 89600 13522
rect 430 12402 89600 12518
rect 350 11734 89600 12402
rect 350 11618 89570 11734
rect 350 11398 89600 11618
rect 430 11282 89600 11398
rect 350 10278 89600 11282
rect 430 10162 89600 10278
rect 350 9606 89600 10162
rect 350 9490 89570 9606
rect 350 9158 89600 9490
rect 430 9042 89600 9158
rect 350 8038 89600 9042
rect 430 7922 89600 8038
rect 350 7478 89600 7922
rect 350 7362 89570 7478
rect 350 6918 89600 7362
rect 430 6802 89600 6918
rect 350 5798 89600 6802
rect 430 5682 89600 5798
rect 350 5350 89600 5682
rect 350 5234 89570 5350
rect 350 4678 89600 5234
rect 430 4562 89600 4678
rect 350 3558 89600 4562
rect 430 3442 89600 3558
rect 350 3222 89600 3442
rect 350 3106 89570 3222
rect 350 2438 89600 3106
rect 430 2322 89600 2438
rect 350 1554 89600 2322
<< metal4 >>
rect 2224 1538 2384 98422
rect 9904 1538 10064 98422
rect 17584 1538 17744 98422
rect 25264 1538 25424 98422
rect 32944 1538 33104 98422
rect 40624 1538 40784 98422
rect 48304 1538 48464 98422
rect 55984 1538 56144 98422
rect 63664 1538 63824 98422
rect 71344 1538 71504 98422
rect 79024 1538 79184 98422
rect 86704 1538 86864 98422
<< obsm4 >>
rect 1694 2473 2194 98215
rect 2414 2473 9874 98215
rect 10094 2473 17554 98215
rect 17774 2473 25234 98215
rect 25454 2473 32914 98215
rect 33134 2473 40594 98215
rect 40814 2473 48274 98215
rect 48494 2473 55954 98215
rect 56174 2473 63634 98215
rect 63854 2473 71314 98215
rect 71534 2473 78994 98215
rect 79214 2473 86674 98215
rect 86894 2473 88802 98215
<< obsm5 >>
rect 2470 21623 81250 98167
<< labels >>
rlabel metal4 s 2224 1538 2384 98422 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 98422 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 98422 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 98422 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 98422 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 98422 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 98422 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 98422 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 98422 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 98422 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 98422 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 98422 6 VSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 4592 400 4648 6 cfg_strap_pad_ctrl
port 3 nsew signal input
rlabel metal3 s 89600 3136 90000 3192 6 digital_io_in[0]
port 4 nsew signal input
rlabel metal3 s 89600 66976 90000 67032 6 digital_io_in[10]
port 5 nsew signal input
rlabel metal3 s 89600 73360 90000 73416 6 digital_io_in[11]
port 6 nsew signal input
rlabel metal3 s 89600 79744 90000 79800 6 digital_io_in[12]
port 7 nsew signal input
rlabel metal3 s 89600 86128 90000 86184 6 digital_io_in[13]
port 8 nsew signal input
rlabel metal3 s 89600 92512 90000 92568 6 digital_io_in[14]
port 9 nsew signal input
rlabel metal2 s 86352 99600 86408 100000 6 digital_io_in[15]
port 10 nsew signal input
rlabel metal2 s 84672 99600 84728 100000 6 digital_io_in[16]
port 11 nsew signal input
rlabel metal2 s 82992 99600 83048 100000 6 digital_io_in[17]
port 12 nsew signal input
rlabel metal2 s 81312 99600 81368 100000 6 digital_io_in[18]
port 13 nsew signal input
rlabel metal2 s 79632 99600 79688 100000 6 digital_io_in[19]
port 14 nsew signal input
rlabel metal3 s 89600 9520 90000 9576 6 digital_io_in[1]
port 15 nsew signal input
rlabel metal2 s 77952 99600 78008 100000 6 digital_io_in[20]
port 16 nsew signal input
rlabel metal2 s 76272 99600 76328 100000 6 digital_io_in[21]
port 17 nsew signal input
rlabel metal2 s 74592 99600 74648 100000 6 digital_io_in[22]
port 18 nsew signal input
rlabel metal2 s 72912 99600 72968 100000 6 digital_io_in[23]
port 19 nsew signal input
rlabel metal2 s 25312 99600 25368 100000 6 digital_io_in[24]
port 20 nsew signal input
rlabel metal2 s 23632 99600 23688 100000 6 digital_io_in[25]
port 21 nsew signal input
rlabel metal2 s 21952 99600 22008 100000 6 digital_io_in[26]
port 22 nsew signal input
rlabel metal2 s 20272 99600 20328 100000 6 digital_io_in[27]
port 23 nsew signal input
rlabel metal2 s 18592 99600 18648 100000 6 digital_io_in[28]
port 24 nsew signal input
rlabel metal2 s 16912 99600 16968 100000 6 digital_io_in[29]
port 25 nsew signal input
rlabel metal3 s 89600 15904 90000 15960 6 digital_io_in[2]
port 26 nsew signal input
rlabel metal2 s 15232 99600 15288 100000 6 digital_io_in[30]
port 27 nsew signal input
rlabel metal2 s 13552 99600 13608 100000 6 digital_io_in[31]
port 28 nsew signal input
rlabel metal2 s 11872 99600 11928 100000 6 digital_io_in[32]
port 29 nsew signal input
rlabel metal2 s 10192 99600 10248 100000 6 digital_io_in[33]
port 30 nsew signal input
rlabel metal2 s 8512 99600 8568 100000 6 digital_io_in[34]
port 31 nsew signal input
rlabel metal2 s 6832 99600 6888 100000 6 digital_io_in[35]
port 32 nsew signal input
rlabel metal2 s 5152 99600 5208 100000 6 digital_io_in[36]
port 33 nsew signal input
rlabel metal2 s 3472 99600 3528 100000 6 digital_io_in[37]
port 34 nsew signal input
rlabel metal3 s 89600 22288 90000 22344 6 digital_io_in[3]
port 35 nsew signal input
rlabel metal3 s 89600 28672 90000 28728 6 digital_io_in[4]
port 36 nsew signal input
rlabel metal3 s 89600 35056 90000 35112 6 digital_io_in[5]
port 37 nsew signal input
rlabel metal3 s 89600 41440 90000 41496 6 digital_io_in[6]
port 38 nsew signal input
rlabel metal3 s 89600 47824 90000 47880 6 digital_io_in[7]
port 39 nsew signal input
rlabel metal3 s 89600 54208 90000 54264 6 digital_io_in[8]
port 40 nsew signal input
rlabel metal3 s 89600 60592 90000 60648 6 digital_io_in[9]
port 41 nsew signal input
rlabel metal3 s 89600 7392 90000 7448 6 digital_io_oen[0]
port 42 nsew signal output
rlabel metal3 s 89600 71232 90000 71288 6 digital_io_oen[10]
port 43 nsew signal output
rlabel metal3 s 89600 77616 90000 77672 6 digital_io_oen[11]
port 44 nsew signal output
rlabel metal3 s 89600 84000 90000 84056 6 digital_io_oen[12]
port 45 nsew signal output
rlabel metal3 s 89600 90384 90000 90440 6 digital_io_oen[13]
port 46 nsew signal output
rlabel metal3 s 89600 96768 90000 96824 6 digital_io_oen[14]
port 47 nsew signal output
rlabel metal2 s 87472 99600 87528 100000 6 digital_io_oen[15]
port 48 nsew signal output
rlabel metal2 s 85792 99600 85848 100000 6 digital_io_oen[16]
port 49 nsew signal output
rlabel metal2 s 84112 99600 84168 100000 6 digital_io_oen[17]
port 50 nsew signal output
rlabel metal2 s 82432 99600 82488 100000 6 digital_io_oen[18]
port 51 nsew signal output
rlabel metal2 s 80752 99600 80808 100000 6 digital_io_oen[19]
port 52 nsew signal output
rlabel metal3 s 89600 13776 90000 13832 6 digital_io_oen[1]
port 53 nsew signal output
rlabel metal2 s 79072 99600 79128 100000 6 digital_io_oen[20]
port 54 nsew signal output
rlabel metal2 s 77392 99600 77448 100000 6 digital_io_oen[21]
port 55 nsew signal output
rlabel metal2 s 75712 99600 75768 100000 6 digital_io_oen[22]
port 56 nsew signal output
rlabel metal2 s 74032 99600 74088 100000 6 digital_io_oen[23]
port 57 nsew signal output
rlabel metal2 s 24192 99600 24248 100000 6 digital_io_oen[24]
port 58 nsew signal output
rlabel metal2 s 22512 99600 22568 100000 6 digital_io_oen[25]
port 59 nsew signal output
rlabel metal2 s 20832 99600 20888 100000 6 digital_io_oen[26]
port 60 nsew signal output
rlabel metal2 s 19152 99600 19208 100000 6 digital_io_oen[27]
port 61 nsew signal output
rlabel metal2 s 17472 99600 17528 100000 6 digital_io_oen[28]
port 62 nsew signal output
rlabel metal2 s 15792 99600 15848 100000 6 digital_io_oen[29]
port 63 nsew signal output
rlabel metal3 s 89600 20160 90000 20216 6 digital_io_oen[2]
port 64 nsew signal output
rlabel metal2 s 14112 99600 14168 100000 6 digital_io_oen[30]
port 65 nsew signal output
rlabel metal2 s 12432 99600 12488 100000 6 digital_io_oen[31]
port 66 nsew signal output
rlabel metal2 s 10752 99600 10808 100000 6 digital_io_oen[32]
port 67 nsew signal output
rlabel metal2 s 9072 99600 9128 100000 6 digital_io_oen[33]
port 68 nsew signal output
rlabel metal2 s 7392 99600 7448 100000 6 digital_io_oen[34]
port 69 nsew signal output
rlabel metal2 s 5712 99600 5768 100000 6 digital_io_oen[35]
port 70 nsew signal output
rlabel metal2 s 4032 99600 4088 100000 6 digital_io_oen[36]
port 71 nsew signal output
rlabel metal2 s 2352 99600 2408 100000 6 digital_io_oen[37]
port 72 nsew signal output
rlabel metal3 s 89600 26544 90000 26600 6 digital_io_oen[3]
port 73 nsew signal output
rlabel metal3 s 89600 32928 90000 32984 6 digital_io_oen[4]
port 74 nsew signal output
rlabel metal3 s 89600 39312 90000 39368 6 digital_io_oen[5]
port 75 nsew signal output
rlabel metal3 s 89600 45696 90000 45752 6 digital_io_oen[6]
port 76 nsew signal output
rlabel metal3 s 89600 52080 90000 52136 6 digital_io_oen[7]
port 77 nsew signal output
rlabel metal3 s 89600 58464 90000 58520 6 digital_io_oen[8]
port 78 nsew signal output
rlabel metal3 s 89600 64848 90000 64904 6 digital_io_oen[9]
port 79 nsew signal output
rlabel metal3 s 89600 5264 90000 5320 6 digital_io_out[0]
port 80 nsew signal output
rlabel metal3 s 89600 69104 90000 69160 6 digital_io_out[10]
port 81 nsew signal output
rlabel metal3 s 89600 75488 90000 75544 6 digital_io_out[11]
port 82 nsew signal output
rlabel metal3 s 89600 81872 90000 81928 6 digital_io_out[12]
port 83 nsew signal output
rlabel metal3 s 89600 88256 90000 88312 6 digital_io_out[13]
port 84 nsew signal output
rlabel metal3 s 89600 94640 90000 94696 6 digital_io_out[14]
port 85 nsew signal output
rlabel metal2 s 86912 99600 86968 100000 6 digital_io_out[15]
port 86 nsew signal output
rlabel metal2 s 85232 99600 85288 100000 6 digital_io_out[16]
port 87 nsew signal output
rlabel metal2 s 83552 99600 83608 100000 6 digital_io_out[17]
port 88 nsew signal output
rlabel metal2 s 81872 99600 81928 100000 6 digital_io_out[18]
port 89 nsew signal output
rlabel metal2 s 80192 99600 80248 100000 6 digital_io_out[19]
port 90 nsew signal output
rlabel metal3 s 89600 11648 90000 11704 6 digital_io_out[1]
port 91 nsew signal output
rlabel metal2 s 78512 99600 78568 100000 6 digital_io_out[20]
port 92 nsew signal output
rlabel metal2 s 76832 99600 76888 100000 6 digital_io_out[21]
port 93 nsew signal output
rlabel metal2 s 75152 99600 75208 100000 6 digital_io_out[22]
port 94 nsew signal output
rlabel metal2 s 73472 99600 73528 100000 6 digital_io_out[23]
port 95 nsew signal output
rlabel metal2 s 24752 99600 24808 100000 6 digital_io_out[24]
port 96 nsew signal output
rlabel metal2 s 23072 99600 23128 100000 6 digital_io_out[25]
port 97 nsew signal output
rlabel metal2 s 21392 99600 21448 100000 6 digital_io_out[26]
port 98 nsew signal output
rlabel metal2 s 19712 99600 19768 100000 6 digital_io_out[27]
port 99 nsew signal output
rlabel metal2 s 18032 99600 18088 100000 6 digital_io_out[28]
port 100 nsew signal output
rlabel metal2 s 16352 99600 16408 100000 6 digital_io_out[29]
port 101 nsew signal output
rlabel metal3 s 89600 18032 90000 18088 6 digital_io_out[2]
port 102 nsew signal output
rlabel metal2 s 14672 99600 14728 100000 6 digital_io_out[30]
port 103 nsew signal output
rlabel metal2 s 12992 99600 13048 100000 6 digital_io_out[31]
port 104 nsew signal output
rlabel metal2 s 11312 99600 11368 100000 6 digital_io_out[32]
port 105 nsew signal output
rlabel metal2 s 9632 99600 9688 100000 6 digital_io_out[33]
port 106 nsew signal output
rlabel metal2 s 7952 99600 8008 100000 6 digital_io_out[34]
port 107 nsew signal output
rlabel metal2 s 6272 99600 6328 100000 6 digital_io_out[35]
port 108 nsew signal output
rlabel metal2 s 4592 99600 4648 100000 6 digital_io_out[36]
port 109 nsew signal output
rlabel metal2 s 2912 99600 2968 100000 6 digital_io_out[37]
port 110 nsew signal output
rlabel metal3 s 89600 24416 90000 24472 6 digital_io_out[3]
port 111 nsew signal output
rlabel metal3 s 89600 30800 90000 30856 6 digital_io_out[4]
port 112 nsew signal output
rlabel metal3 s 89600 37184 90000 37240 6 digital_io_out[5]
port 113 nsew signal output
rlabel metal3 s 89600 43568 90000 43624 6 digital_io_out[6]
port 114 nsew signal output
rlabel metal3 s 89600 49952 90000 50008 6 digital_io_out[7]
port 115 nsew signal output
rlabel metal3 s 89600 56336 90000 56392 6 digital_io_out[8]
port 116 nsew signal output
rlabel metal3 s 89600 62720 90000 62776 6 digital_io_out[9]
port 117 nsew signal output
rlabel metal3 s 0 3472 400 3528 6 e_reset_n
port 118 nsew signal input
rlabel metal2 s 44912 0 44968 400 6 i2cm_clk_i
port 119 nsew signal output
rlabel metal2 s 42560 0 42616 400 6 i2cm_clk_o
port 120 nsew signal input
rlabel metal2 s 47264 0 47320 400 6 i2cm_clk_oen
port 121 nsew signal input
rlabel metal2 s 54320 0 54376 400 6 i2cm_data_i
port 122 nsew signal output
rlabel metal2 s 51968 0 52024 400 6 i2cm_data_o
port 123 nsew signal input
rlabel metal2 s 49616 0 49672 400 6 i2cm_data_oen
port 124 nsew signal input
rlabel metal2 s 75488 0 75544 400 6 i2cm_intr
port 125 nsew signal input
rlabel metal2 s 9632 0 9688 400 6 i2cm_rst_n
port 126 nsew signal output
rlabel metal3 s 0 5712 400 5768 6 mclk
port 127 nsew signal input
rlabel metal3 s 0 2352 400 2408 6 p_reset_n
port 128 nsew signal input
rlabel metal2 s 73136 0 73192 400 6 pulse1m_mclk
port 129 nsew signal output
rlabel metal3 s 0 97552 400 97608 6 reg_ack
port 130 nsew signal output
rlabel metal3 s 0 20272 400 20328 6 reg_addr[0]
port 131 nsew signal input
rlabel metal3 s 0 9072 400 9128 6 reg_addr[10]
port 132 nsew signal input
rlabel metal3 s 0 19152 400 19208 6 reg_addr[1]
port 133 nsew signal input
rlabel metal3 s 0 18032 400 18088 6 reg_addr[2]
port 134 nsew signal input
rlabel metal3 s 0 16912 400 16968 6 reg_addr[3]
port 135 nsew signal input
rlabel metal3 s 0 15792 400 15848 6 reg_addr[4]
port 136 nsew signal input
rlabel metal3 s 0 14672 400 14728 6 reg_addr[5]
port 137 nsew signal input
rlabel metal3 s 0 13552 400 13608 6 reg_addr[6]
port 138 nsew signal input
rlabel metal3 s 0 12432 400 12488 6 reg_addr[7]
port 139 nsew signal input
rlabel metal3 s 0 11312 400 11368 6 reg_addr[8]
port 140 nsew signal input
rlabel metal3 s 0 10192 400 10248 6 reg_addr[9]
port 141 nsew signal input
rlabel metal3 s 0 24752 400 24808 6 reg_be[0]
port 142 nsew signal input
rlabel metal3 s 0 23632 400 23688 6 reg_be[1]
port 143 nsew signal input
rlabel metal3 s 0 22512 400 22568 6 reg_be[2]
port 144 nsew signal input
rlabel metal3 s 0 21392 400 21448 6 reg_be[3]
port 145 nsew signal input
rlabel metal3 s 0 6832 400 6888 6 reg_cs
port 146 nsew signal input
rlabel metal2 s 72352 99600 72408 100000 6 reg_peri_ack
port 147 nsew signal input
rlabel metal2 s 33712 99600 33768 100000 6 reg_peri_addr[0]
port 148 nsew signal output
rlabel metal2 s 28112 99600 28168 100000 6 reg_peri_addr[10]
port 149 nsew signal output
rlabel metal2 s 33152 99600 33208 100000 6 reg_peri_addr[1]
port 150 nsew signal output
rlabel metal2 s 32592 99600 32648 100000 6 reg_peri_addr[2]
port 151 nsew signal output
rlabel metal2 s 32032 99600 32088 100000 6 reg_peri_addr[3]
port 152 nsew signal output
rlabel metal2 s 31472 99600 31528 100000 6 reg_peri_addr[4]
port 153 nsew signal output
rlabel metal2 s 30912 99600 30968 100000 6 reg_peri_addr[5]
port 154 nsew signal output
rlabel metal2 s 30352 99600 30408 100000 6 reg_peri_addr[6]
port 155 nsew signal output
rlabel metal2 s 29792 99600 29848 100000 6 reg_peri_addr[7]
port 156 nsew signal output
rlabel metal2 s 29232 99600 29288 100000 6 reg_peri_addr[8]
port 157 nsew signal output
rlabel metal2 s 28672 99600 28728 100000 6 reg_peri_addr[9]
port 158 nsew signal output
rlabel metal2 s 35952 99600 36008 100000 6 reg_peri_be[0]
port 159 nsew signal output
rlabel metal2 s 35392 99600 35448 100000 6 reg_peri_be[1]
port 160 nsew signal output
rlabel metal2 s 34832 99600 34888 100000 6 reg_peri_be[2]
port 161 nsew signal output
rlabel metal2 s 34272 99600 34328 100000 6 reg_peri_be[3]
port 162 nsew signal output
rlabel metal2 s 26992 99600 27048 100000 6 reg_peri_cs
port 163 nsew signal output
rlabel metal2 s 71792 99600 71848 100000 6 reg_peri_rdata[0]
port 164 nsew signal input
rlabel metal2 s 66192 99600 66248 100000 6 reg_peri_rdata[10]
port 165 nsew signal input
rlabel metal2 s 65632 99600 65688 100000 6 reg_peri_rdata[11]
port 166 nsew signal input
rlabel metal2 s 65072 99600 65128 100000 6 reg_peri_rdata[12]
port 167 nsew signal input
rlabel metal2 s 64512 99600 64568 100000 6 reg_peri_rdata[13]
port 168 nsew signal input
rlabel metal2 s 63952 99600 64008 100000 6 reg_peri_rdata[14]
port 169 nsew signal input
rlabel metal2 s 63392 99600 63448 100000 6 reg_peri_rdata[15]
port 170 nsew signal input
rlabel metal2 s 62832 99600 62888 100000 6 reg_peri_rdata[16]
port 171 nsew signal input
rlabel metal2 s 62272 99600 62328 100000 6 reg_peri_rdata[17]
port 172 nsew signal input
rlabel metal2 s 61712 99600 61768 100000 6 reg_peri_rdata[18]
port 173 nsew signal input
rlabel metal2 s 61152 99600 61208 100000 6 reg_peri_rdata[19]
port 174 nsew signal input
rlabel metal2 s 71232 99600 71288 100000 6 reg_peri_rdata[1]
port 175 nsew signal input
rlabel metal2 s 60592 99600 60648 100000 6 reg_peri_rdata[20]
port 176 nsew signal input
rlabel metal2 s 60032 99600 60088 100000 6 reg_peri_rdata[21]
port 177 nsew signal input
rlabel metal2 s 59472 99600 59528 100000 6 reg_peri_rdata[22]
port 178 nsew signal input
rlabel metal2 s 58912 99600 58968 100000 6 reg_peri_rdata[23]
port 179 nsew signal input
rlabel metal2 s 58352 99600 58408 100000 6 reg_peri_rdata[24]
port 180 nsew signal input
rlabel metal2 s 57792 99600 57848 100000 6 reg_peri_rdata[25]
port 181 nsew signal input
rlabel metal2 s 57232 99600 57288 100000 6 reg_peri_rdata[26]
port 182 nsew signal input
rlabel metal2 s 56672 99600 56728 100000 6 reg_peri_rdata[27]
port 183 nsew signal input
rlabel metal2 s 56112 99600 56168 100000 6 reg_peri_rdata[28]
port 184 nsew signal input
rlabel metal2 s 55552 99600 55608 100000 6 reg_peri_rdata[29]
port 185 nsew signal input
rlabel metal2 s 70672 99600 70728 100000 6 reg_peri_rdata[2]
port 186 nsew signal input
rlabel metal2 s 54992 99600 55048 100000 6 reg_peri_rdata[30]
port 187 nsew signal input
rlabel metal2 s 54432 99600 54488 100000 6 reg_peri_rdata[31]
port 188 nsew signal input
rlabel metal2 s 70112 99600 70168 100000 6 reg_peri_rdata[3]
port 189 nsew signal input
rlabel metal2 s 69552 99600 69608 100000 6 reg_peri_rdata[4]
port 190 nsew signal input
rlabel metal2 s 68992 99600 69048 100000 6 reg_peri_rdata[5]
port 191 nsew signal input
rlabel metal2 s 68432 99600 68488 100000 6 reg_peri_rdata[6]
port 192 nsew signal input
rlabel metal2 s 67872 99600 67928 100000 6 reg_peri_rdata[7]
port 193 nsew signal input
rlabel metal2 s 67312 99600 67368 100000 6 reg_peri_rdata[8]
port 194 nsew signal input
rlabel metal2 s 66752 99600 66808 100000 6 reg_peri_rdata[9]
port 195 nsew signal input
rlabel metal2 s 53872 99600 53928 100000 6 reg_peri_wdata[0]
port 196 nsew signal output
rlabel metal2 s 48272 99600 48328 100000 6 reg_peri_wdata[10]
port 197 nsew signal output
rlabel metal2 s 47712 99600 47768 100000 6 reg_peri_wdata[11]
port 198 nsew signal output
rlabel metal2 s 47152 99600 47208 100000 6 reg_peri_wdata[12]
port 199 nsew signal output
rlabel metal2 s 46592 99600 46648 100000 6 reg_peri_wdata[13]
port 200 nsew signal output
rlabel metal2 s 46032 99600 46088 100000 6 reg_peri_wdata[14]
port 201 nsew signal output
rlabel metal2 s 45472 99600 45528 100000 6 reg_peri_wdata[15]
port 202 nsew signal output
rlabel metal2 s 44912 99600 44968 100000 6 reg_peri_wdata[16]
port 203 nsew signal output
rlabel metal2 s 44352 99600 44408 100000 6 reg_peri_wdata[17]
port 204 nsew signal output
rlabel metal2 s 43792 99600 43848 100000 6 reg_peri_wdata[18]
port 205 nsew signal output
rlabel metal2 s 43232 99600 43288 100000 6 reg_peri_wdata[19]
port 206 nsew signal output
rlabel metal2 s 53312 99600 53368 100000 6 reg_peri_wdata[1]
port 207 nsew signal output
rlabel metal2 s 42672 99600 42728 100000 6 reg_peri_wdata[20]
port 208 nsew signal output
rlabel metal2 s 42112 99600 42168 100000 6 reg_peri_wdata[21]
port 209 nsew signal output
rlabel metal2 s 41552 99600 41608 100000 6 reg_peri_wdata[22]
port 210 nsew signal output
rlabel metal2 s 40992 99600 41048 100000 6 reg_peri_wdata[23]
port 211 nsew signal output
rlabel metal2 s 40432 99600 40488 100000 6 reg_peri_wdata[24]
port 212 nsew signal output
rlabel metal2 s 39872 99600 39928 100000 6 reg_peri_wdata[25]
port 213 nsew signal output
rlabel metal2 s 39312 99600 39368 100000 6 reg_peri_wdata[26]
port 214 nsew signal output
rlabel metal2 s 38752 99600 38808 100000 6 reg_peri_wdata[27]
port 215 nsew signal output
rlabel metal2 s 38192 99600 38248 100000 6 reg_peri_wdata[28]
port 216 nsew signal output
rlabel metal2 s 37632 99600 37688 100000 6 reg_peri_wdata[29]
port 217 nsew signal output
rlabel metal2 s 52752 99600 52808 100000 6 reg_peri_wdata[2]
port 218 nsew signal output
rlabel metal2 s 37072 99600 37128 100000 6 reg_peri_wdata[30]
port 219 nsew signal output
rlabel metal2 s 36512 99600 36568 100000 6 reg_peri_wdata[31]
port 220 nsew signal output
rlabel metal2 s 52192 99600 52248 100000 6 reg_peri_wdata[3]
port 221 nsew signal output
rlabel metal2 s 51632 99600 51688 100000 6 reg_peri_wdata[4]
port 222 nsew signal output
rlabel metal2 s 51072 99600 51128 100000 6 reg_peri_wdata[5]
port 223 nsew signal output
rlabel metal2 s 50512 99600 50568 100000 6 reg_peri_wdata[6]
port 224 nsew signal output
rlabel metal2 s 49952 99600 50008 100000 6 reg_peri_wdata[7]
port 225 nsew signal output
rlabel metal2 s 49392 99600 49448 100000 6 reg_peri_wdata[8]
port 226 nsew signal output
rlabel metal2 s 48832 99600 48888 100000 6 reg_peri_wdata[9]
port 227 nsew signal output
rlabel metal2 s 27552 99600 27608 100000 6 reg_peri_wr
port 228 nsew signal output
rlabel metal3 s 0 96432 400 96488 6 reg_rdata[0]
port 229 nsew signal output
rlabel metal3 s 0 85232 400 85288 6 reg_rdata[10]
port 230 nsew signal output
rlabel metal3 s 0 84112 400 84168 6 reg_rdata[11]
port 231 nsew signal output
rlabel metal3 s 0 82992 400 83048 6 reg_rdata[12]
port 232 nsew signal output
rlabel metal3 s 0 81872 400 81928 6 reg_rdata[13]
port 233 nsew signal output
rlabel metal3 s 0 80752 400 80808 6 reg_rdata[14]
port 234 nsew signal output
rlabel metal3 s 0 79632 400 79688 6 reg_rdata[15]
port 235 nsew signal output
rlabel metal3 s 0 78512 400 78568 6 reg_rdata[16]
port 236 nsew signal output
rlabel metal3 s 0 77392 400 77448 6 reg_rdata[17]
port 237 nsew signal output
rlabel metal3 s 0 76272 400 76328 6 reg_rdata[18]
port 238 nsew signal output
rlabel metal3 s 0 75152 400 75208 6 reg_rdata[19]
port 239 nsew signal output
rlabel metal3 s 0 95312 400 95368 6 reg_rdata[1]
port 240 nsew signal output
rlabel metal3 s 0 74032 400 74088 6 reg_rdata[20]
port 241 nsew signal output
rlabel metal3 s 0 72912 400 72968 6 reg_rdata[21]
port 242 nsew signal output
rlabel metal3 s 0 71792 400 71848 6 reg_rdata[22]
port 243 nsew signal output
rlabel metal3 s 0 70672 400 70728 6 reg_rdata[23]
port 244 nsew signal output
rlabel metal3 s 0 69552 400 69608 6 reg_rdata[24]
port 245 nsew signal output
rlabel metal3 s 0 68432 400 68488 6 reg_rdata[25]
port 246 nsew signal output
rlabel metal3 s 0 67312 400 67368 6 reg_rdata[26]
port 247 nsew signal output
rlabel metal3 s 0 66192 400 66248 6 reg_rdata[27]
port 248 nsew signal output
rlabel metal3 s 0 65072 400 65128 6 reg_rdata[28]
port 249 nsew signal output
rlabel metal3 s 0 63952 400 64008 6 reg_rdata[29]
port 250 nsew signal output
rlabel metal3 s 0 94192 400 94248 6 reg_rdata[2]
port 251 nsew signal output
rlabel metal3 s 0 62832 400 62888 6 reg_rdata[30]
port 252 nsew signal output
rlabel metal3 s 0 61712 400 61768 6 reg_rdata[31]
port 253 nsew signal output
rlabel metal3 s 0 93072 400 93128 6 reg_rdata[3]
port 254 nsew signal output
rlabel metal3 s 0 91952 400 92008 6 reg_rdata[4]
port 255 nsew signal output
rlabel metal3 s 0 90832 400 90888 6 reg_rdata[5]
port 256 nsew signal output
rlabel metal3 s 0 89712 400 89768 6 reg_rdata[6]
port 257 nsew signal output
rlabel metal3 s 0 88592 400 88648 6 reg_rdata[7]
port 258 nsew signal output
rlabel metal3 s 0 87472 400 87528 6 reg_rdata[8]
port 259 nsew signal output
rlabel metal3 s 0 86352 400 86408 6 reg_rdata[9]
port 260 nsew signal output
rlabel metal3 s 0 60592 400 60648 6 reg_wdata[0]
port 261 nsew signal input
rlabel metal3 s 0 49392 400 49448 6 reg_wdata[10]
port 262 nsew signal input
rlabel metal3 s 0 48272 400 48328 6 reg_wdata[11]
port 263 nsew signal input
rlabel metal3 s 0 47152 400 47208 6 reg_wdata[12]
port 264 nsew signal input
rlabel metal3 s 0 46032 400 46088 6 reg_wdata[13]
port 265 nsew signal input
rlabel metal3 s 0 44912 400 44968 6 reg_wdata[14]
port 266 nsew signal input
rlabel metal3 s 0 43792 400 43848 6 reg_wdata[15]
port 267 nsew signal input
rlabel metal3 s 0 42672 400 42728 6 reg_wdata[16]
port 268 nsew signal input
rlabel metal3 s 0 41552 400 41608 6 reg_wdata[17]
port 269 nsew signal input
rlabel metal3 s 0 40432 400 40488 6 reg_wdata[18]
port 270 nsew signal input
rlabel metal3 s 0 39312 400 39368 6 reg_wdata[19]
port 271 nsew signal input
rlabel metal3 s 0 59472 400 59528 6 reg_wdata[1]
port 272 nsew signal input
rlabel metal3 s 0 38192 400 38248 6 reg_wdata[20]
port 273 nsew signal input
rlabel metal3 s 0 37072 400 37128 6 reg_wdata[21]
port 274 nsew signal input
rlabel metal3 s 0 35952 400 36008 6 reg_wdata[22]
port 275 nsew signal input
rlabel metal3 s 0 34832 400 34888 6 reg_wdata[23]
port 276 nsew signal input
rlabel metal3 s 0 33712 400 33768 6 reg_wdata[24]
port 277 nsew signal input
rlabel metal3 s 0 32592 400 32648 6 reg_wdata[25]
port 278 nsew signal input
rlabel metal3 s 0 31472 400 31528 6 reg_wdata[26]
port 279 nsew signal input
rlabel metal3 s 0 30352 400 30408 6 reg_wdata[27]
port 280 nsew signal input
rlabel metal3 s 0 29232 400 29288 6 reg_wdata[28]
port 281 nsew signal input
rlabel metal3 s 0 28112 400 28168 6 reg_wdata[29]
port 282 nsew signal input
rlabel metal3 s 0 58352 400 58408 6 reg_wdata[2]
port 283 nsew signal input
rlabel metal3 s 0 26992 400 27048 6 reg_wdata[30]
port 284 nsew signal input
rlabel metal3 s 0 25872 400 25928 6 reg_wdata[31]
port 285 nsew signal input
rlabel metal3 s 0 57232 400 57288 6 reg_wdata[3]
port 286 nsew signal input
rlabel metal3 s 0 56112 400 56168 6 reg_wdata[4]
port 287 nsew signal input
rlabel metal3 s 0 54992 400 55048 6 reg_wdata[5]
port 288 nsew signal input
rlabel metal3 s 0 53872 400 53928 6 reg_wdata[6]
port 289 nsew signal input
rlabel metal3 s 0 52752 400 52808 6 reg_wdata[7]
port 290 nsew signal input
rlabel metal3 s 0 51632 400 51688 6 reg_wdata[8]
port 291 nsew signal input
rlabel metal3 s 0 50512 400 50568 6 reg_wdata[9]
port 292 nsew signal input
rlabel metal3 s 0 7952 400 8008 6 reg_wr
port 293 nsew signal input
rlabel metal2 s 25872 99600 25928 100000 6 rtc_clk
port 294 nsew signal output
rlabel metal2 s 26432 99600 26488 100000 6 rtc_intr
port 295 nsew signal input
rlabel metal2 s 84896 0 84952 400 6 s_reset_n
port 296 nsew signal input
rlabel metal2 s 68432 0 68488 400 6 spim_miso
port 297 nsew signal input
rlabel metal2 s 70784 0 70840 400 6 spim_mosi
port 298 nsew signal output
rlabel metal2 s 56672 0 56728 400 6 spim_sck
port 299 nsew signal input
rlabel metal2 s 66080 0 66136 400 6 spim_ssn[0]
port 300 nsew signal input
rlabel metal2 s 63728 0 63784 400 6 spim_ssn[1]
port 301 nsew signal input
rlabel metal2 s 61376 0 61432 400 6 spim_ssn[2]
port 302 nsew signal input
rlabel metal2 s 59024 0 59080 400 6 spim_ssn[3]
port 303 nsew signal input
rlabel metal2 s 2576 0 2632 400 6 sspim_rst_n
port 304 nsew signal output
rlabel metal2 s 7280 0 7336 400 6 uart_rst_n[0]
port 305 nsew signal output
rlabel metal2 s 4928 0 4984 400 6 uart_rst_n[1]
port 306 nsew signal output
rlabel metal2 s 40208 0 40264 400 6 uart_rxd[0]
port 307 nsew signal output
rlabel metal2 s 35504 0 35560 400 6 uart_rxd[1]
port 308 nsew signal output
rlabel metal2 s 37856 0 37912 400 6 uart_txd[0]
port 309 nsew signal input
rlabel metal2 s 33152 0 33208 400 6 uart_txd[1]
port 310 nsew signal input
rlabel metal2 s 87248 0 87304 400 6 usb_clk
port 311 nsew signal output
rlabel metal2 s 30800 0 30856 400 6 usb_dn_i
port 312 nsew signal output
rlabel metal2 s 23744 0 23800 400 6 usb_dn_o
port 313 nsew signal input
rlabel metal2 s 28448 0 28504 400 6 usb_dp_i
port 314 nsew signal output
rlabel metal2 s 21392 0 21448 400 6 usb_dp_o
port 315 nsew signal input
rlabel metal2 s 77840 0 77896 400 6 usb_intr
port 316 nsew signal input
rlabel metal2 s 26096 0 26152 400 6 usb_oen
port 317 nsew signal input
rlabel metal2 s 11984 0 12040 400 6 usb_rst_n
port 318 nsew signal output
rlabel metal2 s 80192 0 80248 400 6 user_clock1
port 319 nsew signal input
rlabel metal2 s 82544 0 82600 400 6 user_clock2
port 320 nsew signal input
rlabel metal2 s 14336 0 14392 400 6 user_irq[0]
port 321 nsew signal output
rlabel metal2 s 16688 0 16744 400 6 user_irq[1]
port 322 nsew signal output
rlabel metal2 s 19040 0 19096 400 6 user_irq[2]
port 323 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 90000 100000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 29253984
string GDS_FILE /home/farag/carvel_riscv_soc/gf180mcu_riscv_soc/openlane/pinmux_top/runs/23_11_15_18_38/results/signoff/pinmux_top.magic.gds
string GDS_START 593340
<< end >>

