VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sar_adc
  CLASS BLOCK ;
  FOREIGN sar_adc ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 300.000 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 21.290 15.380 24.790 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 66.290 15.380 69.790 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 111.290 15.380 114.790 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 156.290 15.380 159.790 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 201.290 15.380 204.790 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 246.290 15.380 249.790 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 291.290 15.380 294.790 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 336.290 15.380 339.790 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 381.290 15.380 384.790 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 426.290 15.380 429.790 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 471.290 15.380 474.790 282.540 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 43.790 15.380 47.290 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 88.790 15.380 92.290 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 133.790 15.380 137.290 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 178.790 15.380 182.290 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 223.790 15.380 227.290 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 268.790 15.380 272.290 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 313.790 15.380 317.290 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 358.790 15.380 362.290 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 403.790 15.380 407.290 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 448.790 15.380 452.290 282.540 ;
    END
  END VSS
  PIN analog_dac_out
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 469.280 0.000 469.840 4.000 ;
    END
  END analog_dac_out
  PIN analog_din[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 414.400 0.000 414.960 4.000 ;
    END
  END analog_din[0]
  PIN analog_din[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 359.520 0.000 360.080 4.000 ;
    END
  END analog_din[1]
  PIN analog_din[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 304.640 0.000 305.200 4.000 ;
    END
  END analog_din[2]
  PIN analog_din[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 249.760 0.000 250.320 4.000 ;
    END
  END analog_din[3]
  PIN analog_din[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 194.880 0.000 195.440 4.000 ;
    END
  END analog_din[4]
  PIN analog_din[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 140.000 0.000 140.560 4.000 ;
    END
  END analog_din[5]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 11.020000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 20.160 4.000 20.720 ;
    END
  END clk
  PIN pulse1m_mclk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 85.120 0.000 85.680 4.000 ;
    END
  END pulse1m_mclk
  PIN reg_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 292.320 500.000 292.880 ;
    END
  END reg_ack
  PIN reg_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 76.160 4.000 76.720 ;
    END
  END reg_addr[0]
  PIN reg_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 70.560 4.000 71.120 ;
    END
  END reg_addr[1]
  PIN reg_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 64.960 4.000 65.520 ;
    END
  END reg_addr[2]
  PIN reg_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 59.360 4.000 59.920 ;
    END
  END reg_addr[3]
  PIN reg_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 53.760 4.000 54.320 ;
    END
  END reg_addr[4]
  PIN reg_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 48.160 4.000 48.720 ;
    END
  END reg_addr[5]
  PIN reg_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 42.560 4.000 43.120 ;
    END
  END reg_addr[6]
  PIN reg_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 36.960 4.000 37.520 ;
    END
  END reg_addr[7]
  PIN reg_be[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 98.560 4.000 99.120 ;
    END
  END reg_be[0]
  PIN reg_be[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 92.960 4.000 93.520 ;
    END
  END reg_be[1]
  PIN reg_be[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 87.360 4.000 87.920 ;
    END
  END reg_be[2]
  PIN reg_be[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 81.760 4.000 82.320 ;
    END
  END reg_be[3]
  PIN reg_cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 25.760 4.000 26.320 ;
    END
  END reg_cs
  PIN reg_rdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 283.360 500.000 283.920 ;
    END
  END reg_rdata[0]
  PIN reg_rdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 193.760 500.000 194.320 ;
    END
  END reg_rdata[10]
  PIN reg_rdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 184.800 500.000 185.360 ;
    END
  END reg_rdata[11]
  PIN reg_rdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 175.840 500.000 176.400 ;
    END
  END reg_rdata[12]
  PIN reg_rdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 166.880 500.000 167.440 ;
    END
  END reg_rdata[13]
  PIN reg_rdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 157.920 500.000 158.480 ;
    END
  END reg_rdata[14]
  PIN reg_rdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 148.960 500.000 149.520 ;
    END
  END reg_rdata[15]
  PIN reg_rdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 140.000 500.000 140.560 ;
    END
  END reg_rdata[16]
  PIN reg_rdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 131.040 500.000 131.600 ;
    END
  END reg_rdata[17]
  PIN reg_rdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 122.080 500.000 122.640 ;
    END
  END reg_rdata[18]
  PIN reg_rdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 113.120 500.000 113.680 ;
    END
  END reg_rdata[19]
  PIN reg_rdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 274.400 500.000 274.960 ;
    END
  END reg_rdata[1]
  PIN reg_rdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 104.160 500.000 104.720 ;
    END
  END reg_rdata[20]
  PIN reg_rdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 95.200 500.000 95.760 ;
    END
  END reg_rdata[21]
  PIN reg_rdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 86.240 500.000 86.800 ;
    END
  END reg_rdata[22]
  PIN reg_rdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 77.280 500.000 77.840 ;
    END
  END reg_rdata[23]
  PIN reg_rdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 68.320 500.000 68.880 ;
    END
  END reg_rdata[24]
  PIN reg_rdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 59.360 500.000 59.920 ;
    END
  END reg_rdata[25]
  PIN reg_rdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 50.400 500.000 50.960 ;
    END
  END reg_rdata[26]
  PIN reg_rdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 41.440 500.000 42.000 ;
    END
  END reg_rdata[27]
  PIN reg_rdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 32.480 500.000 33.040 ;
    END
  END reg_rdata[28]
  PIN reg_rdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 23.520 500.000 24.080 ;
    END
  END reg_rdata[29]
  PIN reg_rdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 265.440 500.000 266.000 ;
    END
  END reg_rdata[2]
  PIN reg_rdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 14.560 500.000 15.120 ;
    END
  END reg_rdata[30]
  PIN reg_rdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 5.600 500.000 6.160 ;
    END
  END reg_rdata[31]
  PIN reg_rdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 256.480 500.000 257.040 ;
    END
  END reg_rdata[3]
  PIN reg_rdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 247.520 500.000 248.080 ;
    END
  END reg_rdata[4]
  PIN reg_rdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 238.560 500.000 239.120 ;
    END
  END reg_rdata[5]
  PIN reg_rdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 229.600 500.000 230.160 ;
    END
  END reg_rdata[6]
  PIN reg_rdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 220.640 500.000 221.200 ;
    END
  END reg_rdata[7]
  PIN reg_rdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 211.680 500.000 212.240 ;
    END
  END reg_rdata[8]
  PIN reg_rdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal3 ;
        RECT 496.000 202.720 500.000 203.280 ;
    END
  END reg_rdata[9]
  PIN reg_wdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 277.760 4.000 278.320 ;
    END
  END reg_wdata[0]
  PIN reg_wdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 221.760 4.000 222.320 ;
    END
  END reg_wdata[10]
  PIN reg_wdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 216.160 4.000 216.720 ;
    END
  END reg_wdata[11]
  PIN reg_wdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 210.560 4.000 211.120 ;
    END
  END reg_wdata[12]
  PIN reg_wdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 204.960 4.000 205.520 ;
    END
  END reg_wdata[13]
  PIN reg_wdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 199.360 4.000 199.920 ;
    END
  END reg_wdata[14]
  PIN reg_wdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 193.760 4.000 194.320 ;
    END
  END reg_wdata[15]
  PIN reg_wdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 188.160 4.000 188.720 ;
    END
  END reg_wdata[16]
  PIN reg_wdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 182.560 4.000 183.120 ;
    END
  END reg_wdata[17]
  PIN reg_wdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 176.960 4.000 177.520 ;
    END
  END reg_wdata[18]
  PIN reg_wdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 171.360 4.000 171.920 ;
    END
  END reg_wdata[19]
  PIN reg_wdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 272.160 4.000 272.720 ;
    END
  END reg_wdata[1]
  PIN reg_wdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 165.760 4.000 166.320 ;
    END
  END reg_wdata[20]
  PIN reg_wdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 160.160 4.000 160.720 ;
    END
  END reg_wdata[21]
  PIN reg_wdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 154.560 4.000 155.120 ;
    END
  END reg_wdata[22]
  PIN reg_wdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 148.960 4.000 149.520 ;
    END
  END reg_wdata[23]
  PIN reg_wdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 143.360 4.000 143.920 ;
    END
  END reg_wdata[24]
  PIN reg_wdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 137.760 4.000 138.320 ;
    END
  END reg_wdata[25]
  PIN reg_wdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 132.160 4.000 132.720 ;
    END
  END reg_wdata[26]
  PIN reg_wdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 126.560 4.000 127.120 ;
    END
  END reg_wdata[27]
  PIN reg_wdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 120.960 4.000 121.520 ;
    END
  END reg_wdata[28]
  PIN reg_wdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 115.360 4.000 115.920 ;
    END
  END reg_wdata[29]
  PIN reg_wdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 266.560 4.000 267.120 ;
    END
  END reg_wdata[2]
  PIN reg_wdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 109.760 4.000 110.320 ;
    END
  END reg_wdata[30]
  PIN reg_wdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 104.160 4.000 104.720 ;
    END
  END reg_wdata[31]
  PIN reg_wdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 260.960 4.000 261.520 ;
    END
  END reg_wdata[3]
  PIN reg_wdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 255.360 4.000 255.920 ;
    END
  END reg_wdata[4]
  PIN reg_wdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 249.760 4.000 250.320 ;
    END
  END reg_wdata[5]
  PIN reg_wdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 244.160 4.000 244.720 ;
    END
  END reg_wdata[6]
  PIN reg_wdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 238.560 4.000 239.120 ;
    END
  END reg_wdata[7]
  PIN reg_wdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 232.960 4.000 233.520 ;
    END
  END reg_wdata[8]
  PIN reg_wdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 227.360 4.000 227.920 ;
    END
  END reg_wdata[9]
  PIN reg_wr
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 31.360 4.000 31.920 ;
    END
  END reg_wr
  PIN reset_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 30.240 0.000 30.800 4.000 ;
    END
  END reset_n
  PIN sar2dac[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 464.800 296.000 465.360 300.000 ;
    END
  END sar2dac[0]
  PIN sar2dac[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 403.200 296.000 403.760 300.000 ;
    END
  END sar2dac[1]
  PIN sar2dac[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 341.600 296.000 342.160 300.000 ;
    END
  END sar2dac[2]
  PIN sar2dac[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 280.000 296.000 280.560 300.000 ;
    END
  END sar2dac[3]
  PIN sar2dac[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 218.400 296.000 218.960 300.000 ;
    END
  END sar2dac[4]
  PIN sar2dac[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal2 ;
        RECT 156.800 296.000 157.360 300.000 ;
    END
  END sar2dac[5]
  PIN sar2dac[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 95.200 296.000 95.760 300.000 ;
    END
  END sar2dac[6]
  PIN sar2dac[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.986000 ;
    PORT
      LAYER Metal2 ;
        RECT 33.600 296.000 34.160 300.000 ;
    END
  END sar2dac[7]
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 492.800 283.210 ;
      LAYER Metal2 ;
        RECT 8.540 295.700 33.300 296.000 ;
        RECT 34.460 295.700 94.900 296.000 ;
        RECT 96.060 295.700 156.500 296.000 ;
        RECT 157.660 295.700 218.100 296.000 ;
        RECT 219.260 295.700 279.700 296.000 ;
        RECT 280.860 295.700 341.300 296.000 ;
        RECT 342.460 295.700 402.900 296.000 ;
        RECT 404.060 295.700 464.500 296.000 ;
        RECT 465.660 295.700 490.980 296.000 ;
        RECT 8.540 4.300 490.980 295.700 ;
        RECT 8.540 4.000 29.940 4.300 ;
        RECT 31.100 4.000 84.820 4.300 ;
        RECT 85.980 4.000 139.700 4.300 ;
        RECT 140.860 4.000 194.580 4.300 ;
        RECT 195.740 4.000 249.460 4.300 ;
        RECT 250.620 4.000 304.340 4.300 ;
        RECT 305.500 4.000 359.220 4.300 ;
        RECT 360.380 4.000 414.100 4.300 ;
        RECT 415.260 4.000 468.980 4.300 ;
        RECT 470.140 4.000 490.980 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 292.020 495.700 292.740 ;
        RECT 4.000 284.220 496.000 292.020 ;
        RECT 4.000 283.060 495.700 284.220 ;
        RECT 4.000 278.620 496.000 283.060 ;
        RECT 4.300 277.460 496.000 278.620 ;
        RECT 4.000 275.260 496.000 277.460 ;
        RECT 4.000 274.100 495.700 275.260 ;
        RECT 4.000 273.020 496.000 274.100 ;
        RECT 4.300 271.860 496.000 273.020 ;
        RECT 4.000 267.420 496.000 271.860 ;
        RECT 4.300 266.300 496.000 267.420 ;
        RECT 4.300 266.260 495.700 266.300 ;
        RECT 4.000 265.140 495.700 266.260 ;
        RECT 4.000 261.820 496.000 265.140 ;
        RECT 4.300 260.660 496.000 261.820 ;
        RECT 4.000 257.340 496.000 260.660 ;
        RECT 4.000 256.220 495.700 257.340 ;
        RECT 4.300 256.180 495.700 256.220 ;
        RECT 4.300 255.060 496.000 256.180 ;
        RECT 4.000 250.620 496.000 255.060 ;
        RECT 4.300 249.460 496.000 250.620 ;
        RECT 4.000 248.380 496.000 249.460 ;
        RECT 4.000 247.220 495.700 248.380 ;
        RECT 4.000 245.020 496.000 247.220 ;
        RECT 4.300 243.860 496.000 245.020 ;
        RECT 4.000 239.420 496.000 243.860 ;
        RECT 4.300 238.260 495.700 239.420 ;
        RECT 4.000 233.820 496.000 238.260 ;
        RECT 4.300 232.660 496.000 233.820 ;
        RECT 4.000 230.460 496.000 232.660 ;
        RECT 4.000 229.300 495.700 230.460 ;
        RECT 4.000 228.220 496.000 229.300 ;
        RECT 4.300 227.060 496.000 228.220 ;
        RECT 4.000 222.620 496.000 227.060 ;
        RECT 4.300 221.500 496.000 222.620 ;
        RECT 4.300 221.460 495.700 221.500 ;
        RECT 4.000 220.340 495.700 221.460 ;
        RECT 4.000 217.020 496.000 220.340 ;
        RECT 4.300 215.860 496.000 217.020 ;
        RECT 4.000 212.540 496.000 215.860 ;
        RECT 4.000 211.420 495.700 212.540 ;
        RECT 4.300 211.380 495.700 211.420 ;
        RECT 4.300 210.260 496.000 211.380 ;
        RECT 4.000 205.820 496.000 210.260 ;
        RECT 4.300 204.660 496.000 205.820 ;
        RECT 4.000 203.580 496.000 204.660 ;
        RECT 4.000 202.420 495.700 203.580 ;
        RECT 4.000 200.220 496.000 202.420 ;
        RECT 4.300 199.060 496.000 200.220 ;
        RECT 4.000 194.620 496.000 199.060 ;
        RECT 4.300 193.460 495.700 194.620 ;
        RECT 4.000 189.020 496.000 193.460 ;
        RECT 4.300 187.860 496.000 189.020 ;
        RECT 4.000 185.660 496.000 187.860 ;
        RECT 4.000 184.500 495.700 185.660 ;
        RECT 4.000 183.420 496.000 184.500 ;
        RECT 4.300 182.260 496.000 183.420 ;
        RECT 4.000 177.820 496.000 182.260 ;
        RECT 4.300 176.700 496.000 177.820 ;
        RECT 4.300 176.660 495.700 176.700 ;
        RECT 4.000 175.540 495.700 176.660 ;
        RECT 4.000 172.220 496.000 175.540 ;
        RECT 4.300 171.060 496.000 172.220 ;
        RECT 4.000 167.740 496.000 171.060 ;
        RECT 4.000 166.620 495.700 167.740 ;
        RECT 4.300 166.580 495.700 166.620 ;
        RECT 4.300 165.460 496.000 166.580 ;
        RECT 4.000 161.020 496.000 165.460 ;
        RECT 4.300 159.860 496.000 161.020 ;
        RECT 4.000 158.780 496.000 159.860 ;
        RECT 4.000 157.620 495.700 158.780 ;
        RECT 4.000 155.420 496.000 157.620 ;
        RECT 4.300 154.260 496.000 155.420 ;
        RECT 4.000 149.820 496.000 154.260 ;
        RECT 4.300 148.660 495.700 149.820 ;
        RECT 4.000 144.220 496.000 148.660 ;
        RECT 4.300 143.060 496.000 144.220 ;
        RECT 4.000 140.860 496.000 143.060 ;
        RECT 4.000 139.700 495.700 140.860 ;
        RECT 4.000 138.620 496.000 139.700 ;
        RECT 4.300 137.460 496.000 138.620 ;
        RECT 4.000 133.020 496.000 137.460 ;
        RECT 4.300 131.900 496.000 133.020 ;
        RECT 4.300 131.860 495.700 131.900 ;
        RECT 4.000 130.740 495.700 131.860 ;
        RECT 4.000 127.420 496.000 130.740 ;
        RECT 4.300 126.260 496.000 127.420 ;
        RECT 4.000 122.940 496.000 126.260 ;
        RECT 4.000 121.820 495.700 122.940 ;
        RECT 4.300 121.780 495.700 121.820 ;
        RECT 4.300 120.660 496.000 121.780 ;
        RECT 4.000 116.220 496.000 120.660 ;
        RECT 4.300 115.060 496.000 116.220 ;
        RECT 4.000 113.980 496.000 115.060 ;
        RECT 4.000 112.820 495.700 113.980 ;
        RECT 4.000 110.620 496.000 112.820 ;
        RECT 4.300 109.460 496.000 110.620 ;
        RECT 4.000 105.020 496.000 109.460 ;
        RECT 4.300 103.860 495.700 105.020 ;
        RECT 4.000 99.420 496.000 103.860 ;
        RECT 4.300 98.260 496.000 99.420 ;
        RECT 4.000 96.060 496.000 98.260 ;
        RECT 4.000 94.900 495.700 96.060 ;
        RECT 4.000 93.820 496.000 94.900 ;
        RECT 4.300 92.660 496.000 93.820 ;
        RECT 4.000 88.220 496.000 92.660 ;
        RECT 4.300 87.100 496.000 88.220 ;
        RECT 4.300 87.060 495.700 87.100 ;
        RECT 4.000 85.940 495.700 87.060 ;
        RECT 4.000 82.620 496.000 85.940 ;
        RECT 4.300 81.460 496.000 82.620 ;
        RECT 4.000 78.140 496.000 81.460 ;
        RECT 4.000 77.020 495.700 78.140 ;
        RECT 4.300 76.980 495.700 77.020 ;
        RECT 4.300 75.860 496.000 76.980 ;
        RECT 4.000 71.420 496.000 75.860 ;
        RECT 4.300 70.260 496.000 71.420 ;
        RECT 4.000 69.180 496.000 70.260 ;
        RECT 4.000 68.020 495.700 69.180 ;
        RECT 4.000 65.820 496.000 68.020 ;
        RECT 4.300 64.660 496.000 65.820 ;
        RECT 4.000 60.220 496.000 64.660 ;
        RECT 4.300 59.060 495.700 60.220 ;
        RECT 4.000 54.620 496.000 59.060 ;
        RECT 4.300 53.460 496.000 54.620 ;
        RECT 4.000 51.260 496.000 53.460 ;
        RECT 4.000 50.100 495.700 51.260 ;
        RECT 4.000 49.020 496.000 50.100 ;
        RECT 4.300 47.860 496.000 49.020 ;
        RECT 4.000 43.420 496.000 47.860 ;
        RECT 4.300 42.300 496.000 43.420 ;
        RECT 4.300 42.260 495.700 42.300 ;
        RECT 4.000 41.140 495.700 42.260 ;
        RECT 4.000 37.820 496.000 41.140 ;
        RECT 4.300 36.660 496.000 37.820 ;
        RECT 4.000 33.340 496.000 36.660 ;
        RECT 4.000 32.220 495.700 33.340 ;
        RECT 4.300 32.180 495.700 32.220 ;
        RECT 4.300 31.060 496.000 32.180 ;
        RECT 4.000 26.620 496.000 31.060 ;
        RECT 4.300 25.460 496.000 26.620 ;
        RECT 4.000 24.380 496.000 25.460 ;
        RECT 4.000 23.220 495.700 24.380 ;
        RECT 4.000 21.020 496.000 23.220 ;
        RECT 4.300 19.860 496.000 21.020 ;
        RECT 4.000 15.420 496.000 19.860 ;
        RECT 4.000 14.260 495.700 15.420 ;
        RECT 4.000 6.460 496.000 14.260 ;
        RECT 4.000 5.740 495.700 6.460 ;
      LAYER Metal4 ;
        RECT 244.300 21.930 245.990 210.470 ;
        RECT 250.090 21.930 268.490 210.470 ;
        RECT 272.590 21.930 290.990 210.470 ;
        RECT 295.090 21.930 313.490 210.470 ;
        RECT 317.590 21.930 335.990 210.470 ;
        RECT 340.090 21.930 358.490 210.470 ;
        RECT 362.590 21.930 378.420 210.470 ;
      LAYER Metal5 ;
        RECT 297.980 24.530 378.500 24.970 ;
  END
END sar_adc
END LIBRARY

