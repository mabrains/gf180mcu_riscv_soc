module DSM_core (clk,
    i_wb_cyc,
    i_wb_stb,
    i_wb_we,
    o_wb_ack,
    o_wb_stall,
    reset,
    vdd,
    vss,
    i_wb_addr,
    i_wb_data,
    o_wb_data);
 input clk;
 input i_wb_cyc;
 input i_wb_stb;
 input i_wb_we;
 output o_wb_ack;
 output o_wb_stall;
 input reset;
 input vdd;
 input vss;
 input [31:0] i_wb_addr;
 input [6:0] i_wb_data;
 output [4:0] o_wb_data;

 wire net82;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire \d1.Cout ;
 wire \d1.In_Data[0] ;
 wire \d1.In_Data[1] ;
 wire \d1.In_Data[2] ;
 wire \d1.In_Data[3] ;
 wire \d1.In_Data[4] ;
 wire \d1.In_Data[5] ;
 wire \d1.In_Data[6] ;
 wire \d1.Out_Data[0] ;
 wire \d1.Out_Data[1] ;
 wire \d1.Out_Data[2] ;
 wire \d1.Out_Data[3] ;
 wire \d1.Out_Data[4] ;
 wire \d1.Out_Data[5] ;
 wire \d1.Out_Data[6] ;
 wire \d1.Sum[0] ;
 wire \d1.Sum[1] ;
 wire \d1.Sum[2] ;
 wire \d1.Sum[3] ;
 wire \d1.Sum[4] ;
 wire \d1.Sum[5] ;
 wire \d1.Sum[6] ;
 wire \d1._00_ ;
 wire \d1._01_ ;
 wire \d1._02_ ;
 wire \d1._03_ ;
 wire \d1._04_ ;
 wire \d1._05_ ;
 wire \d1._06_ ;
 wire \d1._07_ ;
 wire \d1._08_ ;
 wire \d1._09_ ;
 wire \d1._10_ ;
 wire \d1._11_ ;
 wire \d1._12_ ;
 wire \d1._13_ ;
 wire \d1._14_ ;
 wire \d1._15_ ;
 wire \d1._16_ ;
 wire \d1._17_ ;
 wire \d1._18_ ;
 wire \d1._19_ ;
 wire \d1._20_ ;
 wire \d1._21_ ;
 wire \d1._22_ ;
 wire \d1._23_ ;
 wire \d1._24_ ;
 wire \d1._25_ ;
 wire \d1._26_ ;
 wire \d1._27_ ;
 wire \d1._28_ ;
 wire \d1._29_ ;
 wire \d1._30_ ;
 wire \d1._31_ ;
 wire \d1._32_ ;
 wire \d1._33_ ;
 wire \d1._34_ ;
 wire \d1._35_ ;
 wire \d1._36_ ;
 wire \d1._37_ ;
 wire \d2.Cout ;
 wire \d2.Out_Data[0] ;
 wire \d2.Out_Data[1] ;
 wire \d2.Out_Data[2] ;
 wire \d2.Out_Data[3] ;
 wire \d2.Out_Data[4] ;
 wire \d2.Out_Data[5] ;
 wire \d2.Out_Data[6] ;
 wire \d2.Sum[0] ;
 wire \d2.Sum[1] ;
 wire \d2.Sum[2] ;
 wire \d2.Sum[3] ;
 wire \d2.Sum[4] ;
 wire \d2.Sum[5] ;
 wire \d2.Sum[6] ;
 wire \d2._00_ ;
 wire \d2._01_ ;
 wire \d2._02_ ;
 wire \d2._03_ ;
 wire \d2._04_ ;
 wire \d2._05_ ;
 wire \d2._06_ ;
 wire \d2._07_ ;
 wire \d2._08_ ;
 wire \d2._09_ ;
 wire \d2._10_ ;
 wire \d2._11_ ;
 wire \d2._12_ ;
 wire \d2._13_ ;
 wire \d2._14_ ;
 wire \d2._15_ ;
 wire \d2._16_ ;
 wire \d2._17_ ;
 wire \d2._18_ ;
 wire \d2._19_ ;
 wire \d2._20_ ;
 wire \d2._21_ ;
 wire \d2._22_ ;
 wire \d2._23_ ;
 wire \d2._24_ ;
 wire \d2._25_ ;
 wire \d2._26_ ;
 wire \d2._27_ ;
 wire \d2._28_ ;
 wire \d2._29_ ;
 wire \d2._30_ ;
 wire \d2._31_ ;
 wire \d2._32_ ;
 wire \d2._33_ ;
 wire \d2._34_ ;
 wire \d2._35_ ;
 wire \d2._36_ ;
 wire \d2._37_ ;
 wire \d3.Cout ;
 wire \d3.Out_Data[0] ;
 wire \d3.Out_Data[1] ;
 wire \d3.Out_Data[2] ;
 wire \d3.Out_Data[3] ;
 wire \d3.Out_Data[4] ;
 wire \d3.Out_Data[5] ;
 wire \d3.Out_Data[6] ;
 wire \d3.Sum[0] ;
 wire \d3.Sum[1] ;
 wire \d3.Sum[2] ;
 wire \d3.Sum[3] ;
 wire \d3.Sum[4] ;
 wire \d3.Sum[5] ;
 wire \d3.Sum[6] ;
 wire \d3._00_ ;
 wire \d3._01_ ;
 wire \d3._02_ ;
 wire \d3._03_ ;
 wire \d3._04_ ;
 wire \d3._05_ ;
 wire \d3._06_ ;
 wire \d3._07_ ;
 wire \d3._08_ ;
 wire \d3._09_ ;
 wire \d3._10_ ;
 wire \d3._11_ ;
 wire \d3._12_ ;
 wire \d3._13_ ;
 wire \d3._14_ ;
 wire \d3._15_ ;
 wire \d3._16_ ;
 wire \d3._17_ ;
 wire \d3._18_ ;
 wire \d3._19_ ;
 wire \d3._20_ ;
 wire \d3._21_ ;
 wire \d3._22_ ;
 wire \d3._23_ ;
 wire \d3._24_ ;
 wire \d3._25_ ;
 wire \d3._26_ ;
 wire \d3._27_ ;
 wire \d3._28_ ;
 wire \d3._29_ ;
 wire \d3._30_ ;
 wire \d3._31_ ;
 wire \d3._32_ ;
 wire \d3._33_ ;
 wire \d3._34_ ;
 wire \d3._35_ ;
 wire \d3._36_ ;
 wire \d3._37_ ;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net9;
 wire \u4.Data3[0] ;
 wire \u4.Out_Data[0] ;
 wire \u4.Out_Data[1] ;
 wire \u4.Out_Data[2] ;
 wire \u4.Out_Data[3] ;
 wire \u4.Out_Data[4] ;
 wire \u4._00_ ;
 wire \u4._01_ ;
 wire \u4._02_ ;
 wire \u4._03_ ;
 wire \u4._04_ ;
 wire \u4._05_ ;
 wire \u4._06_ ;
 wire \u4._07_ ;
 wire \u4._08_ ;
 wire \u4._09_ ;
 wire \u4._10_ ;
 wire \u4._11_ ;
 wire \u4._12_ ;
 wire \u4._13_ ;
 wire \u4._14_ ;
 wire \u4._15_ ;
 wire \u4._16_ ;
 wire \u4._17_ ;
 wire \u4._18_ ;
 wire \u4._19_ ;
 wire \u4._20_ ;
 wire \u4._21_ ;
 wire \u4._22_ ;
 wire \u4._23_ ;
 wire \u4._24_ ;
 wire \u4._25_ ;
 wire \u4._26_ ;
 wire \u4._27_ ;
 wire \u4._28_ ;
 wire \u4._29_ ;
 wire \u4._30_ ;
 wire \u4._31_ ;
 wire \u4._32_ ;
 wire \u5.Data3[0] ;
 wire \u5.Data3[1] ;
 wire \u5.Data3[2] ;
 wire \u5.Data3[3] ;
 wire \u5.Data3[4] ;
 wire \u5.Out_Data[0] ;
 wire \u5.Out_Data[1] ;
 wire \u5.Out_Data[2] ;
 wire \u5.Out_Data[3] ;
 wire \u5.Out_Data[4] ;
 wire \u5._00_ ;
 wire \u5._01_ ;
 wire \u5._02_ ;
 wire \u5._03_ ;
 wire \u5._04_ ;
 wire \u5._05_ ;
 wire \u5._06_ ;
 wire \u5._07_ ;
 wire \u5._08_ ;
 wire \u5._09_ ;
 wire \u5._10_ ;
 wire \u5._11_ ;
 wire \u5._12_ ;
 wire \u5._13_ ;
 wire \u5._14_ ;
 wire \u5._15_ ;
 wire \u5._16_ ;
 wire \u5._17_ ;
 wire \u5._18_ ;
 wire \u5._19_ ;
 wire \u5._20_ ;
 wire \u5._21_ ;
 wire \u5._22_ ;
 wire \u5._23_ ;
 wire \u5._24_ ;
 wire \u5._25_ ;
 wire \u5._26_ ;
 wire \u5._27_ ;
 wire \u5._28_ ;
 wire \u5._29_ ;
 wire \u5._30_ ;
 wire \u5._31_ ;
 wire \u5._32_ ;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__081__I (.I(net44),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__098__A2 (.I(_050_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__099__A2 (.I(_041_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__099__A3 (.I(_049_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__099__A4 (.I(_057_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__104__A1 (.I(_050_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__106__A2 (.I(_063_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__106__B (.I(\d1.In_Data[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__107__A1 (.I(_050_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__111__A2 (.I(_063_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__111__B (.I(\d1.In_Data[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__114__A2 (.I(_063_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__114__B (.I(\d1.In_Data[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__117__A2 (.I(_063_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__120__A2 (.I(_063_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__123__A2 (.I(_063_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__126__A2 (.I(_063_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__131__A2 (.I(_049_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__131__A3 (.I(_057_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__132__A2 (.I(_029_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__132__B (.I(_041_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__133__A1 (.I(_029_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__134__A2 (.I(_049_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__134__A3 (.I(_057_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__135__A2 (.I(_029_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__135__B (.I(_041_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__136__A1 (.I(_029_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__137__A2 (.I(_049_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__137__A3 (.I(_057_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__138__A2 (.I(_029_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__138__B (.I(_041_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__139__A1 (.I(_029_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__140__A2 (.I(_049_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__140__A3 (.I(_057_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__141__A2 (.I(_029_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__141__B (.I(_041_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__142__A1 (.I(_029_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__143__A2 (.I(_049_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__143__A3 (.I(_057_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__144__A2 (.I(_029_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__144__B (.I(_041_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__145__A1 (.I(_029_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__146__CLK (.I(clknet_2_0__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__147__CLK (.I(clknet_2_0__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__147__RN (.I(net44),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__148__CLK (.I(clknet_2_0__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__148__RN (.I(net44),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__149__CLK (.I(clknet_2_0__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__149__RN (.I(net44),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__150__CLK (.I(clknet_2_2__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__150__RN (.I(net44),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__151__CLK (.I(clknet_2_2__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__151__RN (.I(net44),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__152__CLK (.I(clknet_2_2__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__152__RN (.I(net44),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__153__CLK (.I(clknet_2_0__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__154__CLK (.I(clknet_2_0__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__155__CLK (.I(clknet_2_0__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__156__CLK (.I(clknet_2_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__157__CLK (.I(clknet_2_0__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__158__CLK (.I(clknet_2_0__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__159__CLK (.I(clknet_2_0__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__160__CLK (.I(clknet_2_0__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__161__CLK (.I(clknet_2_0__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__162__CLK (.I(clknet_2_2__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__163__CLK (.I(clknet_2_2__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__164__CLK (.I(clknet_2_2__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_clk_I (.I(clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_0__f_clk_I (.I(clknet_0_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_1__f_clk_I (.I(clknet_0_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_2__f_clk_I (.I(clknet_0_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_3__f_clk_I (.I(clknet_0_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d1._38__A2  (.I(\d1.In_Data[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d1._39__A2  (.I(\d1.In_Data[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d1._41__A2  (.I(\d1.In_Data[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d1._42__A2  (.I(\d1.In_Data[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d1._43__A2  (.I(\d1.In_Data[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d1._45__A2  (.I(\d1.In_Data[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d1._48__A2  (.I(\d1.In_Data[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d1._56__C  (.I(\d1.In_Data[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d1._67__A2  (.I(\d1.In_Data[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d1._68__A2  (.I(\d1.In_Data[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d1._79__A2  (.I(\d1.In_Data[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d1._84__CLK  (.I(clknet_2_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d1._84__RN  (.I(net44),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d1._85__CLK  (.I(clknet_2_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d1._85__RN  (.I(net44),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d1._86__CLK  (.I(clknet_2_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d1._86__RN  (.I(net44),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d1._87__CLK  (.I(clknet_2_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d1._87__RN  (.I(net44),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d1._88__CLK  (.I(clknet_2_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d1._88__RN  (.I(net44),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d1._89__CLK  (.I(clknet_2_0__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d1._89__RN  (.I(net44),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d1._90__CLK  (.I(clknet_2_0__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d1._90__RN  (.I(net44),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d2._84__CLK  (.I(clknet_2_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d2._84__RN  (.I(net44),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d2._85__CLK  (.I(clknet_2_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d2._85__RN  (.I(net44),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d2._86__CLK  (.I(clknet_2_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d2._86__RN  (.I(net43),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d2._87__CLK  (.I(clknet_2_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d2._87__RN  (.I(net43),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d2._88__CLK  (.I(clknet_2_3__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d2._88__RN  (.I(net43),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d2._89__CLK  (.I(clknet_2_3__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d2._89__RN  (.I(net44),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d2._90__CLK  (.I(clknet_2_2__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d2._90__RN  (.I(net44),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d3._84__CLK  (.I(clknet_2_3__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d3._84__RN  (.I(net43),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d3._85__CLK  (.I(clknet_2_3__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d3._85__RN  (.I(net43),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d3._86__CLK  (.I(clknet_2_3__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d3._86__RN  (.I(net43),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d3._87__CLK  (.I(clknet_2_3__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d3._87__RN  (.I(net43),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d3._88__CLK  (.I(clknet_2_3__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d3._88__RN  (.I(net43),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d3._89__CLK  (.I(clknet_2_3__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d3._89__RN  (.I(net44),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d3._90__CLK  (.I(clknet_2_3__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_d3._90__RN  (.I(net44),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout44_I (.I(net43),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(i_wb_addr[18]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(i_wb_addr[19]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(i_wb_addr[1]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(i_wb_addr[20]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(i_wb_addr[21]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(i_wb_addr[22]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(i_wb_addr[23]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(i_wb_addr[24]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(i_wb_addr[25]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(i_wb_addr[26]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(i_wb_addr[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(i_wb_addr[27]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(i_wb_addr[28]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(i_wb_addr[29]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(i_wb_addr[2]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(i_wb_addr[30]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(i_wb_addr[31]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(i_wb_addr[3]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(i_wb_addr[4]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(i_wb_addr[5]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(i_wb_addr[6]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(i_wb_addr[10]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(i_wb_addr[7]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(i_wb_addr[8]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(i_wb_addr[9]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(i_wb_cyc),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input34_I (.I(i_wb_data[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input35_I (.I(i_wb_data[1]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input36_I (.I(i_wb_data[2]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input37_I (.I(i_wb_data[3]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input38_I (.I(i_wb_data[4]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input39_I (.I(i_wb_data[5]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(i_wb_addr[11]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input40_I (.I(i_wb_data[6]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input41_I (.I(i_wb_stb),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input42_I (.I(i_wb_we),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input43_I (.I(reset),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(i_wb_addr[12]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(i_wb_addr[13]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(i_wb_addr[14]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(i_wb_addr[15]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(i_wb_addr[16]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(i_wb_addr[17]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel DSM_core_82 (.ZN(net82),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_12 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_16 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_188 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_196 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_200 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_240 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_248 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_252 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_254 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_257 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_265 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_269 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_271 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_308 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_324 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_328 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_330 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_36 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_46 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_50 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_74 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_90 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_98 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_113 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_145 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_161 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_165 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_167 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_19 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_197 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_199 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_224 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_228 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_267 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_280 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_31 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_312 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_14 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_166 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_170 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_214 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_330 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_48 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_52 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_68 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_121 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_153 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_169 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_19 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_201 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_208 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_237 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_27 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_271 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_31 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_323 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_49 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_81 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_97 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_12 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_146 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_150 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_156 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_16 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_163 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_204 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_208 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_220 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_224 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_226 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_233 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_265 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_273 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_298 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_302 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_304 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_328 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_330 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_48 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_64 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_68 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_102 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_115 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_131 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_135 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_149 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_185 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_19 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_225 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_229 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_23 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_231 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_255 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_31 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_78 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_82 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_86 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_94 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_133 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_203 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_226 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_234 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_238 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_28 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_292 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_296 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_316 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_324 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_328 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_330 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_44 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_62 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_82 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_115 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_155 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_19 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_23 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_232 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_240 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_255 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_257 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_269 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_27 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_285 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_49 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_51 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_54 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_86 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_95 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_118 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_224 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_272 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_294 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_30 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_315 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_46 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_50 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_60 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_68 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_76 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_78 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_12 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_14 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_224 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_240 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_31 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_49 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_84 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_97 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_112 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_118 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_12 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_124 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_15 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_200 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_208 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_248 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_270 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_330 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_43 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_47 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_51 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_63 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_115 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_119 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_135 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_146 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_148 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_151 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_163 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_187 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_220 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_224 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_226 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_267 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_271 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_330 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_43 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_57 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_61 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_74 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_77 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_188 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_192 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_233 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_237 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_41 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_252 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_272 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_330 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_47 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_63 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_12 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_129 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_133 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_141 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_149 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_153 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_155 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_170 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_227 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_231 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_239 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_243 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_28 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_85 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_95 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_12 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_125 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_127 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_194 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_198 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_202 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_224 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_232 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_236 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_271 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_275 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_330 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_51 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_55 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_57 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_86 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_88 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_115 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_119 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_12 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_167 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_28 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_294 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_310 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_57 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_114 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_12 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_130 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_132 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_148 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_180 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_196 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_218 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_231 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_273 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_330 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_49 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_57 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_61 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_63 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_82 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_131 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_133 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_154 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_170 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_196 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_214 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_223 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_23 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_239 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_243 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_31 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_61 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_63 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_85 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_124 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_128 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_132 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_134 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_155 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_159 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_194 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_196 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_217 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_230 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_262 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_330 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_77 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_85 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_89 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_12 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_155 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_170 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_195 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_198 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_230 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_240 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_28 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_281 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_285 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_289 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_305 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_85 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_95 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_12 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_120 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_128 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_16 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_330 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_61 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_181 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_219 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_223 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_231 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_233 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_255 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_301 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_309 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_33 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_75 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_79 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_82 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_94 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_12 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_160 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_163 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_201 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_226 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_26 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_297 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_91 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_99 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_101 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_109 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_113 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_146 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_148 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_161 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_203 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_225 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_239 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_243 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_245 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_322 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_330 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_42 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_44 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_85 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_157 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_161 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_168 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_195 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_22 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_259 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_291 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_30 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_307 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_49 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_51 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_87 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_118 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_12 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_122 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_126 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_155 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_16 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_187 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_203 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_207 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_245 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_254 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_270 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_330 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_44 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_52 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_56 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_62 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_12 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_165 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_173 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_225 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_28 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_73 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_109 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_125 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_133 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_152 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_160 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_162 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_201 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_322 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_326 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_328 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_47 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_49 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_77 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_12 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_127 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_140 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_168 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_221 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_237 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_28 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_281 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_285 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_289 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_305 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_57 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_59 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_119 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_12 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_127 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_135 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_220 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_236 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_238 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_245 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_330 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_44 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_60 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_68 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_76 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_102 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_12 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_131 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_170 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_213 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_227 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_243 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_28 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_74 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_90 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_98 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_112 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_116 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_118 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_12 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_157 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_199 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_203 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_234 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_266 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_330 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_44 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_14 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_156 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_194 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_220 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_222 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_225 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_229 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_238 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_245 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_250 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_254 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_256 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_259 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_269 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_277 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_279 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_330 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_46 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_62 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_74 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_84 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_92 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_95 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_131 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_135 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_158 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_160 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_167 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_226 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_23 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_31 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_47 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_12 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_120 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_124 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_128 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_132 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_134 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_16 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_165 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_197 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_205 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_330 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_12 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_131 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_135 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_160 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_168 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_193 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_201 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_210 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_234 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_28 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_34 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_45 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_49 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_60 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_76 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_87 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_148 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_164 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_176 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_184 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_198 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_220 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_224 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_260 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_264 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_268 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_330 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_50 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_6 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_60 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_68 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_127 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_211 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_215 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_219 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_227 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_235 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_243 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_91 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_95 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_99 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_12 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_136 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_182 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_190 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_276 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_314 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_330 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_44 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_52 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_56 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_59 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_104 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_14 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_206 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_22 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_240 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_30 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_308 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_324 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_328 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_330 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_36 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_70 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_118 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_12 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_126 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_130 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_133 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_144 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_160 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_168 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_17 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_172 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_174 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_225 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_229 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_236 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_240 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_242 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_249 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_257 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_261 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_293 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_301 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_309 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_313 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_33 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_41 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_49 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_61 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_83 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_99 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_105 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_124 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_18 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_186 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_202 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_222 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_254 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_270 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_298 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_327 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_56 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_60 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_68 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_74 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_87 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_95 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_99 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_123 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_155 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_171 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_179 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_197 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_232 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_240 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_244 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_263 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_267 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_292 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_300 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_304 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_306 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_311 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_53 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_57 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_89 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_105 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_110 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_126 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_134 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_138 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_170 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_2 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_202 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_227 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_229 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_234 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_266 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_274 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_278 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_298 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_302 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_327 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_4 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_63 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_67 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_69 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_72 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_76 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_92 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_103 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_107 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_111 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_14 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_177 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_241 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_247 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_290 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_294 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_310 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_317 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_325 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_329 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_33 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_37 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_10 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_100 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_102 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_105 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_137 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_139 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_142 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_150 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_152 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_169 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_201 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_209 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_212 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_228 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_236 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_282 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_286 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_292 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_32 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_328 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_330 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_36 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_46 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_58 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_66 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_8 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_80 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_84 (.VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_47 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_57 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_58 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_59 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_60 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_61 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_62 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_63 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_64 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_65 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_66 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_48 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_67 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_68 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_69 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_70 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_71 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_72 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_73 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_74 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_75 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_76 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_49 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_77 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_78 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_79 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_80 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_81 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_82 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_83 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_84 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_85 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_86 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_50 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_87 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_88 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_89 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_90 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_91 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Left_92 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Right_45 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Left_93 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Right_46 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_51 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_52 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_53 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_54 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_55 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_56 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_100 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_101 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_102 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_94 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_95 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_96 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_97 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_98 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_99 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_143 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_144 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_145 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_146 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_147 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_148 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_149 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_150 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_151 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_152 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_153 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_154 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_155 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_156 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_157 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_158 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_159 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_160 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_161 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_162 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_163 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_164 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_165 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_166 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_167 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_168 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_169 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_170 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_171 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_172 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_173 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_174 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_175 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_176 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_177 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_178 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_179 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_180 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_181 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_182 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_183 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_184 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_185 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_186 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_187 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_103 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_104 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_105 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_106 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_188 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_189 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_190 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_191 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_192 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_193 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_194 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_195 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_196 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_197 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_198 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_199 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_200 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_201 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_202 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_203 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_204 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_205 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_206 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_207 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_208 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_209 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_210 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_211 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_212 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_213 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_214 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_215 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_216 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_217 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_218 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_219 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_220 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_221 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_222 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_223 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_224 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_225 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_226 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_227 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_228 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_229 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_230 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_231 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_232 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_107 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_108 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_109 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_110 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_111 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_233 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_234 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_235 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_236 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_237 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_238 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_239 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_240 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_241 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_242 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_243 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_244 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_245 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_246 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_247 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_248 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_249 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_250 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_251 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_252 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_253 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_254 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_255 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_256 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_257 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_258 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_259 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_260 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_261 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_262 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_263 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_264 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_265 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_266 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_267 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_268 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_269 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_270 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_271 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_272 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_273 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_274 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_275 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_276 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_277 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_112 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_113 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_114 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_115 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_278 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_279 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_280 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_281 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_282 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_283 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_284 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_285 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_286 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_287 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_288 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_289 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_290 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_291 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_292 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_293 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_294 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_295 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_296 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_297 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_298 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_299 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_300 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_301 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_302 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_303 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_304 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_305 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_306 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_307 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_308 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_309 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_310 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_311 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_312 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_313 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_116 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_117 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_118 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_119 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_120 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_121 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_122 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_123 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_124 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_125 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_126 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_127 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_128 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_129 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_130 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_131 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_132 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_133 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_134 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_135 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_136 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_137 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_138 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_139 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_140 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_141 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_142 (.VDD(vdd),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _081_ (.I(net44),
    .Z(_040_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _082_ (.I(_040_),
    .ZN(_041_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _083_ (.I(net9),
    .ZN(_042_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _084_ (.A1(net14),
    .A2(net13),
    .A3(net16),
    .A4(net15),
    .ZN(_043_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _085_ (.A1(net11),
    .A2(net10),
    .ZN(_044_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _086_ (.A1(_042_),
    .A2(net8),
    .A3(_043_),
    .A4(_044_),
    .ZN(_045_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _087_ (.A1(net25),
    .A2(net24),
    .ZN(_046_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _088_ (.A1(net22),
    .A2(net21),
    .A3(_046_),
    .ZN(_047_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _089_ (.A1(net18),
    .A2(net17),
    .A3(net20),
    .A4(net19),
    .Z(_048_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _090_ (.A1(_045_),
    .A2(_047_),
    .A3(_048_),
    .ZN(_049_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _091_ (.A1(net5),
    .A2(net4),
    .A3(net7),
    .A4(net6),
    .Z(_050_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _092_ (.I(net1),
    .ZN(_051_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _093_ (.A1(net32),
    .A2(net31),
    .A3(net3),
    .A4(net2),
    .ZN(_052_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _094_ (.A1(net30),
    .A2(net29),
    .ZN(_053_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _095_ (.A1(_051_),
    .A2(net12),
    .A3(_052_),
    .A4(_053_),
    .ZN(_054_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _096_ (.I(net26),
    .ZN(_055_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _097_ (.A1(_055_),
    .A2(net23),
    .A3(net27),
    .ZN(_056_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _098_ (.A1(net28),
    .A2(_050_),
    .A3(_054_),
    .A4(_056_),
    .ZN(_057_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _099_ (.A1(net41),
    .A2(_041_),
    .A3(_049_),
    .A4(_057_),
    .Z(_058_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _100_ (.I(_058_),
    .Z(_000_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _101_ (.I(net23),
    .ZN(_059_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _102_ (.A1(_059_),
    .A2(net27),
    .A3(net28),
    .ZN(_060_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _103_ (.A1(net33),
    .A2(net41),
    .A3(net42),
    .A4(_055_),
    .ZN(_061_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _104_ (.A1(_050_),
    .A2(_054_),
    .A3(_060_),
    .A4(_061_),
    .ZN(_062_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _105_ (.A1(_045_),
    .A2(_047_),
    .A3(_048_),
    .ZN(_063_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _106_ (.A1(_062_),
    .A2(_063_),
    .B(\d1.In_Data[0] ),
    .ZN(_064_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _107_ (.A1(_050_),
    .A2(_054_),
    .A3(_060_),
    .A4(_061_),
    .Z(_013_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _108_ (.A1(_045_),
    .A2(_047_),
    .A3(_048_),
    .Z(_014_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _109_ (.A1(net34),
    .A2(_013_),
    .A3(_014_),
    .ZN(_015_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _110_ (.A1(_040_),
    .A2(_064_),
    .A3(_015_),
    .ZN(_001_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _111_ (.A1(_062_),
    .A2(_063_),
    .B(\d1.In_Data[1] ),
    .ZN(_016_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _112_ (.A1(net35),
    .A2(_013_),
    .A3(_014_),
    .ZN(_017_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _113_ (.A1(_040_),
    .A2(_016_),
    .A3(_017_),
    .ZN(_002_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _114_ (.A1(_062_),
    .A2(_063_),
    .B(\d1.In_Data[2] ),
    .ZN(_018_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _115_ (.A1(net36),
    .A2(_013_),
    .A3(_014_),
    .ZN(_019_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _116_ (.A1(_040_),
    .A2(_018_),
    .A3(_019_),
    .ZN(_003_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _117_ (.A1(_062_),
    .A2(_063_),
    .B(\d1.In_Data[3] ),
    .ZN(_020_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _118_ (.A1(net37),
    .A2(_013_),
    .A3(_014_),
    .ZN(_021_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _119_ (.A1(_040_),
    .A2(_020_),
    .A3(_021_),
    .ZN(_004_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _120_ (.A1(_062_),
    .A2(_063_),
    .B(\d1.In_Data[4] ),
    .ZN(_022_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _121_ (.A1(net38),
    .A2(_013_),
    .A3(_014_),
    .ZN(_023_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _122_ (.A1(_040_),
    .A2(_022_),
    .A3(_023_),
    .ZN(_005_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _123_ (.A1(_062_),
    .A2(_063_),
    .B(\d1.In_Data[5] ),
    .ZN(_024_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _124_ (.A1(net39),
    .A2(_013_),
    .A3(_014_),
    .ZN(_025_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _125_ (.A1(_040_),
    .A2(_024_),
    .A3(_025_),
    .ZN(_006_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _126_ (.A1(_062_),
    .A2(_063_),
    .B(\d1.In_Data[6] ),
    .ZN(_026_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _127_ (.A1(net40),
    .A2(_013_),
    .A3(_014_),
    .ZN(_027_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _128_ (.A1(_040_),
    .A2(_026_),
    .A3(_027_),
    .ZN(_007_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _129_ (.A1(net33),
    .A2(net41),
    .ZN(_028_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _130_ (.A1(net42),
    .A2(_028_),
    .ZN(_029_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _131_ (.A1(\u5.Out_Data[0] ),
    .A2(_049_),
    .A3(_057_),
    .ZN(_030_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _132_ (.A1(o_wb_data[0]),
    .A2(_029_),
    .B(_041_),
    .ZN(_031_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _133_ (.A1(_029_),
    .A2(_030_),
    .B(_031_),
    .ZN(_008_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _134_ (.A1(\u5.Out_Data[1] ),
    .A2(_049_),
    .A3(_057_),
    .ZN(_032_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _135_ (.A1(o_wb_data[1]),
    .A2(_029_),
    .B(_041_),
    .ZN(_033_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _136_ (.A1(_029_),
    .A2(_032_),
    .B(_033_),
    .ZN(_009_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _137_ (.A1(\u5.Out_Data[2] ),
    .A2(_049_),
    .A3(_057_),
    .ZN(_034_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _138_ (.A1(o_wb_data[2]),
    .A2(_029_),
    .B(_041_),
    .ZN(_035_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _139_ (.A1(_029_),
    .A2(_034_),
    .B(_035_),
    .ZN(_010_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _140_ (.A1(\u5.Out_Data[3] ),
    .A2(_049_),
    .A3(_057_),
    .ZN(_036_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _141_ (.A1(o_wb_data[3]),
    .A2(_029_),
    .B(_041_),
    .ZN(_037_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _142_ (.A1(_029_),
    .A2(_036_),
    .B(_037_),
    .ZN(_011_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _143_ (.A1(\u5.Out_Data[4] ),
    .A2(_049_),
    .A3(_057_),
    .ZN(_038_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _144_ (.A1(o_wb_data[4]),
    .A2(_029_),
    .B(_041_),
    .ZN(_039_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _145_ (.A1(_029_),
    .A2(_038_),
    .B(_039_),
    .ZN(_012_),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _146_ (.D(_000_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(o_wb_ack),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _147_ (.D(\d3.Cout ),
    .RN(net44),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\u4.Data3[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _148_ (.D(\u4.Out_Data[0] ),
    .RN(net44),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\u5.Data3[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _149_ (.D(\u4.Out_Data[1] ),
    .RN(net44),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\u5.Data3[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _150_ (.D(\u4.Out_Data[2] ),
    .RN(net44),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\u5.Data3[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _151_ (.D(\u4.Out_Data[3] ),
    .RN(net44),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\u5.Data3[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _152_ (.D(\u4.Out_Data[4] ),
    .RN(net44),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\u5.Data3[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _153_ (.D(_001_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\d1.In_Data[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _154_ (.D(_002_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\d1.In_Data[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _155_ (.D(_003_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\d1.In_Data[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _156_ (.D(_004_),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\d1.In_Data[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _157_ (.D(_005_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\d1.In_Data[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _158_ (.D(_006_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\d1.In_Data[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _159_ (.D(_007_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\d1.In_Data[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _160_ (.D(_008_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(o_wb_data[0]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _161_ (.D(_009_),
    .CLK(clknet_2_0__leaf_clk),
    .Q(o_wb_data[1]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _162_ (.D(_010_),
    .CLK(clknet_2_2__leaf_clk),
    .Q(o_wb_data[2]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _163_ (.D(_011_),
    .CLK(clknet_2_2__leaf_clk),
    .Q(o_wb_data[3]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _164_ (.D(_012_),
    .CLK(clknet_2_2__leaf_clk),
    .Q(o_wb_data[4]),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_0__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_1__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_2__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_2__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_3__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_3__leaf_clk),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \d1._38_  (.A1(\d1.Out_Data[0] ),
    .A2(\d1.In_Data[0] ),
    .Z(\d1._00_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 \d1._39_  (.A1(\d1.Out_Data[1] ),
    .A2(\d1.In_Data[1] ),
    .A3(\d1._00_ ),
    .Z(\d1._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \d1._40_  (.I(\d1._01_ ),
    .Z(\d1.Sum[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \d1._41_  (.A1(\d1.Out_Data[0] ),
    .A2(\d1.In_Data[0] ),
    .ZN(\d1._02_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \d1._42_  (.A1(\d1.Out_Data[1] ),
    .A2(\d1.In_Data[1] ),
    .ZN(\d1._03_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \d1._43_  (.A1(\d1.Out_Data[1] ),
    .A2(\d1.In_Data[1] ),
    .ZN(\d1._04_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 \d1._44_  (.A1(\d1._02_ ),
    .A2(\d1._03_ ),
    .B(\d1._04_ ),
    .ZN(\d1._05_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \d1._45_  (.A1(\d1.Out_Data[2] ),
    .A2(\d1.In_Data[2] ),
    .Z(\d1._06_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \d1._46_  (.A1(\d1._05_ ),
    .A2(\d1._06_ ),
    .Z(\d1._07_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \d1._47_  (.I(\d1._07_ ),
    .Z(\d1.Sum[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \d1._48_  (.A1(\d1.Out_Data[2] ),
    .A2(\d1.In_Data[2] ),
    .ZN(\d1._08_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \d1._49_  (.A1(\d1._05_ ),
    .A2(\d1._06_ ),
    .ZN(\d1._09_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \d1._50_  (.A1(\d1._08_ ),
    .A2(\d1._09_ ),
    .ZN(\d1._10_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \d1._51_  (.A1(\d1.Out_Data[3] ),
    .A2(\d1.In_Data[3] ),
    .Z(\d1._11_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \d1._52_  (.A1(\d1._10_ ),
    .A2(\d1._11_ ),
    .Z(\d1._12_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \d1._53_  (.I(\d1._12_ ),
    .Z(\d1.Sum[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \d1._54_  (.A1(\d1._06_ ),
    .A2(\d1._11_ ),
    .Z(\d1._13_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \d1._55_  (.A1(\d1.Out_Data[3] ),
    .A2(\d1.In_Data[3] ),
    .ZN(\d1._14_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 \d1._56_  (.A1(\d1.Out_Data[3] ),
    .A2(\d1.In_Data[3] ),
    .B(\d1.Out_Data[2] ),
    .C(\d1.In_Data[2] ),
    .ZN(\d1._15_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \d1._57_  (.A1(\d1._14_ ),
    .A2(\d1._15_ ),
    .ZN(\d1._16_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 \d1._58_  (.A1(\d1._05_ ),
    .A2(\d1._13_ ),
    .B(\d1._16_ ),
    .ZN(\d1._17_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 \d1._59_  (.A1(\d1.Out_Data[4] ),
    .A2(\d1.In_Data[4] ),
    .ZN(\d1._18_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \d1._60_  (.A1(\d1._17_ ),
    .A2(\d1._18_ ),
    .Z(\d1._19_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \d1._61_  (.I(\d1._19_ ),
    .Z(\d1.Sum[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \d1._62_  (.A1(\d1.Out_Data[4] ),
    .A2(\d1.In_Data[4] ),
    .ZN(\d1._20_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 \d1._63_  (.A1(\d1._17_ ),
    .A2(\d1._18_ ),
    .B(\d1._20_ ),
    .ZN(\d1._21_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \d1._64_  (.A1(\d1.Out_Data[5] ),
    .A2(\d1.In_Data[5] ),
    .Z(\d1._22_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \d1._65_  (.A1(\d1._21_ ),
    .A2(\d1._22_ ),
    .Z(\d1._23_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \d1._66_  (.I(\d1._23_ ),
    .Z(\d1.Sum[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \d1._67_  (.A1(\d1.Out_Data[1] ),
    .A2(\d1.In_Data[1] ),
    .Z(\d1._24_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \d1._68_  (.A1(\d1.Out_Data[1] ),
    .A2(\d1.In_Data[1] ),
    .Z(\d1._25_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 \d1._69_  (.A1(\d1._00_ ),
    .A2(\d1._24_ ),
    .B(\d1._25_ ),
    .ZN(\d1._26_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \d1._70_  (.A1(\d1._06_ ),
    .A2(\d1._11_ ),
    .ZN(\d1._27_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 \d1._71_  (.A1(\d1._26_ ),
    .A2(\d1._27_ ),
    .B(\d1._15_ ),
    .C(\d1._14_ ),
    .ZN(\d1._28_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \d1._72_  (.I(\d1._22_ ),
    .ZN(\d1._29_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \d1._73_  (.A1(\d1._18_ ),
    .A2(\d1._29_ ),
    .ZN(\d1._30_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \d1._74_  (.A1(\d1.Out_Data[5] ),
    .A2(\d1.In_Data[5] ),
    .ZN(\d1._31_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \d1._75_  (.A1(\d1._20_ ),
    .A2(\d1._31_ ),
    .ZN(\d1._32_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 \d1._76_  (.A1(\d1.Out_Data[5] ),
    .A2(\d1.In_Data[5] ),
    .B1(\d1._28_ ),
    .B2(\d1._30_ ),
    .C(\d1._32_ ),
    .ZN(\d1._33_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 \d1._77_  (.A1(\d1.Out_Data[6] ),
    .A2(\d1.In_Data[6] ),
    .A3(\d1._33_ ),
    .ZN(\d1._34_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \d1._78_  (.I(\d1._34_ ),
    .Z(\d1.Sum[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \d1._79_  (.A1(\d1.Out_Data[0] ),
    .A2(\d1.In_Data[0] ),
    .Z(\d1._35_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \d1._80_  (.I(\d1._35_ ),
    .Z(\d1.Sum[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \d1._81_  (.A1(\d1.Out_Data[6] ),
    .A2(\d1.In_Data[6] ),
    .ZN(\d1._36_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \d1._82_  (.A1(\d1.Out_Data[6] ),
    .A2(\d1.In_Data[6] ),
    .ZN(\d1._37_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 \d1._83_  (.A1(\d1._33_ ),
    .A2(\d1._36_ ),
    .B(\d1._37_ ),
    .ZN(\d1.Cout ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 \d1._84_  (.D(\d1.Sum[0] ),
    .RN(net44),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\d1.Out_Data[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \d1._85_  (.D(\d1.Sum[1] ),
    .RN(net44),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\d1.Out_Data[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \d1._86_  (.D(\d1.Sum[2] ),
    .RN(net44),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\d1.Out_Data[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \d1._87_  (.D(\d1.Sum[3] ),
    .RN(net44),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\d1.Out_Data[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 \d1._88_  (.D(\d1.Sum[4] ),
    .RN(net44),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\d1.Out_Data[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \d1._89_  (.D(\d1.Sum[5] ),
    .RN(net44),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\d1.Out_Data[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 \d1._90_  (.D(\d1.Sum[6] ),
    .RN(net44),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\d1.Out_Data[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \d2._38_  (.A1(\d2.Out_Data[0] ),
    .A2(\d1.Out_Data[0] ),
    .Z(\d2._00_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 \d2._39_  (.A1(\d2.Out_Data[1] ),
    .A2(\d1.Out_Data[1] ),
    .A3(\d2._00_ ),
    .Z(\d2._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \d2._40_  (.I(\d2._01_ ),
    .Z(\d2.Sum[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \d2._41_  (.A1(\d2.Out_Data[0] ),
    .A2(\d1.Out_Data[0] ),
    .ZN(\d2._02_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \d2._42_  (.A1(\d2.Out_Data[1] ),
    .A2(\d1.Out_Data[1] ),
    .ZN(\d2._03_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \d2._43_  (.A1(\d2.Out_Data[1] ),
    .A2(\d1.Out_Data[1] ),
    .ZN(\d2._04_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 \d2._44_  (.A1(\d2._02_ ),
    .A2(\d2._03_ ),
    .B(\d2._04_ ),
    .ZN(\d2._05_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \d2._45_  (.A1(\d2.Out_Data[2] ),
    .A2(\d1.Out_Data[2] ),
    .Z(\d2._06_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \d2._46_  (.A1(\d2._05_ ),
    .A2(\d2._06_ ),
    .Z(\d2._07_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \d2._47_  (.I(\d2._07_ ),
    .Z(\d2.Sum[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \d2._48_  (.A1(\d2.Out_Data[2] ),
    .A2(\d1.Out_Data[2] ),
    .ZN(\d2._08_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \d2._49_  (.A1(\d2._05_ ),
    .A2(\d2._06_ ),
    .ZN(\d2._09_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \d2._50_  (.A1(\d2._08_ ),
    .A2(\d2._09_ ),
    .ZN(\d2._10_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \d2._51_  (.A1(\d2.Out_Data[3] ),
    .A2(\d1.Out_Data[3] ),
    .Z(\d2._11_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \d2._52_  (.A1(\d2._10_ ),
    .A2(\d2._11_ ),
    .Z(\d2._12_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \d2._53_  (.I(\d2._12_ ),
    .Z(\d2.Sum[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \d2._54_  (.A1(\d2._06_ ),
    .A2(\d2._11_ ),
    .Z(\d2._13_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 \d2._55_  (.A1(\d2.Out_Data[3] ),
    .A2(\d1.Out_Data[3] ),
    .ZN(\d2._14_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 \d2._56_  (.A1(\d2.Out_Data[3] ),
    .A2(\d1.Out_Data[3] ),
    .B(\d2.Out_Data[2] ),
    .C(\d1.Out_Data[2] ),
    .ZN(\d2._15_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \d2._57_  (.A1(\d2._14_ ),
    .A2(\d2._15_ ),
    .ZN(\d2._16_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 \d2._58_  (.A1(\d2._05_ ),
    .A2(\d2._13_ ),
    .B(\d2._16_ ),
    .ZN(\d2._17_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 \d2._59_  (.A1(\d2.Out_Data[4] ),
    .A2(\d1.Out_Data[4] ),
    .ZN(\d2._18_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \d2._60_  (.A1(\d2._17_ ),
    .A2(\d2._18_ ),
    .Z(\d2._19_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \d2._61_  (.I(\d2._19_ ),
    .Z(\d2.Sum[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \d2._62_  (.A1(\d2.Out_Data[4] ),
    .A2(\d1.Out_Data[4] ),
    .ZN(\d2._20_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 \d2._63_  (.A1(\d2._17_ ),
    .A2(\d2._18_ ),
    .B(\d2._20_ ),
    .ZN(\d2._21_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \d2._64_  (.A1(\d2.Out_Data[5] ),
    .A2(\d1.Out_Data[5] ),
    .Z(\d2._22_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \d2._65_  (.A1(\d2._21_ ),
    .A2(\d2._22_ ),
    .Z(\d2._23_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \d2._66_  (.I(\d2._23_ ),
    .Z(\d2.Sum[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \d2._67_  (.A1(\d2.Out_Data[1] ),
    .A2(\d1.Out_Data[1] ),
    .Z(\d2._24_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \d2._68_  (.A1(\d2.Out_Data[1] ),
    .A2(\d1.Out_Data[1] ),
    .Z(\d2._25_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 \d2._69_  (.A1(\d2._00_ ),
    .A2(\d2._24_ ),
    .B(\d2._25_ ),
    .ZN(\d2._26_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \d2._70_  (.A1(\d2._06_ ),
    .A2(\d2._11_ ),
    .ZN(\d2._27_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 \d2._71_  (.A1(\d2._26_ ),
    .A2(\d2._27_ ),
    .B(\d2._15_ ),
    .C(\d2._14_ ),
    .ZN(\d2._28_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \d2._72_  (.I(\d2._22_ ),
    .ZN(\d2._29_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \d2._73_  (.A1(\d2._18_ ),
    .A2(\d2._29_ ),
    .ZN(\d2._30_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \d2._74_  (.A1(\d2.Out_Data[5] ),
    .A2(\d1.Out_Data[5] ),
    .ZN(\d2._31_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \d2._75_  (.A1(\d2._20_ ),
    .A2(\d2._31_ ),
    .ZN(\d2._32_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 \d2._76_  (.A1(\d2.Out_Data[5] ),
    .A2(\d1.Out_Data[5] ),
    .B1(\d2._28_ ),
    .B2(\d2._30_ ),
    .C(\d2._32_ ),
    .ZN(\d2._33_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 \d2._77_  (.A1(\d2.Out_Data[6] ),
    .A2(\d1.Out_Data[6] ),
    .A3(\d2._33_ ),
    .ZN(\d2._34_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \d2._78_  (.I(\d2._34_ ),
    .Z(\d2.Sum[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \d2._79_  (.A1(\d2.Out_Data[0] ),
    .A2(\d1.Out_Data[0] ),
    .Z(\d2._35_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \d2._80_  (.I(\d2._35_ ),
    .Z(\d2.Sum[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \d2._81_  (.A1(\d2.Out_Data[6] ),
    .A2(\d1.Out_Data[6] ),
    .ZN(\d2._36_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \d2._82_  (.A1(\d2.Out_Data[6] ),
    .A2(\d1.Out_Data[6] ),
    .ZN(\d2._37_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 \d2._83_  (.A1(\d2._33_ ),
    .A2(\d2._36_ ),
    .B(\d2._37_ ),
    .ZN(\d2.Cout ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 \d2._84_  (.D(\d2.Sum[0] ),
    .RN(net44),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\d2.Out_Data[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \d2._85_  (.D(\d2.Sum[1] ),
    .RN(net44),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\d2.Out_Data[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \d2._86_  (.D(\d2.Sum[2] ),
    .RN(net43),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\d2.Out_Data[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_4 \d2._87_  (.D(\d2.Sum[3] ),
    .RN(net43),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\d2.Out_Data[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 \d2._88_  (.D(\d2.Sum[4] ),
    .RN(net43),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\d2.Out_Data[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 \d2._89_  (.D(\d2.Sum[5] ),
    .RN(net44),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\d2.Out_Data[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 \d2._90_  (.D(\d2.Sum[6] ),
    .RN(net44),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\d2.Out_Data[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \d3._38_  (.A1(\d3.Out_Data[0] ),
    .A2(\d2.Out_Data[0] ),
    .Z(\d3._00_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 \d3._39_  (.A1(\d3.Out_Data[1] ),
    .A2(\d2.Out_Data[1] ),
    .A3(\d3._00_ ),
    .Z(\d3._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \d3._40_  (.I(\d3._01_ ),
    .Z(\d3.Sum[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \d3._41_  (.A1(\d3.Out_Data[0] ),
    .A2(\d2.Out_Data[0] ),
    .ZN(\d3._02_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \d3._42_  (.A1(\d3.Out_Data[1] ),
    .A2(\d2.Out_Data[1] ),
    .ZN(\d3._03_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \d3._43_  (.A1(\d3.Out_Data[1] ),
    .A2(\d2.Out_Data[1] ),
    .ZN(\d3._04_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 \d3._44_  (.A1(\d3._02_ ),
    .A2(\d3._03_ ),
    .B(\d3._04_ ),
    .ZN(\d3._05_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \d3._45_  (.A1(\d3.Out_Data[2] ),
    .A2(\d2.Out_Data[2] ),
    .Z(\d3._06_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \d3._46_  (.A1(\d3._05_ ),
    .A2(\d3._06_ ),
    .Z(\d3._07_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \d3._47_  (.I(\d3._07_ ),
    .Z(\d3.Sum[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \d3._48_  (.A1(\d3.Out_Data[2] ),
    .A2(\d2.Out_Data[2] ),
    .ZN(\d3._08_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \d3._49_  (.A1(\d3._05_ ),
    .A2(\d3._06_ ),
    .ZN(\d3._09_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \d3._50_  (.A1(\d3._08_ ),
    .A2(\d3._09_ ),
    .ZN(\d3._10_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \d3._51_  (.A1(\d3.Out_Data[3] ),
    .A2(\d2.Out_Data[3] ),
    .Z(\d3._11_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \d3._52_  (.A1(\d3._10_ ),
    .A2(\d3._11_ ),
    .Z(\d3._12_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \d3._53_  (.I(\d3._12_ ),
    .Z(\d3.Sum[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \d3._54_  (.A1(\d3._06_ ),
    .A2(\d3._11_ ),
    .Z(\d3._13_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 \d3._55_  (.A1(\d3.Out_Data[3] ),
    .A2(\d2.Out_Data[3] ),
    .ZN(\d3._14_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 \d3._56_  (.A1(\d3.Out_Data[3] ),
    .A2(\d2.Out_Data[3] ),
    .B(\d3.Out_Data[2] ),
    .C(\d2.Out_Data[2] ),
    .ZN(\d3._15_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \d3._57_  (.A1(\d3._14_ ),
    .A2(\d3._15_ ),
    .ZN(\d3._16_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 \d3._58_  (.A1(\d3._05_ ),
    .A2(\d3._13_ ),
    .B(\d3._16_ ),
    .ZN(\d3._17_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 \d3._59_  (.A1(\d3.Out_Data[4] ),
    .A2(\d2.Out_Data[4] ),
    .ZN(\d3._18_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \d3._60_  (.A1(\d3._17_ ),
    .A2(\d3._18_ ),
    .Z(\d3._19_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \d3._61_  (.I(\d3._19_ ),
    .Z(\d3.Sum[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \d3._62_  (.A1(\d3.Out_Data[4] ),
    .A2(\d2.Out_Data[4] ),
    .ZN(\d3._20_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 \d3._63_  (.A1(\d3._17_ ),
    .A2(\d3._18_ ),
    .B(\d3._20_ ),
    .ZN(\d3._21_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \d3._64_  (.A1(\d3.Out_Data[5] ),
    .A2(\d2.Out_Data[5] ),
    .Z(\d3._22_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \d3._65_  (.A1(\d3._21_ ),
    .A2(\d3._22_ ),
    .Z(\d3._23_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \d3._66_  (.I(\d3._23_ ),
    .Z(\d3.Sum[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 \d3._67_  (.A1(\d3.Out_Data[1] ),
    .A2(\d2.Out_Data[1] ),
    .Z(\d3._24_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 \d3._68_  (.A1(\d3.Out_Data[1] ),
    .A2(\d2.Out_Data[1] ),
    .Z(\d3._25_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 \d3._69_  (.A1(\d3._00_ ),
    .A2(\d3._24_ ),
    .B(\d3._25_ ),
    .ZN(\d3._26_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \d3._70_  (.A1(\d3._06_ ),
    .A2(\d3._11_ ),
    .ZN(\d3._27_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 \d3._71_  (.A1(\d3._26_ ),
    .A2(\d3._27_ ),
    .B(\d3._15_ ),
    .C(\d3._14_ ),
    .ZN(\d3._28_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \d3._72_  (.I(\d3._22_ ),
    .ZN(\d3._29_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \d3._73_  (.A1(\d3._18_ ),
    .A2(\d3._29_ ),
    .ZN(\d3._30_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \d3._74_  (.A1(\d3.Out_Data[5] ),
    .A2(\d2.Out_Data[5] ),
    .ZN(\d3._31_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \d3._75_  (.A1(\d3._20_ ),
    .A2(\d3._31_ ),
    .ZN(\d3._32_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 \d3._76_  (.A1(\d3.Out_Data[5] ),
    .A2(\d2.Out_Data[5] ),
    .B1(\d3._28_ ),
    .B2(\d3._30_ ),
    .C(\d3._32_ ),
    .ZN(\d3._33_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 \d3._77_  (.A1(\d3.Out_Data[6] ),
    .A2(\d2.Out_Data[6] ),
    .A3(\d3._33_ ),
    .ZN(\d3._34_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \d3._78_  (.I(\d3._34_ ),
    .Z(\d3.Sum[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \d3._79_  (.A1(\d3.Out_Data[0] ),
    .A2(\d2.Out_Data[0] ),
    .Z(\d3._35_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \d3._80_  (.I(\d3._35_ ),
    .Z(\d3.Sum[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \d3._81_  (.A1(\d3.Out_Data[6] ),
    .A2(\d2.Out_Data[6] ),
    .ZN(\d3._36_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \d3._82_  (.A1(\d3.Out_Data[6] ),
    .A2(\d2.Out_Data[6] ),
    .ZN(\d3._37_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 \d3._83_  (.A1(\d3._33_ ),
    .A2(\d3._36_ ),
    .B(\d3._37_ ),
    .ZN(\d3.Cout ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 \d3._84_  (.D(\d3.Sum[0] ),
    .RN(net43),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\d3.Out_Data[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 \d3._85_  (.D(\d3.Sum[1] ),
    .RN(net43),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\d3.Out_Data[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 \d3._86_  (.D(\d3.Sum[2] ),
    .RN(net43),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\d3.Out_Data[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 \d3._87_  (.D(\d3.Sum[3] ),
    .RN(net43),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\d3.Out_Data[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 \d3._88_  (.D(\d3.Sum[4] ),
    .RN(net43),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\d3.Out_Data[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 \d3._89_  (.D(\d3.Sum[5] ),
    .RN(net44),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\d3.Out_Data[5] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 \d3._90_  (.D(\d3.Sum[6] ),
    .RN(net44),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\d3.Out_Data[6] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 fanout44 (.I(net43),
    .Z(net44),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1 (.I(i_wb_addr[0]),
    .Z(net1),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input10 (.I(i_wb_addr[18]),
    .Z(net10),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input11 (.I(i_wb_addr[19]),
    .Z(net11),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input12 (.I(i_wb_addr[1]),
    .Z(net12),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input13 (.I(i_wb_addr[20]),
    .Z(net13),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input14 (.I(i_wb_addr[21]),
    .Z(net14),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input15 (.I(i_wb_addr[22]),
    .Z(net15),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input16 (.I(i_wb_addr[23]),
    .Z(net16),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input17 (.I(i_wb_addr[24]),
    .Z(net17),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input18 (.I(i_wb_addr[25]),
    .Z(net18),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input19 (.I(i_wb_addr[26]),
    .Z(net19),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input2 (.I(i_wb_addr[10]),
    .Z(net2),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input20 (.I(i_wb_addr[27]),
    .Z(net20),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input21 (.I(i_wb_addr[28]),
    .Z(net21),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input22 (.I(i_wb_addr[29]),
    .Z(net22),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input23 (.I(i_wb_addr[2]),
    .Z(net23),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input24 (.I(i_wb_addr[30]),
    .Z(net24),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input25 (.I(i_wb_addr[31]),
    .Z(net25),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input26 (.I(i_wb_addr[3]),
    .Z(net26),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input27 (.I(i_wb_addr[4]),
    .Z(net27),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input28 (.I(i_wb_addr[5]),
    .Z(net28),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input29 (.I(i_wb_addr[6]),
    .Z(net29),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(i_wb_addr[11]),
    .Z(net3),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input30 (.I(i_wb_addr[7]),
    .Z(net30),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input31 (.I(i_wb_addr[8]),
    .Z(net31),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input32 (.I(i_wb_addr[9]),
    .Z(net32),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input33 (.I(i_wb_cyc),
    .Z(net33),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input34 (.I(i_wb_data[0]),
    .Z(net34),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input35 (.I(i_wb_data[1]),
    .Z(net35),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input36 (.I(i_wb_data[2]),
    .Z(net36),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input37 (.I(i_wb_data[3]),
    .Z(net37),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input38 (.I(i_wb_data[4]),
    .Z(net38),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input39 (.I(i_wb_data[5]),
    .Z(net39),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input4 (.I(i_wb_addr[12]),
    .Z(net4),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input40 (.I(i_wb_data[6]),
    .Z(net40),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input41 (.I(i_wb_stb),
    .Z(net41),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input42 (.I(i_wb_we),
    .Z(net42),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input43 (.I(reset),
    .Z(net43),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(i_wb_addr[13]),
    .Z(net5),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input6 (.I(i_wb_addr[14]),
    .Z(net6),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(i_wb_addr[15]),
    .Z(net7),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(i_wb_addr[16]),
    .Z(net8),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input9 (.I(i_wb_addr[17]),
    .Z(net9),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \u4._33_  (.I(\u4.Data3[0] ),
    .ZN(\u4._00_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \u4._34_  (.A1(\u4._00_ ),
    .A2(\d2.Cout ),
    .ZN(\u4._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \u4._35_  (.A1(\u4.Data3[0] ),
    .A2(\d2.Cout ),
    .Z(\u4._02_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \u4._36_  (.A1(\d3.Cout ),
    .A2(\u4._02_ ),
    .ZN(\u4._03_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 \u4._37_  (.A1(net65),
    .A2(net55),
    .A3(net45),
    .ZN(\u4._04_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u4._37__45  (.ZN(net45),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u4._37__55  (.ZN(net55),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u4._37__65  (.ZN(net65),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 \u4._38_  (.A1(\u4._01_ ),
    .A2(\u4._03_ ),
    .A3(\u4._04_ ),
    .Z(\u4._05_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 \u4._39_  (.I(\u4._05_ ),
    .Z(\u4.Out_Data[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 \u4._40_  (.A1(\u4._00_ ),
    .A2(\d2.Cout ),
    .A3(\u4._04_ ),
    .ZN(\u4._06_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 \u4._41_  (.A1(\u4._00_ ),
    .A2(\d2.Cout ),
    .B(\u4._04_ ),
    .ZN(\u4._07_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 \u4._42_  (.A1(\u4._03_ ),
    .A2(\u4._06_ ),
    .B(\u4._07_ ),
    .ZN(\u4._08_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 \u4._43_  (.A1(net67),
    .A2(net58),
    .A3(net48),
    .ZN(\u4._09_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u4._43__48  (.ZN(net48),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u4._43__58  (.ZN(net58),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u4._43__67  (.ZN(net67),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \u4._44_  (.A1(net56),
    .A2(net46),
    .ZN(\u4._10_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u4._44__46  (.ZN(net46),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u4._44__56  (.ZN(net56),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \u4._45_  (.A1(net57),
    .A2(net47),
    .ZN(\u4._11_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u4._45__47  (.ZN(net47),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u4._45__57  (.ZN(net57),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 \u4._46_  (.A1(net66),
    .A2(\u4._10_ ),
    .B(\u4._11_ ),
    .ZN(\u4._12_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u4._46__66  (.ZN(net66),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \u4._47_  (.A1(\u4._09_ ),
    .A2(\u4._12_ ),
    .Z(\u4._13_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \u4._48_  (.A1(\u4._08_ ),
    .A2(\u4._13_ ),
    .Z(\u4._14_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 \u4._49_  (.I(\u4._14_ ),
    .Z(\u4.Out_Data[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 \u4._50_  (.A1(net69),
    .A2(net61),
    .A3(net51),
    .Z(\u4._15_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u4._50__51  (.ZN(net51),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u4._50__61  (.ZN(net61),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u4._50__69  (.ZN(net69),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \u4._51_  (.I(\u4._15_ ),
    .ZN(\u4._16_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \u4._52_  (.A1(net59),
    .A2(net49),
    .ZN(\u4._17_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u4._52__49  (.ZN(net49),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u4._52__59  (.ZN(net59),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \u4._53_  (.A1(net60),
    .A2(net50),
    .ZN(\u4._18_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u4._53__50  (.ZN(net50),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u4._53__60  (.ZN(net60),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 \u4._54_  (.A1(net68),
    .A2(\u4._17_ ),
    .B(\u4._18_ ),
    .ZN(\u4._19_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u4._54__68  (.ZN(net68),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \u4._55_  (.A1(\u4._09_ ),
    .A2(\u4._12_ ),
    .ZN(\u4._20_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \u4._56_  (.A1(\u4._08_ ),
    .A2(\u4._13_ ),
    .ZN(\u4._21_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \u4._57_  (.A1(\u4._20_ ),
    .A2(\u4._21_ ),
    .ZN(\u4._22_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 \u4._58_  (.A1(\u4._16_ ),
    .A2(\u4._19_ ),
    .A3(\u4._22_ ),
    .Z(\u4._23_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 \u4._59_  (.I(\u4._23_ ),
    .Z(\u4.Out_Data[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \u4._60_  (.A1(net62),
    .A2(net52),
    .ZN(\u4._24_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u4._60__52  (.ZN(net52),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u4._60__62  (.ZN(net62),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \u4._61_  (.A1(net63),
    .A2(net53),
    .ZN(\u4._25_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u4._61__53  (.ZN(net53),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u4._61__63  (.ZN(net63),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 \u4._62_  (.A1(net70),
    .A2(\u4._24_ ),
    .B(\u4._25_ ),
    .ZN(\u4._26_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u4._62__70  (.ZN(net70),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 \u4._63_  (.A1(net64),
    .A2(net54),
    .A3(net71),
    .ZN(\u4._27_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u4._63__54  (.ZN(net54),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u4._63__64  (.ZN(net64),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u4._63__71  (.ZN(net71),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 \u4._64_  (.A1(\u4._09_ ),
    .A2(\u4._12_ ),
    .B1(\u4._16_ ),
    .B2(\u4._19_ ),
    .ZN(\u4._28_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \u4._65_  (.A1(\u4._16_ ),
    .A2(\u4._19_ ),
    .ZN(\u4._29_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \u4._66_  (.A1(\u4._21_ ),
    .A2(\u4._28_ ),
    .B(\u4._29_ ),
    .ZN(\u4._30_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 \u4._67_  (.A1(\u4._26_ ),
    .A2(\u4._27_ ),
    .A3(\u4._30_ ),
    .Z(\u4._31_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \u4._68_  (.I(\u4._31_ ),
    .Z(\u4.Out_Data[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \u4._69_  (.A1(\d3.Cout ),
    .A2(\u4._02_ ),
    .Z(\u4._32_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \u4._70_  (.I(\u4._32_ ),
    .Z(\u4.Out_Data[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \u5._33_  (.I(\u5.Data3[0] ),
    .ZN(\u5._00_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \u5._34_  (.A1(\u5._00_ ),
    .A2(\d1.Cout ),
    .ZN(\u5._01_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \u5._35_  (.A1(\u5.Data3[0] ),
    .A2(\d1.Cout ),
    .Z(\u5._02_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \u5._36_  (.A1(\u4.Out_Data[0] ),
    .A2(\u5._02_ ),
    .ZN(\u5._03_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 \u5._37_  (.A1(\u5.Data3[1] ),
    .A2(\u4.Out_Data[1] ),
    .A3(net72),
    .ZN(\u5._04_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u5._37__72  (.ZN(net72),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 \u5._38_  (.A1(\u5._01_ ),
    .A2(\u5._03_ ),
    .A3(\u5._04_ ),
    .Z(\u5._05_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \u5._39_  (.I(\u5._05_ ),
    .Z(\u5.Out_Data[1] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 \u5._40_  (.A1(\u5._00_ ),
    .A2(\d1.Cout ),
    .A3(\u5._04_ ),
    .ZN(\u5._06_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 \u5._41_  (.A1(\u5._00_ ),
    .A2(\d1.Cout ),
    .B(\u5._04_ ),
    .ZN(\u5._07_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 \u5._42_  (.A1(\u5._03_ ),
    .A2(\u5._06_ ),
    .B(\u5._07_ ),
    .ZN(\u5._08_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 \u5._43_  (.A1(\u5.Data3[2] ),
    .A2(\u4.Out_Data[2] ),
    .A3(net75),
    .ZN(\u5._09_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u5._43__75  (.ZN(net75),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \u5._44_  (.A1(\u4.Out_Data[1] ),
    .A2(net73),
    .ZN(\u5._10_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u5._44__73  (.ZN(net73),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \u5._45_  (.A1(\u4.Out_Data[1] ),
    .A2(net74),
    .ZN(\u5._11_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u5._45__74  (.ZN(net74),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 \u5._46_  (.A1(\u5.Data3[1] ),
    .A2(\u5._10_ ),
    .B(\u5._11_ ),
    .ZN(\u5._12_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \u5._47_  (.A1(\u5._09_ ),
    .A2(\u5._12_ ),
    .Z(\u5._13_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \u5._48_  (.A1(\u5._08_ ),
    .A2(\u5._13_ ),
    .Z(\u5._14_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \u5._49_  (.I(\u5._14_ ),
    .Z(\u5.Out_Data[2] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 \u5._50_  (.A1(\u5.Data3[3] ),
    .A2(\u4.Out_Data[3] ),
    .A3(net78),
    .Z(\u5._15_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u5._50__78  (.ZN(net78),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 \u5._51_  (.I(\u5._15_ ),
    .ZN(\u5._16_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \u5._52_  (.A1(\u4.Out_Data[2] ),
    .A2(net76),
    .ZN(\u5._17_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u5._52__76  (.ZN(net76),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \u5._53_  (.A1(\u4.Out_Data[2] ),
    .A2(net77),
    .ZN(\u5._18_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u5._53__77  (.ZN(net77),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 \u5._54_  (.A1(\u5.Data3[2] ),
    .A2(\u5._17_ ),
    .B(\u5._18_ ),
    .ZN(\u5._19_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \u5._55_  (.A1(\u5._09_ ),
    .A2(\u5._12_ ),
    .ZN(\u5._20_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \u5._56_  (.A1(\u5._08_ ),
    .A2(\u5._13_ ),
    .ZN(\u5._21_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \u5._57_  (.A1(\u5._20_ ),
    .A2(\u5._21_ ),
    .ZN(\u5._22_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 \u5._58_  (.A1(\u5._16_ ),
    .A2(\u5._19_ ),
    .A3(\u5._22_ ),
    .Z(\u5._23_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \u5._59_  (.I(\u5._23_ ),
    .Z(\u5.Out_Data[3] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \u5._60_  (.A1(\u4.Out_Data[3] ),
    .A2(net79),
    .ZN(\u5._24_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u5._60__79  (.ZN(net79),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 \u5._61_  (.A1(\u4.Out_Data[3] ),
    .A2(net80),
    .ZN(\u5._25_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u5._61__80  (.ZN(net80),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 \u5._62_  (.A1(\u5.Data3[3] ),
    .A2(\u5._24_ ),
    .B(\u5._25_ ),
    .ZN(\u5._26_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 \u5._63_  (.A1(\u4.Out_Data[4] ),
    .A2(net81),
    .A3(\u5.Data3[4] ),
    .ZN(\u5._27_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__tiel \u5._63__81  (.ZN(net81),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 \u5._64_  (.A1(\u5._09_ ),
    .A2(\u5._12_ ),
    .B1(\u5._16_ ),
    .B2(\u5._19_ ),
    .ZN(\u5._28_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 \u5._65_  (.A1(\u5._16_ ),
    .A2(\u5._19_ ),
    .ZN(\u5._29_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 \u5._66_  (.A1(\u5._21_ ),
    .A2(\u5._28_ ),
    .B(\u5._29_ ),
    .ZN(\u5._30_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 \u5._67_  (.A1(\u5._26_ ),
    .A2(\u5._27_ ),
    .A3(\u5._30_ ),
    .Z(\u5._31_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \u5._68_  (.I(\u5._31_ ),
    .Z(\u5.Out_Data[4] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 \u5._69_  (.A1(\u4.Out_Data[0] ),
    .A2(\u5._02_ ),
    .Z(\u5._32_ ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 \u5._70_  (.I(\u5._32_ ),
    .Z(\u5.Out_Data[0] ),
    .VDD(vdd),
    .VNW(vdd),
    .VPW(vss),
    .VSS(vss));
 assign o_wb_stall = net82;
endmodule
