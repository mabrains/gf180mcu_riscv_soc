module user_project_wrapper (user_clock2,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    vss,
    vdd,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    user_irq,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input user_clock2;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input vss;
 input vdd;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [63:0] la_data_in;
 output [63:0] la_data_out;
 input [63:0] la_oenb;
 output [2:0] user_irq;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire i2c_rst_n;
 wire i2cm_clk_i;
 wire i2cm_clk_o;
 wire i2cm_clk_oen;
 wire i2cm_data_i;
 wire i2cm_data_o;
 wire i2cm_data_oen;
 wire i2cm_intr_o;
 wire pulse1m_mclk;
 wire reg_peri_ack;
 wire \reg_peri_addr[0] ;
 wire \reg_peri_addr[10] ;
 wire \reg_peri_addr[1] ;
 wire \reg_peri_addr[2] ;
 wire \reg_peri_addr[3] ;
 wire \reg_peri_addr[4] ;
 wire \reg_peri_addr[5] ;
 wire \reg_peri_addr[6] ;
 wire \reg_peri_addr[7] ;
 wire \reg_peri_addr[8] ;
 wire \reg_peri_addr[9] ;
 wire \reg_peri_be[0] ;
 wire \reg_peri_be[1] ;
 wire \reg_peri_be[2] ;
 wire \reg_peri_be[3] ;
 wire reg_peri_cs;
 wire \reg_peri_rdata[0] ;
 wire \reg_peri_rdata[10] ;
 wire \reg_peri_rdata[11] ;
 wire \reg_peri_rdata[12] ;
 wire \reg_peri_rdata[13] ;
 wire \reg_peri_rdata[14] ;
 wire \reg_peri_rdata[15] ;
 wire \reg_peri_rdata[16] ;
 wire \reg_peri_rdata[17] ;
 wire \reg_peri_rdata[18] ;
 wire \reg_peri_rdata[19] ;
 wire \reg_peri_rdata[1] ;
 wire \reg_peri_rdata[20] ;
 wire \reg_peri_rdata[21] ;
 wire \reg_peri_rdata[22] ;
 wire \reg_peri_rdata[23] ;
 wire \reg_peri_rdata[24] ;
 wire \reg_peri_rdata[25] ;
 wire \reg_peri_rdata[26] ;
 wire \reg_peri_rdata[27] ;
 wire \reg_peri_rdata[28] ;
 wire \reg_peri_rdata[29] ;
 wire \reg_peri_rdata[2] ;
 wire \reg_peri_rdata[30] ;
 wire \reg_peri_rdata[31] ;
 wire \reg_peri_rdata[3] ;
 wire \reg_peri_rdata[4] ;
 wire \reg_peri_rdata[5] ;
 wire \reg_peri_rdata[6] ;
 wire \reg_peri_rdata[7] ;
 wire \reg_peri_rdata[8] ;
 wire \reg_peri_rdata[9] ;
 wire \reg_peri_wdata[0] ;
 wire \reg_peri_wdata[10] ;
 wire \reg_peri_wdata[11] ;
 wire \reg_peri_wdata[12] ;
 wire \reg_peri_wdata[13] ;
 wire \reg_peri_wdata[14] ;
 wire \reg_peri_wdata[15] ;
 wire \reg_peri_wdata[16] ;
 wire \reg_peri_wdata[17] ;
 wire \reg_peri_wdata[18] ;
 wire \reg_peri_wdata[19] ;
 wire \reg_peri_wdata[1] ;
 wire \reg_peri_wdata[20] ;
 wire \reg_peri_wdata[21] ;
 wire \reg_peri_wdata[22] ;
 wire \reg_peri_wdata[23] ;
 wire \reg_peri_wdata[24] ;
 wire \reg_peri_wdata[25] ;
 wire \reg_peri_wdata[26] ;
 wire \reg_peri_wdata[27] ;
 wire \reg_peri_wdata[28] ;
 wire \reg_peri_wdata[29] ;
 wire \reg_peri_wdata[2] ;
 wire \reg_peri_wdata[30] ;
 wire \reg_peri_wdata[31] ;
 wire \reg_peri_wdata[3] ;
 wire \reg_peri_wdata[4] ;
 wire \reg_peri_wdata[5] ;
 wire \reg_peri_wdata[6] ;
 wire \reg_peri_wdata[7] ;
 wire \reg_peri_wdata[8] ;
 wire \reg_peri_wdata[9] ;
 wire reg_peri_wr;
 wire rtc_clk;
 wire rtc_intr;
 wire sspim_rst_n;
 wire sspim_sck;
 wire sspim_si;
 wire sspim_so;
 wire \sspim_ssn[0] ;
 wire \sspim_ssn[1] ;
 wire \sspim_ssn[2] ;
 wire \sspim_ssn[3] ;
 wire \uart_rst_n[0] ;
 wire \uart_rst_n[1] ;
 wire \uart_rxd[0] ;
 wire \uart_rxd[1] ;
 wire \uart_txd[0] ;
 wire \uart_txd[1] ;
 wire usb_clk;
 wire usb_dn_i;
 wire usb_dn_o;
 wire usb_dp_i;
 wire usb_dp_o;
 wire usb_intr_o;
 wire usb_oen;
 wire usb_rst_n;

 DSM_core DSM_core (.clk(wb_clk_i),
    .i_wb_cyc(wbs_cyc_i),
    .i_wb_stb(wbs_stb_i),
    .i_wb_we(wbs_we_i),
    .o_wb_ack(wbs_ack_o),
    .reset(wb_rst_i),
    .i_wb_addr({wbs_adr_i[31],
    wbs_adr_i[30],
    wbs_adr_i[29],
    wbs_adr_i[28],
    wbs_adr_i[27],
    wbs_adr_i[26],
    wbs_adr_i[25],
    wbs_adr_i[24],
    wbs_adr_i[23],
    wbs_adr_i[22],
    wbs_adr_i[21],
    wbs_adr_i[20],
    wbs_adr_i[19],
    wbs_adr_i[18],
    wbs_adr_i[17],
    wbs_adr_i[16],
    wbs_adr_i[15],
    wbs_adr_i[14],
    wbs_adr_i[13],
    wbs_adr_i[12],
    wbs_adr_i[11],
    wbs_adr_i[10],
    wbs_adr_i[9],
    wbs_adr_i[8],
    wbs_adr_i[7],
    wbs_adr_i[6],
    wbs_adr_i[5],
    wbs_adr_i[4],
    wbs_adr_i[3],
    wbs_adr_i[2],
    wbs_adr_i[1],
    wbs_adr_i[0]}),
    .i_wb_data({wbs_dat_i[6],
    wbs_dat_i[5],
    wbs_dat_i[4],
    wbs_dat_i[3],
    wbs_dat_i[2],
    wbs_dat_i[1],
    wbs_dat_i[0]}),
    .o_wb_data({wbs_dat_o[4],
    wbs_dat_o[3],
    wbs_dat_o[2],
    wbs_dat_o[1],
    wbs_dat_o[0]}));
 analog_wrapper analog_wrapper ();
 mabrains_logo mabrains_logo ();
 temp_sensor temp_sensor (.clk(user_clock2),
    .i_wb_cyc(wbs_cyc_i),
    .i_wb_stb(wbs_stb_i),
    .i_wb_we(wbs_we_i),
    .o_wb_ack(wbs_ack_o),
    .reset(wb_rst_i),
    .vdd(vdd),
    .vss(vss),
    .i_wb_addr({wbs_adr_i[31],
    wbs_adr_i[30],
    wbs_adr_i[29],
    wbs_adr_i[28],
    wbs_adr_i[27],
    wbs_adr_i[26],
    wbs_adr_i[25],
    wbs_adr_i[24],
    wbs_adr_i[23],
    wbs_adr_i[22],
    wbs_adr_i[21],
    wbs_adr_i[20],
    wbs_adr_i[19],
    wbs_adr_i[18],
    wbs_adr_i[17],
    wbs_adr_i[16],
    wbs_adr_i[15],
    wbs_adr_i[14],
    wbs_adr_i[13],
    wbs_adr_i[12],
    wbs_adr_i[11],
    wbs_adr_i[10],
    wbs_adr_i[9],
    wbs_adr_i[8],
    wbs_adr_i[7],
    wbs_adr_i[6],
    wbs_adr_i[5],
    wbs_adr_i[4],
    wbs_adr_i[3],
    wbs_adr_i[2],
    wbs_adr_i[1],
    wbs_adr_i[0]}),
    .i_wb_data({wbs_dat_i[31],
    wbs_dat_i[30],
    wbs_dat_i[29],
    wbs_dat_i[28],
    wbs_dat_i[27],
    wbs_dat_i[26],
    wbs_dat_i[25],
    wbs_dat_i[24],
    wbs_dat_i[23],
    wbs_dat_i[22],
    wbs_dat_i[21],
    wbs_dat_i[20],
    wbs_dat_i[19],
    wbs_dat_i[18],
    wbs_dat_i[17],
    wbs_dat_i[16],
    wbs_dat_i[15],
    wbs_dat_i[14],
    wbs_dat_i[13],
    wbs_dat_i[12],
    wbs_dat_i[11],
    wbs_dat_i[10],
    wbs_dat_i[9],
    wbs_dat_i[8],
    wbs_dat_i[7],
    wbs_dat_i[6],
    wbs_dat_i[5],
    wbs_dat_i[4],
    wbs_dat_i[3],
    wbs_dat_i[2],
    wbs_dat_i[1],
    wbs_dat_i[0]}),
    .io_oeb({io_oeb[20],
    io_oeb[19],
    io_oeb[18],
    io_oeb[17],
    io_oeb[16],
    io_oeb[15],
    io_oeb[14],
    io_oeb[13]}),
    .io_out({io_out[20],
    io_out[19],
    io_out[18],
    io_out[17],
    io_out[16],
    io_out[15],
    io_out[14],
    io_out[13]}),
    .o_wb_data({wbs_dat_o[7],
    wbs_dat_o[6],
    wbs_dat_o[5],
    wbs_dat_o[4],
    wbs_dat_o[3],
    wbs_dat_o[2],
    wbs_dat_o[1],
    wbs_dat_o[0]}));
 peri_top u_peri (.mclk(wb_clk_i),
    .reg_ack(reg_peri_ack),
    .reg_cs(reg_peri_cs),
    .reg_wr(reg_peri_wr),
    .rtc_clk(rtc_clk),
    .rtc_intr(rtc_intr),
    .s_reset_n(wb_rst_i),
    .vdd(vdd),
    .vss(vss),
    .reg_addr({\reg_peri_addr[10] ,
    \reg_peri_addr[9] ,
    \reg_peri_addr[8] ,
    \reg_peri_addr[7] ,
    \reg_peri_addr[6] ,
    \reg_peri_addr[5] ,
    \reg_peri_addr[4] ,
    \reg_peri_addr[3] ,
    \reg_peri_addr[2] ,
    \reg_peri_addr[1] ,
    \reg_peri_addr[0] }),
    .reg_be({\reg_peri_be[3] ,
    \reg_peri_be[2] ,
    \reg_peri_be[1] ,
    \reg_peri_be[0] }),
    .reg_rdata({\reg_peri_rdata[31] ,
    \reg_peri_rdata[30] ,
    \reg_peri_rdata[29] ,
    \reg_peri_rdata[28] ,
    \reg_peri_rdata[27] ,
    \reg_peri_rdata[26] ,
    \reg_peri_rdata[25] ,
    \reg_peri_rdata[24] ,
    \reg_peri_rdata[23] ,
    \reg_peri_rdata[22] ,
    \reg_peri_rdata[21] ,
    \reg_peri_rdata[20] ,
    \reg_peri_rdata[19] ,
    \reg_peri_rdata[18] ,
    \reg_peri_rdata[17] ,
    \reg_peri_rdata[16] ,
    \reg_peri_rdata[15] ,
    \reg_peri_rdata[14] ,
    \reg_peri_rdata[13] ,
    \reg_peri_rdata[12] ,
    \reg_peri_rdata[11] ,
    \reg_peri_rdata[10] ,
    \reg_peri_rdata[9] ,
    \reg_peri_rdata[8] ,
    \reg_peri_rdata[7] ,
    \reg_peri_rdata[6] ,
    \reg_peri_rdata[5] ,
    \reg_peri_rdata[4] ,
    \reg_peri_rdata[3] ,
    \reg_peri_rdata[2] ,
    \reg_peri_rdata[1] ,
    \reg_peri_rdata[0] }),
    .reg_wdata({\reg_peri_wdata[31] ,
    \reg_peri_wdata[30] ,
    \reg_peri_wdata[29] ,
    \reg_peri_wdata[28] ,
    \reg_peri_wdata[27] ,
    \reg_peri_wdata[26] ,
    \reg_peri_wdata[25] ,
    \reg_peri_wdata[24] ,
    \reg_peri_wdata[23] ,
    \reg_peri_wdata[22] ,
    \reg_peri_wdata[21] ,
    \reg_peri_wdata[20] ,
    \reg_peri_wdata[19] ,
    \reg_peri_wdata[18] ,
    \reg_peri_wdata[17] ,
    \reg_peri_wdata[16] ,
    \reg_peri_wdata[15] ,
    \reg_peri_wdata[14] ,
    \reg_peri_wdata[13] ,
    \reg_peri_wdata[12] ,
    \reg_peri_wdata[11] ,
    \reg_peri_wdata[10] ,
    \reg_peri_wdata[9] ,
    \reg_peri_wdata[8] ,
    \reg_peri_wdata[7] ,
    \reg_peri_wdata[6] ,
    \reg_peri_wdata[5] ,
    \reg_peri_wdata[4] ,
    \reg_peri_wdata[3] ,
    \reg_peri_wdata[2] ,
    \reg_peri_wdata[1] ,
    \reg_peri_wdata[0] }));
 pinmux_top u_pinmux (.e_reset_n(wb_rst_i),
    .i2cm_clk_i(i2cm_clk_i),
    .i2cm_clk_o(i2cm_clk_o),
    .i2cm_clk_oen(i2cm_clk_oen),
    .i2cm_data_i(i2cm_data_i),
    .i2cm_data_o(i2cm_data_o),
    .i2cm_data_oen(i2cm_data_oen),
    .i2cm_intr(i2cm_intr_o),
    .i2cm_rst_n(i2c_rst_n),
    .mclk(wb_clk_i),
    .p_reset_n(wb_rst_i),
    .pulse1m_mclk(pulse1m_mclk),
    .reg_ack(wbs_ack_o),
    .reg_cs(wbs_stb_i),
    .reg_peri_ack(reg_peri_ack),
    .reg_peri_cs(reg_peri_cs),
    .reg_peri_wr(reg_peri_wr),
    .reg_wr(wbs_we_i),
    .rtc_clk(rtc_clk),
    .rtc_intr(rtc_intr),
    .s_reset_n(wb_rst_i),
    .spim_miso(sspim_so),
    .spim_mosi(sspim_si),
    .spim_sck(sspim_sck),
    .sspim_rst_n(sspim_rst_n),
    .usb_clk(usb_clk),
    .usb_dn_i(usb_dn_i),
    .usb_dn_o(usb_dn_o),
    .usb_dp_i(usb_dp_i),
    .usb_dp_o(usb_dp_o),
    .usb_intr(usb_intr_o),
    .usb_oen(usb_oen),
    .usb_rst_n(usb_rst_n),
    .user_clock1(wb_clk_i),
    .user_clock2(user_clock2),
    .vdd(vdd),
    .vss(vss),
    .digital_io_in({io_in[37],
    io_in[36],
    io_in[35],
    io_in[34],
    io_in[33],
    io_in[32],
    io_in[31],
    io_in[30],
    io_in[29],
    io_in[28],
    io_in[27],
    io_in[26],
    io_in[25],
    io_in[24],
    io_in[23],
    io_in[22],
    io_in[21]}),
    .digital_io_oen({io_oeb[37],
    io_oeb[36],
    io_oeb[35],
    io_oeb[34],
    io_oeb[33],
    io_oeb[32],
    io_oeb[31],
    io_oeb[30],
    io_oeb[29],
    io_oeb[28],
    io_oeb[27],
    io_oeb[26],
    io_oeb[25],
    io_oeb[24],
    io_oeb[23],
    io_oeb[22],
    io_oeb[21]}),
    .digital_io_out({io_out[37],
    io_out[36],
    io_out[35],
    io_out[34],
    io_out[33],
    io_out[32],
    io_out[31],
    io_out[30],
    io_out[29],
    io_out[28],
    io_out[27],
    io_out[26],
    io_out[25],
    io_out[24],
    io_out[23],
    io_out[22],
    io_out[21]}),
    .reg_addr({wbs_adr_i[10],
    wbs_adr_i[9],
    wbs_adr_i[8],
    wbs_adr_i[7],
    wbs_adr_i[6],
    wbs_adr_i[5],
    wbs_adr_i[4],
    wbs_adr_i[3],
    wbs_adr_i[2],
    wbs_adr_i[1],
    wbs_adr_i[0]}),
    .reg_be({wbs_sel_i[3],
    wbs_sel_i[2],
    wbs_sel_i[1],
    wbs_sel_i[0]}),
    .reg_peri_addr({\reg_peri_addr[10] ,
    \reg_peri_addr[9] ,
    \reg_peri_addr[8] ,
    \reg_peri_addr[7] ,
    \reg_peri_addr[6] ,
    \reg_peri_addr[5] ,
    \reg_peri_addr[4] ,
    \reg_peri_addr[3] ,
    \reg_peri_addr[2] ,
    \reg_peri_addr[1] ,
    \reg_peri_addr[0] }),
    .reg_peri_be({\reg_peri_be[3] ,
    \reg_peri_be[2] ,
    \reg_peri_be[1] ,
    \reg_peri_be[0] }),
    .reg_peri_rdata({\reg_peri_rdata[31] ,
    \reg_peri_rdata[30] ,
    \reg_peri_rdata[29] ,
    \reg_peri_rdata[28] ,
    \reg_peri_rdata[27] ,
    \reg_peri_rdata[26] ,
    \reg_peri_rdata[25] ,
    \reg_peri_rdata[24] ,
    \reg_peri_rdata[23] ,
    \reg_peri_rdata[22] ,
    \reg_peri_rdata[21] ,
    \reg_peri_rdata[20] ,
    \reg_peri_rdata[19] ,
    \reg_peri_rdata[18] ,
    \reg_peri_rdata[17] ,
    \reg_peri_rdata[16] ,
    \reg_peri_rdata[15] ,
    \reg_peri_rdata[14] ,
    \reg_peri_rdata[13] ,
    \reg_peri_rdata[12] ,
    \reg_peri_rdata[11] ,
    \reg_peri_rdata[10] ,
    \reg_peri_rdata[9] ,
    \reg_peri_rdata[8] ,
    \reg_peri_rdata[7] ,
    \reg_peri_rdata[6] ,
    \reg_peri_rdata[5] ,
    \reg_peri_rdata[4] ,
    \reg_peri_rdata[3] ,
    \reg_peri_rdata[2] ,
    \reg_peri_rdata[1] ,
    \reg_peri_rdata[0] }),
    .reg_peri_wdata({\reg_peri_wdata[31] ,
    \reg_peri_wdata[30] ,
    \reg_peri_wdata[29] ,
    \reg_peri_wdata[28] ,
    \reg_peri_wdata[27] ,
    \reg_peri_wdata[26] ,
    \reg_peri_wdata[25] ,
    \reg_peri_wdata[24] ,
    \reg_peri_wdata[23] ,
    \reg_peri_wdata[22] ,
    \reg_peri_wdata[21] ,
    \reg_peri_wdata[20] ,
    \reg_peri_wdata[19] ,
    \reg_peri_wdata[18] ,
    \reg_peri_wdata[17] ,
    \reg_peri_wdata[16] ,
    \reg_peri_wdata[15] ,
    \reg_peri_wdata[14] ,
    \reg_peri_wdata[13] ,
    \reg_peri_wdata[12] ,
    \reg_peri_wdata[11] ,
    \reg_peri_wdata[10] ,
    \reg_peri_wdata[9] ,
    \reg_peri_wdata[8] ,
    \reg_peri_wdata[7] ,
    \reg_peri_wdata[6] ,
    \reg_peri_wdata[5] ,
    \reg_peri_wdata[4] ,
    \reg_peri_wdata[3] ,
    \reg_peri_wdata[2] ,
    \reg_peri_wdata[1] ,
    \reg_peri_wdata[0] }),
    .reg_rdata({wbs_dat_o[31],
    wbs_dat_o[30],
    wbs_dat_o[29],
    wbs_dat_o[28],
    wbs_dat_o[27],
    wbs_dat_o[26],
    wbs_dat_o[25],
    wbs_dat_o[24],
    wbs_dat_o[23],
    wbs_dat_o[22],
    wbs_dat_o[21],
    wbs_dat_o[20],
    wbs_dat_o[19],
    wbs_dat_o[18],
    wbs_dat_o[17],
    wbs_dat_o[16],
    wbs_dat_o[15],
    wbs_dat_o[14],
    wbs_dat_o[13],
    wbs_dat_o[12],
    wbs_dat_o[11],
    wbs_dat_o[10],
    wbs_dat_o[9],
    wbs_dat_o[8],
    wbs_dat_o[7],
    wbs_dat_o[6],
    wbs_dat_o[5],
    wbs_dat_o[4],
    wbs_dat_o[3],
    wbs_dat_o[2],
    wbs_dat_o[1],
    wbs_dat_o[0]}),
    .reg_wdata({wbs_dat_i[31],
    wbs_dat_i[30],
    wbs_dat_i[29],
    wbs_dat_i[28],
    wbs_dat_i[27],
    wbs_dat_i[26],
    wbs_dat_i[25],
    wbs_dat_i[24],
    wbs_dat_i[23],
    wbs_dat_i[22],
    wbs_dat_i[21],
    wbs_dat_i[20],
    wbs_dat_i[19],
    wbs_dat_i[18],
    wbs_dat_i[17],
    wbs_dat_i[16],
    wbs_dat_i[15],
    wbs_dat_i[14],
    wbs_dat_i[13],
    wbs_dat_i[12],
    wbs_dat_i[11],
    wbs_dat_i[10],
    wbs_dat_i[9],
    wbs_dat_i[8],
    wbs_dat_i[7],
    wbs_dat_i[6],
    wbs_dat_i[5],
    wbs_dat_i[4],
    wbs_dat_i[3],
    wbs_dat_i[2],
    wbs_dat_i[1],
    wbs_dat_i[0]}),
    .spim_ssn({\sspim_ssn[3] ,
    \sspim_ssn[2] ,
    \sspim_ssn[1] ,
    \sspim_ssn[0] }),
    .uart_rst_n({\uart_rst_n[1] ,
    \uart_rst_n[0] }),
    .uart_rxd({\uart_rxd[1] ,
    \uart_rxd[0] }),
    .uart_txd({\uart_txd[1] ,
    \uart_txd[0] }),
    .user_irq({user_irq[2],
    user_irq[1],
    user_irq[0]}));
 uart_i2c_usb_spi_top u_uart_i2c_usb_spi (.app_clk(wb_clk_i),
    .i2c_rstn(i2c_rst_n),
    .i2cm_intr_o(i2cm_intr_o),
    .reg_ack(wbs_ack_o),
    .reg_cs(wbs_stb_i),
    .reg_wr(wbs_we_i),
    .scl_pad_i(i2cm_clk_i),
    .scl_pad_o(i2cm_clk_o),
    .scl_pad_oen_o(i2cm_clk_oen),
    .sda_pad_i(i2cm_data_i),
    .sda_pad_o(i2cm_data_o),
    .sda_padoen_o(i2cm_data_oen),
    .spi_rstn(sspim_rst_n),
    .sspim_sck(sspim_sck),
    .sspim_si(sspim_si),
    .sspim_so(sspim_so),
    .usb_clk(usb_clk),
    .usb_in_dn(usb_dn_i),
    .usb_in_dp(usb_dp_i),
    .usb_intr_o(usb_intr_o),
    .usb_out_dn(usb_dn_o),
    .usb_out_dp(usb_dp_o),
    .usb_out_tx_oen(usb_oen),
    .usb_rstn(usb_rst_n),
    .vdd(vdd),
    .vss(vss),
    .reg_addr({wbs_adr_i[8],
    wbs_adr_i[7],
    wbs_adr_i[6],
    wbs_adr_i[5],
    wbs_adr_i[4],
    wbs_adr_i[3],
    wbs_adr_i[2],
    wbs_adr_i[1],
    wbs_adr_i[0]}),
    .reg_be({wbs_sel_i[3],
    wbs_sel_i[2],
    wbs_sel_i[1],
    wbs_sel_i[0]}),
    .reg_rdata({wbs_dat_o[31],
    wbs_dat_o[30],
    wbs_dat_o[29],
    wbs_dat_o[28],
    wbs_dat_o[27],
    wbs_dat_o[26],
    wbs_dat_o[25],
    wbs_dat_o[24],
    wbs_dat_o[23],
    wbs_dat_o[22],
    wbs_dat_o[21],
    wbs_dat_o[20],
    wbs_dat_o[19],
    wbs_dat_o[18],
    wbs_dat_o[17],
    wbs_dat_o[16],
    wbs_dat_o[15],
    wbs_dat_o[14],
    wbs_dat_o[13],
    wbs_dat_o[12],
    wbs_dat_o[11],
    wbs_dat_o[10],
    wbs_dat_o[9],
    wbs_dat_o[8],
    wbs_dat_o[7],
    wbs_dat_o[6],
    wbs_dat_o[5],
    wbs_dat_o[4],
    wbs_dat_o[3],
    wbs_dat_o[2],
    wbs_dat_o[1],
    wbs_dat_o[0]}),
    .reg_wdata({wbs_dat_i[31],
    wbs_dat_i[30],
    wbs_dat_i[29],
    wbs_dat_i[28],
    wbs_dat_i[27],
    wbs_dat_i[26],
    wbs_dat_i[25],
    wbs_dat_i[24],
    wbs_dat_i[23],
    wbs_dat_i[22],
    wbs_dat_i[21],
    wbs_dat_i[20],
    wbs_dat_i[19],
    wbs_dat_i[18],
    wbs_dat_i[17],
    wbs_dat_i[16],
    wbs_dat_i[15],
    wbs_dat_i[14],
    wbs_dat_i[13],
    wbs_dat_i[12],
    wbs_dat_i[11],
    wbs_dat_i[10],
    wbs_dat_i[9],
    wbs_dat_i[8],
    wbs_dat_i[7],
    wbs_dat_i[6],
    wbs_dat_i[5],
    wbs_dat_i[4],
    wbs_dat_i[3],
    wbs_dat_i[2],
    wbs_dat_i[1],
    wbs_dat_i[0]}),
    .sspim_ssn({\sspim_ssn[3] ,
    \sspim_ssn[2] ,
    \sspim_ssn[1] ,
    \sspim_ssn[0] }),
    .uart_rstn({\uart_rst_n[1] ,
    \uart_rst_n[0] }),
    .uart_rxd({\uart_rxd[1] ,
    \uart_rxd[0] }),
    .uart_txd({\uart_txd[1] ,
    \uart_txd[0] }));
 wb_buttons_leds wb_buttons_leds (.clk(wb_clk_i),
    .clk2(user_clock2),
    .i_wb_cyc(wbs_cyc_i),
    .i_wb_stb(wbs_stb_i),
    .i_wb_we(wbs_we_i),
    .o_wb_ack(wbs_ack_o),
    .reset(wb_rst_i),
    .vdd(vdd),
    .vss(vss),
    .buttons({io_in[6],
    io_in[5]}),
    .buttons_enb({io_oeb[6],
    io_oeb[5]}),
    .i_wb_addr({wbs_adr_i[31],
    wbs_adr_i[30],
    wbs_adr_i[29],
    wbs_adr_i[28],
    wbs_adr_i[27],
    wbs_adr_i[26],
    wbs_adr_i[25],
    wbs_adr_i[24],
    wbs_adr_i[23],
    wbs_adr_i[22],
    wbs_adr_i[21],
    wbs_adr_i[20],
    wbs_adr_i[19],
    wbs_adr_i[18],
    wbs_adr_i[17],
    wbs_adr_i[16],
    wbs_adr_i[15],
    wbs_adr_i[14],
    wbs_adr_i[13],
    wbs_adr_i[12],
    wbs_adr_i[11],
    wbs_adr_i[10],
    wbs_adr_i[9],
    wbs_adr_i[8],
    wbs_adr_i[7],
    wbs_adr_i[6],
    wbs_adr_i[5],
    wbs_adr_i[4],
    wbs_adr_i[3],
    wbs_adr_i[2],
    wbs_adr_i[1],
    wbs_adr_i[0]}),
    .i_wb_data({wbs_dat_i[1],
    wbs_dat_i[0]}),
    .led_enb({io_oeb[8],
    io_oeb[7]}),
    .leds({io_out[8],
    io_out[7]}),
    .o_wb_data({wbs_dat_o[31],
    wbs_dat_o[30],
    wbs_dat_o[29],
    wbs_dat_o[28],
    wbs_dat_o[27],
    wbs_dat_o[26],
    wbs_dat_o[25],
    wbs_dat_o[24],
    wbs_dat_o[23],
    wbs_dat_o[22],
    wbs_dat_o[21],
    wbs_dat_o[20],
    wbs_dat_o[19],
    wbs_dat_o[18],
    wbs_dat_o[17],
    wbs_dat_o[16],
    wbs_dat_o[15],
    wbs_dat_o[14],
    wbs_dat_o[13],
    wbs_dat_o[12],
    wbs_dat_o[11],
    wbs_dat_o[10],
    wbs_dat_o[9],
    wbs_dat_o[8],
    wbs_dat_o[7],
    wbs_dat_o[6],
    wbs_dat_o[5],
    wbs_dat_o[4],
    wbs_dat_o[3],
    wbs_dat_o[2],
    wbs_dat_o[1],
    wbs_dat_o[0]}),
    .xtal_clk({io_out[10],
    io_out[9]}),
    .xtal_clk_enb({io_oeb[10],
    io_oeb[9]}));
endmodule
